
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_rem IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END mgc_rem;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_rem IS
BEGIN
  z <= std_logic_vector(unsigned(a) rem unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) rem   signed(b));
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_div IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END mgc_div;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_div IS
BEGIN
  z <= std_logic_vector(unsigned(a) / unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) /   signed(b));
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Thu Jul  1 00:56:08 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen;

ARCHITECTURE v43 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
    STAGE_LOOP_C_8_tr0 : IN STD_LOGIC;
    modExp_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_1_tr0 : IN STD_LOGIC;
    COMP_LOOP_1_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_62_tr0 : IN STD_LOGIC;
    COMP_LOOP_2_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_124_tr0 : IN STD_LOGIC;
    COMP_LOOP_3_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_186_tr0 : IN STD_LOGIC;
    COMP_LOOP_4_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_248_tr0 : IN STD_LOGIC;
    COMP_LOOP_5_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_310_tr0 : IN STD_LOGIC;
    COMP_LOOP_6_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_372_tr0 : IN STD_LOGIC;
    COMP_LOOP_7_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_434_tr0 : IN STD_LOGIC;
    COMP_LOOP_8_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_496_tr0 : IN STD_LOGIC;
    COMP_LOOP_9_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_558_tr0 : IN STD_LOGIC;
    COMP_LOOP_10_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_620_tr0 : IN STD_LOGIC;
    COMP_LOOP_11_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_682_tr0 : IN STD_LOGIC;
    COMP_LOOP_12_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_744_tr0 : IN STD_LOGIC;
    COMP_LOOP_13_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_806_tr0 : IN STD_LOGIC;
    COMP_LOOP_14_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_868_tr0 : IN STD_LOGIC;
    COMP_LOOP_15_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_930_tr0 : IN STD_LOGIC;
    COMP_LOOP_16_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_992_tr0 : IN STD_LOGIC;
    VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_9_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIT_core_core_fsm;

ARCHITECTURE v43 OF inPlaceNTT_DIT_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  TYPE inPlaceNTT_DIT_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, STAGE_LOOP_C_1,
      STAGE_LOOP_C_2, STAGE_LOOP_C_3, STAGE_LOOP_C_4, STAGE_LOOP_C_5, STAGE_LOOP_C_6,
      STAGE_LOOP_C_7, STAGE_LOOP_C_8, modExp_while_C_0, modExp_while_C_1, modExp_while_C_2,
      modExp_while_C_3, modExp_while_C_4, modExp_while_C_5, modExp_while_C_6, modExp_while_C_7,
      modExp_while_C_8, modExp_while_C_9, modExp_while_C_10, modExp_while_C_11, modExp_while_C_12,
      modExp_while_C_13, modExp_while_C_14, modExp_while_C_15, modExp_while_C_16,
      modExp_while_C_17, modExp_while_C_18, modExp_while_C_19, modExp_while_C_20,
      modExp_while_C_21, modExp_while_C_22, modExp_while_C_23, modExp_while_C_24,
      modExp_while_C_25, modExp_while_C_26, modExp_while_C_27, modExp_while_C_28,
      modExp_while_C_29, modExp_while_C_30, modExp_while_C_31, modExp_while_C_32,
      modExp_while_C_33, modExp_while_C_34, modExp_while_C_35, modExp_while_C_36,
      modExp_while_C_37, modExp_while_C_38, COMP_LOOP_C_0, COMP_LOOP_C_1, COMP_LOOP_1_modExp_1_while_C_0,
      COMP_LOOP_1_modExp_1_while_C_1, COMP_LOOP_1_modExp_1_while_C_2, COMP_LOOP_1_modExp_1_while_C_3,
      COMP_LOOP_1_modExp_1_while_C_4, COMP_LOOP_1_modExp_1_while_C_5, COMP_LOOP_1_modExp_1_while_C_6,
      COMP_LOOP_1_modExp_1_while_C_7, COMP_LOOP_1_modExp_1_while_C_8, COMP_LOOP_1_modExp_1_while_C_9,
      COMP_LOOP_1_modExp_1_while_C_10, COMP_LOOP_1_modExp_1_while_C_11, COMP_LOOP_1_modExp_1_while_C_12,
      COMP_LOOP_1_modExp_1_while_C_13, COMP_LOOP_1_modExp_1_while_C_14, COMP_LOOP_1_modExp_1_while_C_15,
      COMP_LOOP_1_modExp_1_while_C_16, COMP_LOOP_1_modExp_1_while_C_17, COMP_LOOP_1_modExp_1_while_C_18,
      COMP_LOOP_1_modExp_1_while_C_19, COMP_LOOP_1_modExp_1_while_C_20, COMP_LOOP_1_modExp_1_while_C_21,
      COMP_LOOP_1_modExp_1_while_C_22, COMP_LOOP_1_modExp_1_while_C_23, COMP_LOOP_1_modExp_1_while_C_24,
      COMP_LOOP_1_modExp_1_while_C_25, COMP_LOOP_1_modExp_1_while_C_26, COMP_LOOP_1_modExp_1_while_C_27,
      COMP_LOOP_1_modExp_1_while_C_28, COMP_LOOP_1_modExp_1_while_C_29, COMP_LOOP_1_modExp_1_while_C_30,
      COMP_LOOP_1_modExp_1_while_C_31, COMP_LOOP_1_modExp_1_while_C_32, COMP_LOOP_1_modExp_1_while_C_33,
      COMP_LOOP_1_modExp_1_while_C_34, COMP_LOOP_1_modExp_1_while_C_35, COMP_LOOP_1_modExp_1_while_C_36,
      COMP_LOOP_1_modExp_1_while_C_37, COMP_LOOP_1_modExp_1_while_C_38, COMP_LOOP_C_2,
      COMP_LOOP_C_3, COMP_LOOP_C_4, COMP_LOOP_C_5, COMP_LOOP_C_6, COMP_LOOP_C_7,
      COMP_LOOP_C_8, COMP_LOOP_C_9, COMP_LOOP_C_10, COMP_LOOP_C_11, COMP_LOOP_C_12,
      COMP_LOOP_C_13, COMP_LOOP_C_14, COMP_LOOP_C_15, COMP_LOOP_C_16, COMP_LOOP_C_17,
      COMP_LOOP_C_18, COMP_LOOP_C_19, COMP_LOOP_C_20, COMP_LOOP_C_21, COMP_LOOP_C_22,
      COMP_LOOP_C_23, COMP_LOOP_C_24, COMP_LOOP_C_25, COMP_LOOP_C_26, COMP_LOOP_C_27,
      COMP_LOOP_C_28, COMP_LOOP_C_29, COMP_LOOP_C_30, COMP_LOOP_C_31, COMP_LOOP_C_32,
      COMP_LOOP_C_33, COMP_LOOP_C_34, COMP_LOOP_C_35, COMP_LOOP_C_36, COMP_LOOP_C_37,
      COMP_LOOP_C_38, COMP_LOOP_C_39, COMP_LOOP_C_40, COMP_LOOP_C_41, COMP_LOOP_C_42,
      COMP_LOOP_C_43, COMP_LOOP_C_44, COMP_LOOP_C_45, COMP_LOOP_C_46, COMP_LOOP_C_47,
      COMP_LOOP_C_48, COMP_LOOP_C_49, COMP_LOOP_C_50, COMP_LOOP_C_51, COMP_LOOP_C_52,
      COMP_LOOP_C_53, COMP_LOOP_C_54, COMP_LOOP_C_55, COMP_LOOP_C_56, COMP_LOOP_C_57,
      COMP_LOOP_C_58, COMP_LOOP_C_59, COMP_LOOP_C_60, COMP_LOOP_C_61, COMP_LOOP_C_62,
      COMP_LOOP_C_63, COMP_LOOP_2_modExp_1_while_C_0, COMP_LOOP_2_modExp_1_while_C_1,
      COMP_LOOP_2_modExp_1_while_C_2, COMP_LOOP_2_modExp_1_while_C_3, COMP_LOOP_2_modExp_1_while_C_4,
      COMP_LOOP_2_modExp_1_while_C_5, COMP_LOOP_2_modExp_1_while_C_6, COMP_LOOP_2_modExp_1_while_C_7,
      COMP_LOOP_2_modExp_1_while_C_8, COMP_LOOP_2_modExp_1_while_C_9, COMP_LOOP_2_modExp_1_while_C_10,
      COMP_LOOP_2_modExp_1_while_C_11, COMP_LOOP_2_modExp_1_while_C_12, COMP_LOOP_2_modExp_1_while_C_13,
      COMP_LOOP_2_modExp_1_while_C_14, COMP_LOOP_2_modExp_1_while_C_15, COMP_LOOP_2_modExp_1_while_C_16,
      COMP_LOOP_2_modExp_1_while_C_17, COMP_LOOP_2_modExp_1_while_C_18, COMP_LOOP_2_modExp_1_while_C_19,
      COMP_LOOP_2_modExp_1_while_C_20, COMP_LOOP_2_modExp_1_while_C_21, COMP_LOOP_2_modExp_1_while_C_22,
      COMP_LOOP_2_modExp_1_while_C_23, COMP_LOOP_2_modExp_1_while_C_24, COMP_LOOP_2_modExp_1_while_C_25,
      COMP_LOOP_2_modExp_1_while_C_26, COMP_LOOP_2_modExp_1_while_C_27, COMP_LOOP_2_modExp_1_while_C_28,
      COMP_LOOP_2_modExp_1_while_C_29, COMP_LOOP_2_modExp_1_while_C_30, COMP_LOOP_2_modExp_1_while_C_31,
      COMP_LOOP_2_modExp_1_while_C_32, COMP_LOOP_2_modExp_1_while_C_33, COMP_LOOP_2_modExp_1_while_C_34,
      COMP_LOOP_2_modExp_1_while_C_35, COMP_LOOP_2_modExp_1_while_C_36, COMP_LOOP_2_modExp_1_while_C_37,
      COMP_LOOP_2_modExp_1_while_C_38, COMP_LOOP_C_64, COMP_LOOP_C_65, COMP_LOOP_C_66,
      COMP_LOOP_C_67, COMP_LOOP_C_68, COMP_LOOP_C_69, COMP_LOOP_C_70, COMP_LOOP_C_71,
      COMP_LOOP_C_72, COMP_LOOP_C_73, COMP_LOOP_C_74, COMP_LOOP_C_75, COMP_LOOP_C_76,
      COMP_LOOP_C_77, COMP_LOOP_C_78, COMP_LOOP_C_79, COMP_LOOP_C_80, COMP_LOOP_C_81,
      COMP_LOOP_C_82, COMP_LOOP_C_83, COMP_LOOP_C_84, COMP_LOOP_C_85, COMP_LOOP_C_86,
      COMP_LOOP_C_87, COMP_LOOP_C_88, COMP_LOOP_C_89, COMP_LOOP_C_90, COMP_LOOP_C_91,
      COMP_LOOP_C_92, COMP_LOOP_C_93, COMP_LOOP_C_94, COMP_LOOP_C_95, COMP_LOOP_C_96,
      COMP_LOOP_C_97, COMP_LOOP_C_98, COMP_LOOP_C_99, COMP_LOOP_C_100, COMP_LOOP_C_101,
      COMP_LOOP_C_102, COMP_LOOP_C_103, COMP_LOOP_C_104, COMP_LOOP_C_105, COMP_LOOP_C_106,
      COMP_LOOP_C_107, COMP_LOOP_C_108, COMP_LOOP_C_109, COMP_LOOP_C_110, COMP_LOOP_C_111,
      COMP_LOOP_C_112, COMP_LOOP_C_113, COMP_LOOP_C_114, COMP_LOOP_C_115, COMP_LOOP_C_116,
      COMP_LOOP_C_117, COMP_LOOP_C_118, COMP_LOOP_C_119, COMP_LOOP_C_120, COMP_LOOP_C_121,
      COMP_LOOP_C_122, COMP_LOOP_C_123, COMP_LOOP_C_124, COMP_LOOP_C_125, COMP_LOOP_3_modExp_1_while_C_0,
      COMP_LOOP_3_modExp_1_while_C_1, COMP_LOOP_3_modExp_1_while_C_2, COMP_LOOP_3_modExp_1_while_C_3,
      COMP_LOOP_3_modExp_1_while_C_4, COMP_LOOP_3_modExp_1_while_C_5, COMP_LOOP_3_modExp_1_while_C_6,
      COMP_LOOP_3_modExp_1_while_C_7, COMP_LOOP_3_modExp_1_while_C_8, COMP_LOOP_3_modExp_1_while_C_9,
      COMP_LOOP_3_modExp_1_while_C_10, COMP_LOOP_3_modExp_1_while_C_11, COMP_LOOP_3_modExp_1_while_C_12,
      COMP_LOOP_3_modExp_1_while_C_13, COMP_LOOP_3_modExp_1_while_C_14, COMP_LOOP_3_modExp_1_while_C_15,
      COMP_LOOP_3_modExp_1_while_C_16, COMP_LOOP_3_modExp_1_while_C_17, COMP_LOOP_3_modExp_1_while_C_18,
      COMP_LOOP_3_modExp_1_while_C_19, COMP_LOOP_3_modExp_1_while_C_20, COMP_LOOP_3_modExp_1_while_C_21,
      COMP_LOOP_3_modExp_1_while_C_22, COMP_LOOP_3_modExp_1_while_C_23, COMP_LOOP_3_modExp_1_while_C_24,
      COMP_LOOP_3_modExp_1_while_C_25, COMP_LOOP_3_modExp_1_while_C_26, COMP_LOOP_3_modExp_1_while_C_27,
      COMP_LOOP_3_modExp_1_while_C_28, COMP_LOOP_3_modExp_1_while_C_29, COMP_LOOP_3_modExp_1_while_C_30,
      COMP_LOOP_3_modExp_1_while_C_31, COMP_LOOP_3_modExp_1_while_C_32, COMP_LOOP_3_modExp_1_while_C_33,
      COMP_LOOP_3_modExp_1_while_C_34, COMP_LOOP_3_modExp_1_while_C_35, COMP_LOOP_3_modExp_1_while_C_36,
      COMP_LOOP_3_modExp_1_while_C_37, COMP_LOOP_3_modExp_1_while_C_38, COMP_LOOP_C_126,
      COMP_LOOP_C_127, COMP_LOOP_C_128, COMP_LOOP_C_129, COMP_LOOP_C_130, COMP_LOOP_C_131,
      COMP_LOOP_C_132, COMP_LOOP_C_133, COMP_LOOP_C_134, COMP_LOOP_C_135, COMP_LOOP_C_136,
      COMP_LOOP_C_137, COMP_LOOP_C_138, COMP_LOOP_C_139, COMP_LOOP_C_140, COMP_LOOP_C_141,
      COMP_LOOP_C_142, COMP_LOOP_C_143, COMP_LOOP_C_144, COMP_LOOP_C_145, COMP_LOOP_C_146,
      COMP_LOOP_C_147, COMP_LOOP_C_148, COMP_LOOP_C_149, COMP_LOOP_C_150, COMP_LOOP_C_151,
      COMP_LOOP_C_152, COMP_LOOP_C_153, COMP_LOOP_C_154, COMP_LOOP_C_155, COMP_LOOP_C_156,
      COMP_LOOP_C_157, COMP_LOOP_C_158, COMP_LOOP_C_159, COMP_LOOP_C_160, COMP_LOOP_C_161,
      COMP_LOOP_C_162, COMP_LOOP_C_163, COMP_LOOP_C_164, COMP_LOOP_C_165, COMP_LOOP_C_166,
      COMP_LOOP_C_167, COMP_LOOP_C_168, COMP_LOOP_C_169, COMP_LOOP_C_170, COMP_LOOP_C_171,
      COMP_LOOP_C_172, COMP_LOOP_C_173, COMP_LOOP_C_174, COMP_LOOP_C_175, COMP_LOOP_C_176,
      COMP_LOOP_C_177, COMP_LOOP_C_178, COMP_LOOP_C_179, COMP_LOOP_C_180, COMP_LOOP_C_181,
      COMP_LOOP_C_182, COMP_LOOP_C_183, COMP_LOOP_C_184, COMP_LOOP_C_185, COMP_LOOP_C_186,
      COMP_LOOP_C_187, COMP_LOOP_4_modExp_1_while_C_0, COMP_LOOP_4_modExp_1_while_C_1,
      COMP_LOOP_4_modExp_1_while_C_2, COMP_LOOP_4_modExp_1_while_C_3, COMP_LOOP_4_modExp_1_while_C_4,
      COMP_LOOP_4_modExp_1_while_C_5, COMP_LOOP_4_modExp_1_while_C_6, COMP_LOOP_4_modExp_1_while_C_7,
      COMP_LOOP_4_modExp_1_while_C_8, COMP_LOOP_4_modExp_1_while_C_9, COMP_LOOP_4_modExp_1_while_C_10,
      COMP_LOOP_4_modExp_1_while_C_11, COMP_LOOP_4_modExp_1_while_C_12, COMP_LOOP_4_modExp_1_while_C_13,
      COMP_LOOP_4_modExp_1_while_C_14, COMP_LOOP_4_modExp_1_while_C_15, COMP_LOOP_4_modExp_1_while_C_16,
      COMP_LOOP_4_modExp_1_while_C_17, COMP_LOOP_4_modExp_1_while_C_18, COMP_LOOP_4_modExp_1_while_C_19,
      COMP_LOOP_4_modExp_1_while_C_20, COMP_LOOP_4_modExp_1_while_C_21, COMP_LOOP_4_modExp_1_while_C_22,
      COMP_LOOP_4_modExp_1_while_C_23, COMP_LOOP_4_modExp_1_while_C_24, COMP_LOOP_4_modExp_1_while_C_25,
      COMP_LOOP_4_modExp_1_while_C_26, COMP_LOOP_4_modExp_1_while_C_27, COMP_LOOP_4_modExp_1_while_C_28,
      COMP_LOOP_4_modExp_1_while_C_29, COMP_LOOP_4_modExp_1_while_C_30, COMP_LOOP_4_modExp_1_while_C_31,
      COMP_LOOP_4_modExp_1_while_C_32, COMP_LOOP_4_modExp_1_while_C_33, COMP_LOOP_4_modExp_1_while_C_34,
      COMP_LOOP_4_modExp_1_while_C_35, COMP_LOOP_4_modExp_1_while_C_36, COMP_LOOP_4_modExp_1_while_C_37,
      COMP_LOOP_4_modExp_1_while_C_38, COMP_LOOP_C_188, COMP_LOOP_C_189, COMP_LOOP_C_190,
      COMP_LOOP_C_191, COMP_LOOP_C_192, COMP_LOOP_C_193, COMP_LOOP_C_194, COMP_LOOP_C_195,
      COMP_LOOP_C_196, COMP_LOOP_C_197, COMP_LOOP_C_198, COMP_LOOP_C_199, COMP_LOOP_C_200,
      COMP_LOOP_C_201, COMP_LOOP_C_202, COMP_LOOP_C_203, COMP_LOOP_C_204, COMP_LOOP_C_205,
      COMP_LOOP_C_206, COMP_LOOP_C_207, COMP_LOOP_C_208, COMP_LOOP_C_209, COMP_LOOP_C_210,
      COMP_LOOP_C_211, COMP_LOOP_C_212, COMP_LOOP_C_213, COMP_LOOP_C_214, COMP_LOOP_C_215,
      COMP_LOOP_C_216, COMP_LOOP_C_217, COMP_LOOP_C_218, COMP_LOOP_C_219, COMP_LOOP_C_220,
      COMP_LOOP_C_221, COMP_LOOP_C_222, COMP_LOOP_C_223, COMP_LOOP_C_224, COMP_LOOP_C_225,
      COMP_LOOP_C_226, COMP_LOOP_C_227, COMP_LOOP_C_228, COMP_LOOP_C_229, COMP_LOOP_C_230,
      COMP_LOOP_C_231, COMP_LOOP_C_232, COMP_LOOP_C_233, COMP_LOOP_C_234, COMP_LOOP_C_235,
      COMP_LOOP_C_236, COMP_LOOP_C_237, COMP_LOOP_C_238, COMP_LOOP_C_239, COMP_LOOP_C_240,
      COMP_LOOP_C_241, COMP_LOOP_C_242, COMP_LOOP_C_243, COMP_LOOP_C_244, COMP_LOOP_C_245,
      COMP_LOOP_C_246, COMP_LOOP_C_247, COMP_LOOP_C_248, COMP_LOOP_C_249, COMP_LOOP_5_modExp_1_while_C_0,
      COMP_LOOP_5_modExp_1_while_C_1, COMP_LOOP_5_modExp_1_while_C_2, COMP_LOOP_5_modExp_1_while_C_3,
      COMP_LOOP_5_modExp_1_while_C_4, COMP_LOOP_5_modExp_1_while_C_5, COMP_LOOP_5_modExp_1_while_C_6,
      COMP_LOOP_5_modExp_1_while_C_7, COMP_LOOP_5_modExp_1_while_C_8, COMP_LOOP_5_modExp_1_while_C_9,
      COMP_LOOP_5_modExp_1_while_C_10, COMP_LOOP_5_modExp_1_while_C_11, COMP_LOOP_5_modExp_1_while_C_12,
      COMP_LOOP_5_modExp_1_while_C_13, COMP_LOOP_5_modExp_1_while_C_14, COMP_LOOP_5_modExp_1_while_C_15,
      COMP_LOOP_5_modExp_1_while_C_16, COMP_LOOP_5_modExp_1_while_C_17, COMP_LOOP_5_modExp_1_while_C_18,
      COMP_LOOP_5_modExp_1_while_C_19, COMP_LOOP_5_modExp_1_while_C_20, COMP_LOOP_5_modExp_1_while_C_21,
      COMP_LOOP_5_modExp_1_while_C_22, COMP_LOOP_5_modExp_1_while_C_23, COMP_LOOP_5_modExp_1_while_C_24,
      COMP_LOOP_5_modExp_1_while_C_25, COMP_LOOP_5_modExp_1_while_C_26, COMP_LOOP_5_modExp_1_while_C_27,
      COMP_LOOP_5_modExp_1_while_C_28, COMP_LOOP_5_modExp_1_while_C_29, COMP_LOOP_5_modExp_1_while_C_30,
      COMP_LOOP_5_modExp_1_while_C_31, COMP_LOOP_5_modExp_1_while_C_32, COMP_LOOP_5_modExp_1_while_C_33,
      COMP_LOOP_5_modExp_1_while_C_34, COMP_LOOP_5_modExp_1_while_C_35, COMP_LOOP_5_modExp_1_while_C_36,
      COMP_LOOP_5_modExp_1_while_C_37, COMP_LOOP_5_modExp_1_while_C_38, COMP_LOOP_C_250,
      COMP_LOOP_C_251, COMP_LOOP_C_252, COMP_LOOP_C_253, COMP_LOOP_C_254, COMP_LOOP_C_255,
      COMP_LOOP_C_256, COMP_LOOP_C_257, COMP_LOOP_C_258, COMP_LOOP_C_259, COMP_LOOP_C_260,
      COMP_LOOP_C_261, COMP_LOOP_C_262, COMP_LOOP_C_263, COMP_LOOP_C_264, COMP_LOOP_C_265,
      COMP_LOOP_C_266, COMP_LOOP_C_267, COMP_LOOP_C_268, COMP_LOOP_C_269, COMP_LOOP_C_270,
      COMP_LOOP_C_271, COMP_LOOP_C_272, COMP_LOOP_C_273, COMP_LOOP_C_274, COMP_LOOP_C_275,
      COMP_LOOP_C_276, COMP_LOOP_C_277, COMP_LOOP_C_278, COMP_LOOP_C_279, COMP_LOOP_C_280,
      COMP_LOOP_C_281, COMP_LOOP_C_282, COMP_LOOP_C_283, COMP_LOOP_C_284, COMP_LOOP_C_285,
      COMP_LOOP_C_286, COMP_LOOP_C_287, COMP_LOOP_C_288, COMP_LOOP_C_289, COMP_LOOP_C_290,
      COMP_LOOP_C_291, COMP_LOOP_C_292, COMP_LOOP_C_293, COMP_LOOP_C_294, COMP_LOOP_C_295,
      COMP_LOOP_C_296, COMP_LOOP_C_297, COMP_LOOP_C_298, COMP_LOOP_C_299, COMP_LOOP_C_300,
      COMP_LOOP_C_301, COMP_LOOP_C_302, COMP_LOOP_C_303, COMP_LOOP_C_304, COMP_LOOP_C_305,
      COMP_LOOP_C_306, COMP_LOOP_C_307, COMP_LOOP_C_308, COMP_LOOP_C_309, COMP_LOOP_C_310,
      COMP_LOOP_C_311, COMP_LOOP_6_modExp_1_while_C_0, COMP_LOOP_6_modExp_1_while_C_1,
      COMP_LOOP_6_modExp_1_while_C_2, COMP_LOOP_6_modExp_1_while_C_3, COMP_LOOP_6_modExp_1_while_C_4,
      COMP_LOOP_6_modExp_1_while_C_5, COMP_LOOP_6_modExp_1_while_C_6, COMP_LOOP_6_modExp_1_while_C_7,
      COMP_LOOP_6_modExp_1_while_C_8, COMP_LOOP_6_modExp_1_while_C_9, COMP_LOOP_6_modExp_1_while_C_10,
      COMP_LOOP_6_modExp_1_while_C_11, COMP_LOOP_6_modExp_1_while_C_12, COMP_LOOP_6_modExp_1_while_C_13,
      COMP_LOOP_6_modExp_1_while_C_14, COMP_LOOP_6_modExp_1_while_C_15, COMP_LOOP_6_modExp_1_while_C_16,
      COMP_LOOP_6_modExp_1_while_C_17, COMP_LOOP_6_modExp_1_while_C_18, COMP_LOOP_6_modExp_1_while_C_19,
      COMP_LOOP_6_modExp_1_while_C_20, COMP_LOOP_6_modExp_1_while_C_21, COMP_LOOP_6_modExp_1_while_C_22,
      COMP_LOOP_6_modExp_1_while_C_23, COMP_LOOP_6_modExp_1_while_C_24, COMP_LOOP_6_modExp_1_while_C_25,
      COMP_LOOP_6_modExp_1_while_C_26, COMP_LOOP_6_modExp_1_while_C_27, COMP_LOOP_6_modExp_1_while_C_28,
      COMP_LOOP_6_modExp_1_while_C_29, COMP_LOOP_6_modExp_1_while_C_30, COMP_LOOP_6_modExp_1_while_C_31,
      COMP_LOOP_6_modExp_1_while_C_32, COMP_LOOP_6_modExp_1_while_C_33, COMP_LOOP_6_modExp_1_while_C_34,
      COMP_LOOP_6_modExp_1_while_C_35, COMP_LOOP_6_modExp_1_while_C_36, COMP_LOOP_6_modExp_1_while_C_37,
      COMP_LOOP_6_modExp_1_while_C_38, COMP_LOOP_C_312, COMP_LOOP_C_313, COMP_LOOP_C_314,
      COMP_LOOP_C_315, COMP_LOOP_C_316, COMP_LOOP_C_317, COMP_LOOP_C_318, COMP_LOOP_C_319,
      COMP_LOOP_C_320, COMP_LOOP_C_321, COMP_LOOP_C_322, COMP_LOOP_C_323, COMP_LOOP_C_324,
      COMP_LOOP_C_325, COMP_LOOP_C_326, COMP_LOOP_C_327, COMP_LOOP_C_328, COMP_LOOP_C_329,
      COMP_LOOP_C_330, COMP_LOOP_C_331, COMP_LOOP_C_332, COMP_LOOP_C_333, COMP_LOOP_C_334,
      COMP_LOOP_C_335, COMP_LOOP_C_336, COMP_LOOP_C_337, COMP_LOOP_C_338, COMP_LOOP_C_339,
      COMP_LOOP_C_340, COMP_LOOP_C_341, COMP_LOOP_C_342, COMP_LOOP_C_343, COMP_LOOP_C_344,
      COMP_LOOP_C_345, COMP_LOOP_C_346, COMP_LOOP_C_347, COMP_LOOP_C_348, COMP_LOOP_C_349,
      COMP_LOOP_C_350, COMP_LOOP_C_351, COMP_LOOP_C_352, COMP_LOOP_C_353, COMP_LOOP_C_354,
      COMP_LOOP_C_355, COMP_LOOP_C_356, COMP_LOOP_C_357, COMP_LOOP_C_358, COMP_LOOP_C_359,
      COMP_LOOP_C_360, COMP_LOOP_C_361, COMP_LOOP_C_362, COMP_LOOP_C_363, COMP_LOOP_C_364,
      COMP_LOOP_C_365, COMP_LOOP_C_366, COMP_LOOP_C_367, COMP_LOOP_C_368, COMP_LOOP_C_369,
      COMP_LOOP_C_370, COMP_LOOP_C_371, COMP_LOOP_C_372, COMP_LOOP_C_373, COMP_LOOP_7_modExp_1_while_C_0,
      COMP_LOOP_7_modExp_1_while_C_1, COMP_LOOP_7_modExp_1_while_C_2, COMP_LOOP_7_modExp_1_while_C_3,
      COMP_LOOP_7_modExp_1_while_C_4, COMP_LOOP_7_modExp_1_while_C_5, COMP_LOOP_7_modExp_1_while_C_6,
      COMP_LOOP_7_modExp_1_while_C_7, COMP_LOOP_7_modExp_1_while_C_8, COMP_LOOP_7_modExp_1_while_C_9,
      COMP_LOOP_7_modExp_1_while_C_10, COMP_LOOP_7_modExp_1_while_C_11, COMP_LOOP_7_modExp_1_while_C_12,
      COMP_LOOP_7_modExp_1_while_C_13, COMP_LOOP_7_modExp_1_while_C_14, COMP_LOOP_7_modExp_1_while_C_15,
      COMP_LOOP_7_modExp_1_while_C_16, COMP_LOOP_7_modExp_1_while_C_17, COMP_LOOP_7_modExp_1_while_C_18,
      COMP_LOOP_7_modExp_1_while_C_19, COMP_LOOP_7_modExp_1_while_C_20, COMP_LOOP_7_modExp_1_while_C_21,
      COMP_LOOP_7_modExp_1_while_C_22, COMP_LOOP_7_modExp_1_while_C_23, COMP_LOOP_7_modExp_1_while_C_24,
      COMP_LOOP_7_modExp_1_while_C_25, COMP_LOOP_7_modExp_1_while_C_26, COMP_LOOP_7_modExp_1_while_C_27,
      COMP_LOOP_7_modExp_1_while_C_28, COMP_LOOP_7_modExp_1_while_C_29, COMP_LOOP_7_modExp_1_while_C_30,
      COMP_LOOP_7_modExp_1_while_C_31, COMP_LOOP_7_modExp_1_while_C_32, COMP_LOOP_7_modExp_1_while_C_33,
      COMP_LOOP_7_modExp_1_while_C_34, COMP_LOOP_7_modExp_1_while_C_35, COMP_LOOP_7_modExp_1_while_C_36,
      COMP_LOOP_7_modExp_1_while_C_37, COMP_LOOP_7_modExp_1_while_C_38, COMP_LOOP_C_374,
      COMP_LOOP_C_375, COMP_LOOP_C_376, COMP_LOOP_C_377, COMP_LOOP_C_378, COMP_LOOP_C_379,
      COMP_LOOP_C_380, COMP_LOOP_C_381, COMP_LOOP_C_382, COMP_LOOP_C_383, COMP_LOOP_C_384,
      COMP_LOOP_C_385, COMP_LOOP_C_386, COMP_LOOP_C_387, COMP_LOOP_C_388, COMP_LOOP_C_389,
      COMP_LOOP_C_390, COMP_LOOP_C_391, COMP_LOOP_C_392, COMP_LOOP_C_393, COMP_LOOP_C_394,
      COMP_LOOP_C_395, COMP_LOOP_C_396, COMP_LOOP_C_397, COMP_LOOP_C_398, COMP_LOOP_C_399,
      COMP_LOOP_C_400, COMP_LOOP_C_401, COMP_LOOP_C_402, COMP_LOOP_C_403, COMP_LOOP_C_404,
      COMP_LOOP_C_405, COMP_LOOP_C_406, COMP_LOOP_C_407, COMP_LOOP_C_408, COMP_LOOP_C_409,
      COMP_LOOP_C_410, COMP_LOOP_C_411, COMP_LOOP_C_412, COMP_LOOP_C_413, COMP_LOOP_C_414,
      COMP_LOOP_C_415, COMP_LOOP_C_416, COMP_LOOP_C_417, COMP_LOOP_C_418, COMP_LOOP_C_419,
      COMP_LOOP_C_420, COMP_LOOP_C_421, COMP_LOOP_C_422, COMP_LOOP_C_423, COMP_LOOP_C_424,
      COMP_LOOP_C_425, COMP_LOOP_C_426, COMP_LOOP_C_427, COMP_LOOP_C_428, COMP_LOOP_C_429,
      COMP_LOOP_C_430, COMP_LOOP_C_431, COMP_LOOP_C_432, COMP_LOOP_C_433, COMP_LOOP_C_434,
      COMP_LOOP_C_435, COMP_LOOP_8_modExp_1_while_C_0, COMP_LOOP_8_modExp_1_while_C_1,
      COMP_LOOP_8_modExp_1_while_C_2, COMP_LOOP_8_modExp_1_while_C_3, COMP_LOOP_8_modExp_1_while_C_4,
      COMP_LOOP_8_modExp_1_while_C_5, COMP_LOOP_8_modExp_1_while_C_6, COMP_LOOP_8_modExp_1_while_C_7,
      COMP_LOOP_8_modExp_1_while_C_8, COMP_LOOP_8_modExp_1_while_C_9, COMP_LOOP_8_modExp_1_while_C_10,
      COMP_LOOP_8_modExp_1_while_C_11, COMP_LOOP_8_modExp_1_while_C_12, COMP_LOOP_8_modExp_1_while_C_13,
      COMP_LOOP_8_modExp_1_while_C_14, COMP_LOOP_8_modExp_1_while_C_15, COMP_LOOP_8_modExp_1_while_C_16,
      COMP_LOOP_8_modExp_1_while_C_17, COMP_LOOP_8_modExp_1_while_C_18, COMP_LOOP_8_modExp_1_while_C_19,
      COMP_LOOP_8_modExp_1_while_C_20, COMP_LOOP_8_modExp_1_while_C_21, COMP_LOOP_8_modExp_1_while_C_22,
      COMP_LOOP_8_modExp_1_while_C_23, COMP_LOOP_8_modExp_1_while_C_24, COMP_LOOP_8_modExp_1_while_C_25,
      COMP_LOOP_8_modExp_1_while_C_26, COMP_LOOP_8_modExp_1_while_C_27, COMP_LOOP_8_modExp_1_while_C_28,
      COMP_LOOP_8_modExp_1_while_C_29, COMP_LOOP_8_modExp_1_while_C_30, COMP_LOOP_8_modExp_1_while_C_31,
      COMP_LOOP_8_modExp_1_while_C_32, COMP_LOOP_8_modExp_1_while_C_33, COMP_LOOP_8_modExp_1_while_C_34,
      COMP_LOOP_8_modExp_1_while_C_35, COMP_LOOP_8_modExp_1_while_C_36, COMP_LOOP_8_modExp_1_while_C_37,
      COMP_LOOP_8_modExp_1_while_C_38, COMP_LOOP_C_436, COMP_LOOP_C_437, COMP_LOOP_C_438,
      COMP_LOOP_C_439, COMP_LOOP_C_440, COMP_LOOP_C_441, COMP_LOOP_C_442, COMP_LOOP_C_443,
      COMP_LOOP_C_444, COMP_LOOP_C_445, COMP_LOOP_C_446, COMP_LOOP_C_447, COMP_LOOP_C_448,
      COMP_LOOP_C_449, COMP_LOOP_C_450, COMP_LOOP_C_451, COMP_LOOP_C_452, COMP_LOOP_C_453,
      COMP_LOOP_C_454, COMP_LOOP_C_455, COMP_LOOP_C_456, COMP_LOOP_C_457, COMP_LOOP_C_458,
      COMP_LOOP_C_459, COMP_LOOP_C_460, COMP_LOOP_C_461, COMP_LOOP_C_462, COMP_LOOP_C_463,
      COMP_LOOP_C_464, COMP_LOOP_C_465, COMP_LOOP_C_466, COMP_LOOP_C_467, COMP_LOOP_C_468,
      COMP_LOOP_C_469, COMP_LOOP_C_470, COMP_LOOP_C_471, COMP_LOOP_C_472, COMP_LOOP_C_473,
      COMP_LOOP_C_474, COMP_LOOP_C_475, COMP_LOOP_C_476, COMP_LOOP_C_477, COMP_LOOP_C_478,
      COMP_LOOP_C_479, COMP_LOOP_C_480, COMP_LOOP_C_481, COMP_LOOP_C_482, COMP_LOOP_C_483,
      COMP_LOOP_C_484, COMP_LOOP_C_485, COMP_LOOP_C_486, COMP_LOOP_C_487, COMP_LOOP_C_488,
      COMP_LOOP_C_489, COMP_LOOP_C_490, COMP_LOOP_C_491, COMP_LOOP_C_492, COMP_LOOP_C_493,
      COMP_LOOP_C_494, COMP_LOOP_C_495, COMP_LOOP_C_496, COMP_LOOP_C_497, COMP_LOOP_9_modExp_1_while_C_0,
      COMP_LOOP_9_modExp_1_while_C_1, COMP_LOOP_9_modExp_1_while_C_2, COMP_LOOP_9_modExp_1_while_C_3,
      COMP_LOOP_9_modExp_1_while_C_4, COMP_LOOP_9_modExp_1_while_C_5, COMP_LOOP_9_modExp_1_while_C_6,
      COMP_LOOP_9_modExp_1_while_C_7, COMP_LOOP_9_modExp_1_while_C_8, COMP_LOOP_9_modExp_1_while_C_9,
      COMP_LOOP_9_modExp_1_while_C_10, COMP_LOOP_9_modExp_1_while_C_11, COMP_LOOP_9_modExp_1_while_C_12,
      COMP_LOOP_9_modExp_1_while_C_13, COMP_LOOP_9_modExp_1_while_C_14, COMP_LOOP_9_modExp_1_while_C_15,
      COMP_LOOP_9_modExp_1_while_C_16, COMP_LOOP_9_modExp_1_while_C_17, COMP_LOOP_9_modExp_1_while_C_18,
      COMP_LOOP_9_modExp_1_while_C_19, COMP_LOOP_9_modExp_1_while_C_20, COMP_LOOP_9_modExp_1_while_C_21,
      COMP_LOOP_9_modExp_1_while_C_22, COMP_LOOP_9_modExp_1_while_C_23, COMP_LOOP_9_modExp_1_while_C_24,
      COMP_LOOP_9_modExp_1_while_C_25, COMP_LOOP_9_modExp_1_while_C_26, COMP_LOOP_9_modExp_1_while_C_27,
      COMP_LOOP_9_modExp_1_while_C_28, COMP_LOOP_9_modExp_1_while_C_29, COMP_LOOP_9_modExp_1_while_C_30,
      COMP_LOOP_9_modExp_1_while_C_31, COMP_LOOP_9_modExp_1_while_C_32, COMP_LOOP_9_modExp_1_while_C_33,
      COMP_LOOP_9_modExp_1_while_C_34, COMP_LOOP_9_modExp_1_while_C_35, COMP_LOOP_9_modExp_1_while_C_36,
      COMP_LOOP_9_modExp_1_while_C_37, COMP_LOOP_9_modExp_1_while_C_38, COMP_LOOP_C_498,
      COMP_LOOP_C_499, COMP_LOOP_C_500, COMP_LOOP_C_501, COMP_LOOP_C_502, COMP_LOOP_C_503,
      COMP_LOOP_C_504, COMP_LOOP_C_505, COMP_LOOP_C_506, COMP_LOOP_C_507, COMP_LOOP_C_508,
      COMP_LOOP_C_509, COMP_LOOP_C_510, COMP_LOOP_C_511, COMP_LOOP_C_512, COMP_LOOP_C_513,
      COMP_LOOP_C_514, COMP_LOOP_C_515, COMP_LOOP_C_516, COMP_LOOP_C_517, COMP_LOOP_C_518,
      COMP_LOOP_C_519, COMP_LOOP_C_520, COMP_LOOP_C_521, COMP_LOOP_C_522, COMP_LOOP_C_523,
      COMP_LOOP_C_524, COMP_LOOP_C_525, COMP_LOOP_C_526, COMP_LOOP_C_527, COMP_LOOP_C_528,
      COMP_LOOP_C_529, COMP_LOOP_C_530, COMP_LOOP_C_531, COMP_LOOP_C_532, COMP_LOOP_C_533,
      COMP_LOOP_C_534, COMP_LOOP_C_535, COMP_LOOP_C_536, COMP_LOOP_C_537, COMP_LOOP_C_538,
      COMP_LOOP_C_539, COMP_LOOP_C_540, COMP_LOOP_C_541, COMP_LOOP_C_542, COMP_LOOP_C_543,
      COMP_LOOP_C_544, COMP_LOOP_C_545, COMP_LOOP_C_546, COMP_LOOP_C_547, COMP_LOOP_C_548,
      COMP_LOOP_C_549, COMP_LOOP_C_550, COMP_LOOP_C_551, COMP_LOOP_C_552, COMP_LOOP_C_553,
      COMP_LOOP_C_554, COMP_LOOP_C_555, COMP_LOOP_C_556, COMP_LOOP_C_557, COMP_LOOP_C_558,
      COMP_LOOP_C_559, COMP_LOOP_10_modExp_1_while_C_0, COMP_LOOP_10_modExp_1_while_C_1,
      COMP_LOOP_10_modExp_1_while_C_2, COMP_LOOP_10_modExp_1_while_C_3, COMP_LOOP_10_modExp_1_while_C_4,
      COMP_LOOP_10_modExp_1_while_C_5, COMP_LOOP_10_modExp_1_while_C_6, COMP_LOOP_10_modExp_1_while_C_7,
      COMP_LOOP_10_modExp_1_while_C_8, COMP_LOOP_10_modExp_1_while_C_9, COMP_LOOP_10_modExp_1_while_C_10,
      COMP_LOOP_10_modExp_1_while_C_11, COMP_LOOP_10_modExp_1_while_C_12, COMP_LOOP_10_modExp_1_while_C_13,
      COMP_LOOP_10_modExp_1_while_C_14, COMP_LOOP_10_modExp_1_while_C_15, COMP_LOOP_10_modExp_1_while_C_16,
      COMP_LOOP_10_modExp_1_while_C_17, COMP_LOOP_10_modExp_1_while_C_18, COMP_LOOP_10_modExp_1_while_C_19,
      COMP_LOOP_10_modExp_1_while_C_20, COMP_LOOP_10_modExp_1_while_C_21, COMP_LOOP_10_modExp_1_while_C_22,
      COMP_LOOP_10_modExp_1_while_C_23, COMP_LOOP_10_modExp_1_while_C_24, COMP_LOOP_10_modExp_1_while_C_25,
      COMP_LOOP_10_modExp_1_while_C_26, COMP_LOOP_10_modExp_1_while_C_27, COMP_LOOP_10_modExp_1_while_C_28,
      COMP_LOOP_10_modExp_1_while_C_29, COMP_LOOP_10_modExp_1_while_C_30, COMP_LOOP_10_modExp_1_while_C_31,
      COMP_LOOP_10_modExp_1_while_C_32, COMP_LOOP_10_modExp_1_while_C_33, COMP_LOOP_10_modExp_1_while_C_34,
      COMP_LOOP_10_modExp_1_while_C_35, COMP_LOOP_10_modExp_1_while_C_36, COMP_LOOP_10_modExp_1_while_C_37,
      COMP_LOOP_10_modExp_1_while_C_38, COMP_LOOP_C_560, COMP_LOOP_C_561, COMP_LOOP_C_562,
      COMP_LOOP_C_563, COMP_LOOP_C_564, COMP_LOOP_C_565, COMP_LOOP_C_566, COMP_LOOP_C_567,
      COMP_LOOP_C_568, COMP_LOOP_C_569, COMP_LOOP_C_570, COMP_LOOP_C_571, COMP_LOOP_C_572,
      COMP_LOOP_C_573, COMP_LOOP_C_574, COMP_LOOP_C_575, COMP_LOOP_C_576, COMP_LOOP_C_577,
      COMP_LOOP_C_578, COMP_LOOP_C_579, COMP_LOOP_C_580, COMP_LOOP_C_581, COMP_LOOP_C_582,
      COMP_LOOP_C_583, COMP_LOOP_C_584, COMP_LOOP_C_585, COMP_LOOP_C_586, COMP_LOOP_C_587,
      COMP_LOOP_C_588, COMP_LOOP_C_589, COMP_LOOP_C_590, COMP_LOOP_C_591, COMP_LOOP_C_592,
      COMP_LOOP_C_593, COMP_LOOP_C_594, COMP_LOOP_C_595, COMP_LOOP_C_596, COMP_LOOP_C_597,
      COMP_LOOP_C_598, COMP_LOOP_C_599, COMP_LOOP_C_600, COMP_LOOP_C_601, COMP_LOOP_C_602,
      COMP_LOOP_C_603, COMP_LOOP_C_604, COMP_LOOP_C_605, COMP_LOOP_C_606, COMP_LOOP_C_607,
      COMP_LOOP_C_608, COMP_LOOP_C_609, COMP_LOOP_C_610, COMP_LOOP_C_611, COMP_LOOP_C_612,
      COMP_LOOP_C_613, COMP_LOOP_C_614, COMP_LOOP_C_615, COMP_LOOP_C_616, COMP_LOOP_C_617,
      COMP_LOOP_C_618, COMP_LOOP_C_619, COMP_LOOP_C_620, COMP_LOOP_C_621, COMP_LOOP_11_modExp_1_while_C_0,
      COMP_LOOP_11_modExp_1_while_C_1, COMP_LOOP_11_modExp_1_while_C_2, COMP_LOOP_11_modExp_1_while_C_3,
      COMP_LOOP_11_modExp_1_while_C_4, COMP_LOOP_11_modExp_1_while_C_5, COMP_LOOP_11_modExp_1_while_C_6,
      COMP_LOOP_11_modExp_1_while_C_7, COMP_LOOP_11_modExp_1_while_C_8, COMP_LOOP_11_modExp_1_while_C_9,
      COMP_LOOP_11_modExp_1_while_C_10, COMP_LOOP_11_modExp_1_while_C_11, COMP_LOOP_11_modExp_1_while_C_12,
      COMP_LOOP_11_modExp_1_while_C_13, COMP_LOOP_11_modExp_1_while_C_14, COMP_LOOP_11_modExp_1_while_C_15,
      COMP_LOOP_11_modExp_1_while_C_16, COMP_LOOP_11_modExp_1_while_C_17, COMP_LOOP_11_modExp_1_while_C_18,
      COMP_LOOP_11_modExp_1_while_C_19, COMP_LOOP_11_modExp_1_while_C_20, COMP_LOOP_11_modExp_1_while_C_21,
      COMP_LOOP_11_modExp_1_while_C_22, COMP_LOOP_11_modExp_1_while_C_23, COMP_LOOP_11_modExp_1_while_C_24,
      COMP_LOOP_11_modExp_1_while_C_25, COMP_LOOP_11_modExp_1_while_C_26, COMP_LOOP_11_modExp_1_while_C_27,
      COMP_LOOP_11_modExp_1_while_C_28, COMP_LOOP_11_modExp_1_while_C_29, COMP_LOOP_11_modExp_1_while_C_30,
      COMP_LOOP_11_modExp_1_while_C_31, COMP_LOOP_11_modExp_1_while_C_32, COMP_LOOP_11_modExp_1_while_C_33,
      COMP_LOOP_11_modExp_1_while_C_34, COMP_LOOP_11_modExp_1_while_C_35, COMP_LOOP_11_modExp_1_while_C_36,
      COMP_LOOP_11_modExp_1_while_C_37, COMP_LOOP_11_modExp_1_while_C_38, COMP_LOOP_C_622,
      COMP_LOOP_C_623, COMP_LOOP_C_624, COMP_LOOP_C_625, COMP_LOOP_C_626, COMP_LOOP_C_627,
      COMP_LOOP_C_628, COMP_LOOP_C_629, COMP_LOOP_C_630, COMP_LOOP_C_631, COMP_LOOP_C_632,
      COMP_LOOP_C_633, COMP_LOOP_C_634, COMP_LOOP_C_635, COMP_LOOP_C_636, COMP_LOOP_C_637,
      COMP_LOOP_C_638, COMP_LOOP_C_639, COMP_LOOP_C_640, COMP_LOOP_C_641, COMP_LOOP_C_642,
      COMP_LOOP_C_643, COMP_LOOP_C_644, COMP_LOOP_C_645, COMP_LOOP_C_646, COMP_LOOP_C_647,
      COMP_LOOP_C_648, COMP_LOOP_C_649, COMP_LOOP_C_650, COMP_LOOP_C_651, COMP_LOOP_C_652,
      COMP_LOOP_C_653, COMP_LOOP_C_654, COMP_LOOP_C_655, COMP_LOOP_C_656, COMP_LOOP_C_657,
      COMP_LOOP_C_658, COMP_LOOP_C_659, COMP_LOOP_C_660, COMP_LOOP_C_661, COMP_LOOP_C_662,
      COMP_LOOP_C_663, COMP_LOOP_C_664, COMP_LOOP_C_665, COMP_LOOP_C_666, COMP_LOOP_C_667,
      COMP_LOOP_C_668, COMP_LOOP_C_669, COMP_LOOP_C_670, COMP_LOOP_C_671, COMP_LOOP_C_672,
      COMP_LOOP_C_673, COMP_LOOP_C_674, COMP_LOOP_C_675, COMP_LOOP_C_676, COMP_LOOP_C_677,
      COMP_LOOP_C_678, COMP_LOOP_C_679, COMP_LOOP_C_680, COMP_LOOP_C_681, COMP_LOOP_C_682,
      COMP_LOOP_C_683, COMP_LOOP_12_modExp_1_while_C_0, COMP_LOOP_12_modExp_1_while_C_1,
      COMP_LOOP_12_modExp_1_while_C_2, COMP_LOOP_12_modExp_1_while_C_3, COMP_LOOP_12_modExp_1_while_C_4,
      COMP_LOOP_12_modExp_1_while_C_5, COMP_LOOP_12_modExp_1_while_C_6, COMP_LOOP_12_modExp_1_while_C_7,
      COMP_LOOP_12_modExp_1_while_C_8, COMP_LOOP_12_modExp_1_while_C_9, COMP_LOOP_12_modExp_1_while_C_10,
      COMP_LOOP_12_modExp_1_while_C_11, COMP_LOOP_12_modExp_1_while_C_12, COMP_LOOP_12_modExp_1_while_C_13,
      COMP_LOOP_12_modExp_1_while_C_14, COMP_LOOP_12_modExp_1_while_C_15, COMP_LOOP_12_modExp_1_while_C_16,
      COMP_LOOP_12_modExp_1_while_C_17, COMP_LOOP_12_modExp_1_while_C_18, COMP_LOOP_12_modExp_1_while_C_19,
      COMP_LOOP_12_modExp_1_while_C_20, COMP_LOOP_12_modExp_1_while_C_21, COMP_LOOP_12_modExp_1_while_C_22,
      COMP_LOOP_12_modExp_1_while_C_23, COMP_LOOP_12_modExp_1_while_C_24, COMP_LOOP_12_modExp_1_while_C_25,
      COMP_LOOP_12_modExp_1_while_C_26, COMP_LOOP_12_modExp_1_while_C_27, COMP_LOOP_12_modExp_1_while_C_28,
      COMP_LOOP_12_modExp_1_while_C_29, COMP_LOOP_12_modExp_1_while_C_30, COMP_LOOP_12_modExp_1_while_C_31,
      COMP_LOOP_12_modExp_1_while_C_32, COMP_LOOP_12_modExp_1_while_C_33, COMP_LOOP_12_modExp_1_while_C_34,
      COMP_LOOP_12_modExp_1_while_C_35, COMP_LOOP_12_modExp_1_while_C_36, COMP_LOOP_12_modExp_1_while_C_37,
      COMP_LOOP_12_modExp_1_while_C_38, COMP_LOOP_C_684, COMP_LOOP_C_685, COMP_LOOP_C_686,
      COMP_LOOP_C_687, COMP_LOOP_C_688, COMP_LOOP_C_689, COMP_LOOP_C_690, COMP_LOOP_C_691,
      COMP_LOOP_C_692, COMP_LOOP_C_693, COMP_LOOP_C_694, COMP_LOOP_C_695, COMP_LOOP_C_696,
      COMP_LOOP_C_697, COMP_LOOP_C_698, COMP_LOOP_C_699, COMP_LOOP_C_700, COMP_LOOP_C_701,
      COMP_LOOP_C_702, COMP_LOOP_C_703, COMP_LOOP_C_704, COMP_LOOP_C_705, COMP_LOOP_C_706,
      COMP_LOOP_C_707, COMP_LOOP_C_708, COMP_LOOP_C_709, COMP_LOOP_C_710, COMP_LOOP_C_711,
      COMP_LOOP_C_712, COMP_LOOP_C_713, COMP_LOOP_C_714, COMP_LOOP_C_715, COMP_LOOP_C_716,
      COMP_LOOP_C_717, COMP_LOOP_C_718, COMP_LOOP_C_719, COMP_LOOP_C_720, COMP_LOOP_C_721,
      COMP_LOOP_C_722, COMP_LOOP_C_723, COMP_LOOP_C_724, COMP_LOOP_C_725, COMP_LOOP_C_726,
      COMP_LOOP_C_727, COMP_LOOP_C_728, COMP_LOOP_C_729, COMP_LOOP_C_730, COMP_LOOP_C_731,
      COMP_LOOP_C_732, COMP_LOOP_C_733, COMP_LOOP_C_734, COMP_LOOP_C_735, COMP_LOOP_C_736,
      COMP_LOOP_C_737, COMP_LOOP_C_738, COMP_LOOP_C_739, COMP_LOOP_C_740, COMP_LOOP_C_741,
      COMP_LOOP_C_742, COMP_LOOP_C_743, COMP_LOOP_C_744, COMP_LOOP_C_745, COMP_LOOP_13_modExp_1_while_C_0,
      COMP_LOOP_13_modExp_1_while_C_1, COMP_LOOP_13_modExp_1_while_C_2, COMP_LOOP_13_modExp_1_while_C_3,
      COMP_LOOP_13_modExp_1_while_C_4, COMP_LOOP_13_modExp_1_while_C_5, COMP_LOOP_13_modExp_1_while_C_6,
      COMP_LOOP_13_modExp_1_while_C_7, COMP_LOOP_13_modExp_1_while_C_8, COMP_LOOP_13_modExp_1_while_C_9,
      COMP_LOOP_13_modExp_1_while_C_10, COMP_LOOP_13_modExp_1_while_C_11, COMP_LOOP_13_modExp_1_while_C_12,
      COMP_LOOP_13_modExp_1_while_C_13, COMP_LOOP_13_modExp_1_while_C_14, COMP_LOOP_13_modExp_1_while_C_15,
      COMP_LOOP_13_modExp_1_while_C_16, COMP_LOOP_13_modExp_1_while_C_17, COMP_LOOP_13_modExp_1_while_C_18,
      COMP_LOOP_13_modExp_1_while_C_19, COMP_LOOP_13_modExp_1_while_C_20, COMP_LOOP_13_modExp_1_while_C_21,
      COMP_LOOP_13_modExp_1_while_C_22, COMP_LOOP_13_modExp_1_while_C_23, COMP_LOOP_13_modExp_1_while_C_24,
      COMP_LOOP_13_modExp_1_while_C_25, COMP_LOOP_13_modExp_1_while_C_26, COMP_LOOP_13_modExp_1_while_C_27,
      COMP_LOOP_13_modExp_1_while_C_28, COMP_LOOP_13_modExp_1_while_C_29, COMP_LOOP_13_modExp_1_while_C_30,
      COMP_LOOP_13_modExp_1_while_C_31, COMP_LOOP_13_modExp_1_while_C_32, COMP_LOOP_13_modExp_1_while_C_33,
      COMP_LOOP_13_modExp_1_while_C_34, COMP_LOOP_13_modExp_1_while_C_35, COMP_LOOP_13_modExp_1_while_C_36,
      COMP_LOOP_13_modExp_1_while_C_37, COMP_LOOP_13_modExp_1_while_C_38, COMP_LOOP_C_746,
      COMP_LOOP_C_747, COMP_LOOP_C_748, COMP_LOOP_C_749, COMP_LOOP_C_750, COMP_LOOP_C_751,
      COMP_LOOP_C_752, COMP_LOOP_C_753, COMP_LOOP_C_754, COMP_LOOP_C_755, COMP_LOOP_C_756,
      COMP_LOOP_C_757, COMP_LOOP_C_758, COMP_LOOP_C_759, COMP_LOOP_C_760, COMP_LOOP_C_761,
      COMP_LOOP_C_762, COMP_LOOP_C_763, COMP_LOOP_C_764, COMP_LOOP_C_765, COMP_LOOP_C_766,
      COMP_LOOP_C_767, COMP_LOOP_C_768, COMP_LOOP_C_769, COMP_LOOP_C_770, COMP_LOOP_C_771,
      COMP_LOOP_C_772, COMP_LOOP_C_773, COMP_LOOP_C_774, COMP_LOOP_C_775, COMP_LOOP_C_776,
      COMP_LOOP_C_777, COMP_LOOP_C_778, COMP_LOOP_C_779, COMP_LOOP_C_780, COMP_LOOP_C_781,
      COMP_LOOP_C_782, COMP_LOOP_C_783, COMP_LOOP_C_784, COMP_LOOP_C_785, COMP_LOOP_C_786,
      COMP_LOOP_C_787, COMP_LOOP_C_788, COMP_LOOP_C_789, COMP_LOOP_C_790, COMP_LOOP_C_791,
      COMP_LOOP_C_792, COMP_LOOP_C_793, COMP_LOOP_C_794, COMP_LOOP_C_795, COMP_LOOP_C_796,
      COMP_LOOP_C_797, COMP_LOOP_C_798, COMP_LOOP_C_799, COMP_LOOP_C_800, COMP_LOOP_C_801,
      COMP_LOOP_C_802, COMP_LOOP_C_803, COMP_LOOP_C_804, COMP_LOOP_C_805, COMP_LOOP_C_806,
      COMP_LOOP_C_807, COMP_LOOP_14_modExp_1_while_C_0, COMP_LOOP_14_modExp_1_while_C_1,
      COMP_LOOP_14_modExp_1_while_C_2, COMP_LOOP_14_modExp_1_while_C_3, COMP_LOOP_14_modExp_1_while_C_4,
      COMP_LOOP_14_modExp_1_while_C_5, COMP_LOOP_14_modExp_1_while_C_6, COMP_LOOP_14_modExp_1_while_C_7,
      COMP_LOOP_14_modExp_1_while_C_8, COMP_LOOP_14_modExp_1_while_C_9, COMP_LOOP_14_modExp_1_while_C_10,
      COMP_LOOP_14_modExp_1_while_C_11, COMP_LOOP_14_modExp_1_while_C_12, COMP_LOOP_14_modExp_1_while_C_13,
      COMP_LOOP_14_modExp_1_while_C_14, COMP_LOOP_14_modExp_1_while_C_15, COMP_LOOP_14_modExp_1_while_C_16,
      COMP_LOOP_14_modExp_1_while_C_17, COMP_LOOP_14_modExp_1_while_C_18, COMP_LOOP_14_modExp_1_while_C_19,
      COMP_LOOP_14_modExp_1_while_C_20, COMP_LOOP_14_modExp_1_while_C_21, COMP_LOOP_14_modExp_1_while_C_22,
      COMP_LOOP_14_modExp_1_while_C_23, COMP_LOOP_14_modExp_1_while_C_24, COMP_LOOP_14_modExp_1_while_C_25,
      COMP_LOOP_14_modExp_1_while_C_26, COMP_LOOP_14_modExp_1_while_C_27, COMP_LOOP_14_modExp_1_while_C_28,
      COMP_LOOP_14_modExp_1_while_C_29, COMP_LOOP_14_modExp_1_while_C_30, COMP_LOOP_14_modExp_1_while_C_31,
      COMP_LOOP_14_modExp_1_while_C_32, COMP_LOOP_14_modExp_1_while_C_33, COMP_LOOP_14_modExp_1_while_C_34,
      COMP_LOOP_14_modExp_1_while_C_35, COMP_LOOP_14_modExp_1_while_C_36, COMP_LOOP_14_modExp_1_while_C_37,
      COMP_LOOP_14_modExp_1_while_C_38, COMP_LOOP_C_808, COMP_LOOP_C_809, COMP_LOOP_C_810,
      COMP_LOOP_C_811, COMP_LOOP_C_812, COMP_LOOP_C_813, COMP_LOOP_C_814, COMP_LOOP_C_815,
      COMP_LOOP_C_816, COMP_LOOP_C_817, COMP_LOOP_C_818, COMP_LOOP_C_819, COMP_LOOP_C_820,
      COMP_LOOP_C_821, COMP_LOOP_C_822, COMP_LOOP_C_823, COMP_LOOP_C_824, COMP_LOOP_C_825,
      COMP_LOOP_C_826, COMP_LOOP_C_827, COMP_LOOP_C_828, COMP_LOOP_C_829, COMP_LOOP_C_830,
      COMP_LOOP_C_831, COMP_LOOP_C_832, COMP_LOOP_C_833, COMP_LOOP_C_834, COMP_LOOP_C_835,
      COMP_LOOP_C_836, COMP_LOOP_C_837, COMP_LOOP_C_838, COMP_LOOP_C_839, COMP_LOOP_C_840,
      COMP_LOOP_C_841, COMP_LOOP_C_842, COMP_LOOP_C_843, COMP_LOOP_C_844, COMP_LOOP_C_845,
      COMP_LOOP_C_846, COMP_LOOP_C_847, COMP_LOOP_C_848, COMP_LOOP_C_849, COMP_LOOP_C_850,
      COMP_LOOP_C_851, COMP_LOOP_C_852, COMP_LOOP_C_853, COMP_LOOP_C_854, COMP_LOOP_C_855,
      COMP_LOOP_C_856, COMP_LOOP_C_857, COMP_LOOP_C_858, COMP_LOOP_C_859, COMP_LOOP_C_860,
      COMP_LOOP_C_861, COMP_LOOP_C_862, COMP_LOOP_C_863, COMP_LOOP_C_864, COMP_LOOP_C_865,
      COMP_LOOP_C_866, COMP_LOOP_C_867, COMP_LOOP_C_868, COMP_LOOP_C_869, COMP_LOOP_15_modExp_1_while_C_0,
      COMP_LOOP_15_modExp_1_while_C_1, COMP_LOOP_15_modExp_1_while_C_2, COMP_LOOP_15_modExp_1_while_C_3,
      COMP_LOOP_15_modExp_1_while_C_4, COMP_LOOP_15_modExp_1_while_C_5, COMP_LOOP_15_modExp_1_while_C_6,
      COMP_LOOP_15_modExp_1_while_C_7, COMP_LOOP_15_modExp_1_while_C_8, COMP_LOOP_15_modExp_1_while_C_9,
      COMP_LOOP_15_modExp_1_while_C_10, COMP_LOOP_15_modExp_1_while_C_11, COMP_LOOP_15_modExp_1_while_C_12,
      COMP_LOOP_15_modExp_1_while_C_13, COMP_LOOP_15_modExp_1_while_C_14, COMP_LOOP_15_modExp_1_while_C_15,
      COMP_LOOP_15_modExp_1_while_C_16, COMP_LOOP_15_modExp_1_while_C_17, COMP_LOOP_15_modExp_1_while_C_18,
      COMP_LOOP_15_modExp_1_while_C_19, COMP_LOOP_15_modExp_1_while_C_20, COMP_LOOP_15_modExp_1_while_C_21,
      COMP_LOOP_15_modExp_1_while_C_22, COMP_LOOP_15_modExp_1_while_C_23, COMP_LOOP_15_modExp_1_while_C_24,
      COMP_LOOP_15_modExp_1_while_C_25, COMP_LOOP_15_modExp_1_while_C_26, COMP_LOOP_15_modExp_1_while_C_27,
      COMP_LOOP_15_modExp_1_while_C_28, COMP_LOOP_15_modExp_1_while_C_29, COMP_LOOP_15_modExp_1_while_C_30,
      COMP_LOOP_15_modExp_1_while_C_31, COMP_LOOP_15_modExp_1_while_C_32, COMP_LOOP_15_modExp_1_while_C_33,
      COMP_LOOP_15_modExp_1_while_C_34, COMP_LOOP_15_modExp_1_while_C_35, COMP_LOOP_15_modExp_1_while_C_36,
      COMP_LOOP_15_modExp_1_while_C_37, COMP_LOOP_15_modExp_1_while_C_38, COMP_LOOP_C_870,
      COMP_LOOP_C_871, COMP_LOOP_C_872, COMP_LOOP_C_873, COMP_LOOP_C_874, COMP_LOOP_C_875,
      COMP_LOOP_C_876, COMP_LOOP_C_877, COMP_LOOP_C_878, COMP_LOOP_C_879, COMP_LOOP_C_880,
      COMP_LOOP_C_881, COMP_LOOP_C_882, COMP_LOOP_C_883, COMP_LOOP_C_884, COMP_LOOP_C_885,
      COMP_LOOP_C_886, COMP_LOOP_C_887, COMP_LOOP_C_888, COMP_LOOP_C_889, COMP_LOOP_C_890,
      COMP_LOOP_C_891, COMP_LOOP_C_892, COMP_LOOP_C_893, COMP_LOOP_C_894, COMP_LOOP_C_895,
      COMP_LOOP_C_896, COMP_LOOP_C_897, COMP_LOOP_C_898, COMP_LOOP_C_899, COMP_LOOP_C_900,
      COMP_LOOP_C_901, COMP_LOOP_C_902, COMP_LOOP_C_903, COMP_LOOP_C_904, COMP_LOOP_C_905,
      COMP_LOOP_C_906, COMP_LOOP_C_907, COMP_LOOP_C_908, COMP_LOOP_C_909, COMP_LOOP_C_910,
      COMP_LOOP_C_911, COMP_LOOP_C_912, COMP_LOOP_C_913, COMP_LOOP_C_914, COMP_LOOP_C_915,
      COMP_LOOP_C_916, COMP_LOOP_C_917, COMP_LOOP_C_918, COMP_LOOP_C_919, COMP_LOOP_C_920,
      COMP_LOOP_C_921, COMP_LOOP_C_922, COMP_LOOP_C_923, COMP_LOOP_C_924, COMP_LOOP_C_925,
      COMP_LOOP_C_926, COMP_LOOP_C_927, COMP_LOOP_C_928, COMP_LOOP_C_929, COMP_LOOP_C_930,
      COMP_LOOP_C_931, COMP_LOOP_16_modExp_1_while_C_0, COMP_LOOP_16_modExp_1_while_C_1,
      COMP_LOOP_16_modExp_1_while_C_2, COMP_LOOP_16_modExp_1_while_C_3, COMP_LOOP_16_modExp_1_while_C_4,
      COMP_LOOP_16_modExp_1_while_C_5, COMP_LOOP_16_modExp_1_while_C_6, COMP_LOOP_16_modExp_1_while_C_7,
      COMP_LOOP_16_modExp_1_while_C_8, COMP_LOOP_16_modExp_1_while_C_9, COMP_LOOP_16_modExp_1_while_C_10,
      COMP_LOOP_16_modExp_1_while_C_11, COMP_LOOP_16_modExp_1_while_C_12, COMP_LOOP_16_modExp_1_while_C_13,
      COMP_LOOP_16_modExp_1_while_C_14, COMP_LOOP_16_modExp_1_while_C_15, COMP_LOOP_16_modExp_1_while_C_16,
      COMP_LOOP_16_modExp_1_while_C_17, COMP_LOOP_16_modExp_1_while_C_18, COMP_LOOP_16_modExp_1_while_C_19,
      COMP_LOOP_16_modExp_1_while_C_20, COMP_LOOP_16_modExp_1_while_C_21, COMP_LOOP_16_modExp_1_while_C_22,
      COMP_LOOP_16_modExp_1_while_C_23, COMP_LOOP_16_modExp_1_while_C_24, COMP_LOOP_16_modExp_1_while_C_25,
      COMP_LOOP_16_modExp_1_while_C_26, COMP_LOOP_16_modExp_1_while_C_27, COMP_LOOP_16_modExp_1_while_C_28,
      COMP_LOOP_16_modExp_1_while_C_29, COMP_LOOP_16_modExp_1_while_C_30, COMP_LOOP_16_modExp_1_while_C_31,
      COMP_LOOP_16_modExp_1_while_C_32, COMP_LOOP_16_modExp_1_while_C_33, COMP_LOOP_16_modExp_1_while_C_34,
      COMP_LOOP_16_modExp_1_while_C_35, COMP_LOOP_16_modExp_1_while_C_36, COMP_LOOP_16_modExp_1_while_C_37,
      COMP_LOOP_16_modExp_1_while_C_38, COMP_LOOP_C_932, COMP_LOOP_C_933, COMP_LOOP_C_934,
      COMP_LOOP_C_935, COMP_LOOP_C_936, COMP_LOOP_C_937, COMP_LOOP_C_938, COMP_LOOP_C_939,
      COMP_LOOP_C_940, COMP_LOOP_C_941, COMP_LOOP_C_942, COMP_LOOP_C_943, COMP_LOOP_C_944,
      COMP_LOOP_C_945, COMP_LOOP_C_946, COMP_LOOP_C_947, COMP_LOOP_C_948, COMP_LOOP_C_949,
      COMP_LOOP_C_950, COMP_LOOP_C_951, COMP_LOOP_C_952, COMP_LOOP_C_953, COMP_LOOP_C_954,
      COMP_LOOP_C_955, COMP_LOOP_C_956, COMP_LOOP_C_957, COMP_LOOP_C_958, COMP_LOOP_C_959,
      COMP_LOOP_C_960, COMP_LOOP_C_961, COMP_LOOP_C_962, COMP_LOOP_C_963, COMP_LOOP_C_964,
      COMP_LOOP_C_965, COMP_LOOP_C_966, COMP_LOOP_C_967, COMP_LOOP_C_968, COMP_LOOP_C_969,
      COMP_LOOP_C_970, COMP_LOOP_C_971, COMP_LOOP_C_972, COMP_LOOP_C_973, COMP_LOOP_C_974,
      COMP_LOOP_C_975, COMP_LOOP_C_976, COMP_LOOP_C_977, COMP_LOOP_C_978, COMP_LOOP_C_979,
      COMP_LOOP_C_980, COMP_LOOP_C_981, COMP_LOOP_C_982, COMP_LOOP_C_983, COMP_LOOP_C_984,
      COMP_LOOP_C_985, COMP_LOOP_C_986, COMP_LOOP_C_987, COMP_LOOP_C_988, COMP_LOOP_C_989,
      COMP_LOOP_C_990, COMP_LOOP_C_991, COMP_LOOP_C_992, VEC_LOOP_C_0, STAGE_LOOP_C_9,
      main_C_1);

  SIGNAL state_var : inPlaceNTT_DIT_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIT_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIT_core_core_fsm_1 : PROCESS (STAGE_LOOP_C_8_tr0, modExp_while_C_38_tr0,
      COMP_LOOP_C_1_tr0, COMP_LOOP_1_modExp_1_while_C_38_tr0, COMP_LOOP_C_62_tr0,
      COMP_LOOP_2_modExp_1_while_C_38_tr0, COMP_LOOP_C_124_tr0, COMP_LOOP_3_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_186_tr0, COMP_LOOP_4_modExp_1_while_C_38_tr0, COMP_LOOP_C_248_tr0,
      COMP_LOOP_5_modExp_1_while_C_38_tr0, COMP_LOOP_C_310_tr0, COMP_LOOP_6_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_372_tr0, COMP_LOOP_7_modExp_1_while_C_38_tr0, COMP_LOOP_C_434_tr0,
      COMP_LOOP_8_modExp_1_while_C_38_tr0, COMP_LOOP_C_496_tr0, COMP_LOOP_9_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_558_tr0, COMP_LOOP_10_modExp_1_while_C_38_tr0, COMP_LOOP_C_620_tr0,
      COMP_LOOP_11_modExp_1_while_C_38_tr0, COMP_LOOP_C_682_tr0, COMP_LOOP_12_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_744_tr0, COMP_LOOP_13_modExp_1_while_C_38_tr0, COMP_LOOP_C_806_tr0,
      COMP_LOOP_14_modExp_1_while_C_38_tr0, COMP_LOOP_C_868_tr0, COMP_LOOP_15_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_930_tr0, COMP_LOOP_16_modExp_1_while_C_38_tr0, COMP_LOOP_C_992_tr0,
      VEC_LOOP_C_0_tr0, STAGE_LOOP_C_9_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000001");
        state_var_NS <= STAGE_LOOP_C_1;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000010");
        state_var_NS <= STAGE_LOOP_C_2;
      WHEN STAGE_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000011");
        state_var_NS <= STAGE_LOOP_C_3;
      WHEN STAGE_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000100");
        state_var_NS <= STAGE_LOOP_C_4;
      WHEN STAGE_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000101");
        state_var_NS <= STAGE_LOOP_C_5;
      WHEN STAGE_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000110");
        state_var_NS <= STAGE_LOOP_C_6;
      WHEN STAGE_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000111");
        state_var_NS <= STAGE_LOOP_C_7;
      WHEN STAGE_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001000");
        state_var_NS <= STAGE_LOOP_C_8;
      WHEN STAGE_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001001");
        IF ( STAGE_LOOP_C_8_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_while_C_0;
        END IF;
      WHEN modExp_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001010");
        state_var_NS <= modExp_while_C_1;
      WHEN modExp_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001011");
        state_var_NS <= modExp_while_C_2;
      WHEN modExp_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001100");
        state_var_NS <= modExp_while_C_3;
      WHEN modExp_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001101");
        state_var_NS <= modExp_while_C_4;
      WHEN modExp_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001110");
        state_var_NS <= modExp_while_C_5;
      WHEN modExp_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001111");
        state_var_NS <= modExp_while_C_6;
      WHEN modExp_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010000");
        state_var_NS <= modExp_while_C_7;
      WHEN modExp_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010001");
        state_var_NS <= modExp_while_C_8;
      WHEN modExp_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010010");
        state_var_NS <= modExp_while_C_9;
      WHEN modExp_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010011");
        state_var_NS <= modExp_while_C_10;
      WHEN modExp_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010100");
        state_var_NS <= modExp_while_C_11;
      WHEN modExp_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010101");
        state_var_NS <= modExp_while_C_12;
      WHEN modExp_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010110");
        state_var_NS <= modExp_while_C_13;
      WHEN modExp_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010111");
        state_var_NS <= modExp_while_C_14;
      WHEN modExp_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011000");
        state_var_NS <= modExp_while_C_15;
      WHEN modExp_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011001");
        state_var_NS <= modExp_while_C_16;
      WHEN modExp_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011010");
        state_var_NS <= modExp_while_C_17;
      WHEN modExp_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011011");
        state_var_NS <= modExp_while_C_18;
      WHEN modExp_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011100");
        state_var_NS <= modExp_while_C_19;
      WHEN modExp_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011101");
        state_var_NS <= modExp_while_C_20;
      WHEN modExp_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011110");
        state_var_NS <= modExp_while_C_21;
      WHEN modExp_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011111");
        state_var_NS <= modExp_while_C_22;
      WHEN modExp_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100000");
        state_var_NS <= modExp_while_C_23;
      WHEN modExp_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100001");
        state_var_NS <= modExp_while_C_24;
      WHEN modExp_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100010");
        state_var_NS <= modExp_while_C_25;
      WHEN modExp_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100011");
        state_var_NS <= modExp_while_C_26;
      WHEN modExp_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100100");
        state_var_NS <= modExp_while_C_27;
      WHEN modExp_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100101");
        state_var_NS <= modExp_while_C_28;
      WHEN modExp_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100110");
        state_var_NS <= modExp_while_C_29;
      WHEN modExp_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100111");
        state_var_NS <= modExp_while_C_30;
      WHEN modExp_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101000");
        state_var_NS <= modExp_while_C_31;
      WHEN modExp_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101001");
        state_var_NS <= modExp_while_C_32;
      WHEN modExp_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101010");
        state_var_NS <= modExp_while_C_33;
      WHEN modExp_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101011");
        state_var_NS <= modExp_while_C_34;
      WHEN modExp_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101100");
        state_var_NS <= modExp_while_C_35;
      WHEN modExp_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101101");
        state_var_NS <= modExp_while_C_36;
      WHEN modExp_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101110");
        state_var_NS <= modExp_while_C_37;
      WHEN modExp_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101111");
        state_var_NS <= modExp_while_C_38;
      WHEN modExp_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110000");
        IF ( modExp_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110001");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110010");
        IF ( COMP_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_2;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_1_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_1;
      WHEN COMP_LOOP_1_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_2;
      WHEN COMP_LOOP_1_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_3;
      WHEN COMP_LOOP_1_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_4;
      WHEN COMP_LOOP_1_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_5;
      WHEN COMP_LOOP_1_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_6;
      WHEN COMP_LOOP_1_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_7;
      WHEN COMP_LOOP_1_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_8;
      WHEN COMP_LOOP_1_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_9;
      WHEN COMP_LOOP_1_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_10;
      WHEN COMP_LOOP_1_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_11;
      WHEN COMP_LOOP_1_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_12;
      WHEN COMP_LOOP_1_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_13;
      WHEN COMP_LOOP_1_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_14;
      WHEN COMP_LOOP_1_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_15;
      WHEN COMP_LOOP_1_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_16;
      WHEN COMP_LOOP_1_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_17;
      WHEN COMP_LOOP_1_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_18;
      WHEN COMP_LOOP_1_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_19;
      WHEN COMP_LOOP_1_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_20;
      WHEN COMP_LOOP_1_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_21;
      WHEN COMP_LOOP_1_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_22;
      WHEN COMP_LOOP_1_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_23;
      WHEN COMP_LOOP_1_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_24;
      WHEN COMP_LOOP_1_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_25;
      WHEN COMP_LOOP_1_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_26;
      WHEN COMP_LOOP_1_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_27;
      WHEN COMP_LOOP_1_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_28;
      WHEN COMP_LOOP_1_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_29;
      WHEN COMP_LOOP_1_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_30;
      WHEN COMP_LOOP_1_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010001");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_31;
      WHEN COMP_LOOP_1_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010010");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_32;
      WHEN COMP_LOOP_1_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010011");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_33;
      WHEN COMP_LOOP_1_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010100");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_34;
      WHEN COMP_LOOP_1_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010101");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_35;
      WHEN COMP_LOOP_1_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010110");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_36;
      WHEN COMP_LOOP_1_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010111");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_37;
      WHEN COMP_LOOP_1_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011000");
        state_var_NS <= COMP_LOOP_1_modExp_1_while_C_38;
      WHEN COMP_LOOP_1_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011001");
        IF ( COMP_LOOP_1_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_2;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011010");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011011");
        state_var_NS <= COMP_LOOP_C_4;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011100");
        state_var_NS <= COMP_LOOP_C_5;
      WHEN COMP_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011101");
        state_var_NS <= COMP_LOOP_C_6;
      WHEN COMP_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011110");
        state_var_NS <= COMP_LOOP_C_7;
      WHEN COMP_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011111");
        state_var_NS <= COMP_LOOP_C_8;
      WHEN COMP_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100000");
        state_var_NS <= COMP_LOOP_C_9;
      WHEN COMP_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100001");
        state_var_NS <= COMP_LOOP_C_10;
      WHEN COMP_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100010");
        state_var_NS <= COMP_LOOP_C_11;
      WHEN COMP_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100011");
        state_var_NS <= COMP_LOOP_C_12;
      WHEN COMP_LOOP_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100100");
        state_var_NS <= COMP_LOOP_C_13;
      WHEN COMP_LOOP_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100101");
        state_var_NS <= COMP_LOOP_C_14;
      WHEN COMP_LOOP_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100110");
        state_var_NS <= COMP_LOOP_C_15;
      WHEN COMP_LOOP_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100111");
        state_var_NS <= COMP_LOOP_C_16;
      WHEN COMP_LOOP_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101000");
        state_var_NS <= COMP_LOOP_C_17;
      WHEN COMP_LOOP_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101001");
        state_var_NS <= COMP_LOOP_C_18;
      WHEN COMP_LOOP_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101010");
        state_var_NS <= COMP_LOOP_C_19;
      WHEN COMP_LOOP_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101011");
        state_var_NS <= COMP_LOOP_C_20;
      WHEN COMP_LOOP_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101100");
        state_var_NS <= COMP_LOOP_C_21;
      WHEN COMP_LOOP_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101101");
        state_var_NS <= COMP_LOOP_C_22;
      WHEN COMP_LOOP_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101110");
        state_var_NS <= COMP_LOOP_C_23;
      WHEN COMP_LOOP_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101111");
        state_var_NS <= COMP_LOOP_C_24;
      WHEN COMP_LOOP_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110000");
        state_var_NS <= COMP_LOOP_C_25;
      WHEN COMP_LOOP_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110001");
        state_var_NS <= COMP_LOOP_C_26;
      WHEN COMP_LOOP_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110010");
        state_var_NS <= COMP_LOOP_C_27;
      WHEN COMP_LOOP_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110011");
        state_var_NS <= COMP_LOOP_C_28;
      WHEN COMP_LOOP_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110100");
        state_var_NS <= COMP_LOOP_C_29;
      WHEN COMP_LOOP_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110101");
        state_var_NS <= COMP_LOOP_C_30;
      WHEN COMP_LOOP_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110110");
        state_var_NS <= COMP_LOOP_C_31;
      WHEN COMP_LOOP_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110111");
        state_var_NS <= COMP_LOOP_C_32;
      WHEN COMP_LOOP_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111000");
        state_var_NS <= COMP_LOOP_C_33;
      WHEN COMP_LOOP_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111001");
        state_var_NS <= COMP_LOOP_C_34;
      WHEN COMP_LOOP_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111010");
        state_var_NS <= COMP_LOOP_C_35;
      WHEN COMP_LOOP_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111011");
        state_var_NS <= COMP_LOOP_C_36;
      WHEN COMP_LOOP_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111100");
        state_var_NS <= COMP_LOOP_C_37;
      WHEN COMP_LOOP_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111101");
        state_var_NS <= COMP_LOOP_C_38;
      WHEN COMP_LOOP_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111110");
        state_var_NS <= COMP_LOOP_C_39;
      WHEN COMP_LOOP_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111111");
        state_var_NS <= COMP_LOOP_C_40;
      WHEN COMP_LOOP_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000000");
        state_var_NS <= COMP_LOOP_C_41;
      WHEN COMP_LOOP_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000001");
        state_var_NS <= COMP_LOOP_C_42;
      WHEN COMP_LOOP_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000010");
        state_var_NS <= COMP_LOOP_C_43;
      WHEN COMP_LOOP_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000011");
        state_var_NS <= COMP_LOOP_C_44;
      WHEN COMP_LOOP_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000100");
        state_var_NS <= COMP_LOOP_C_45;
      WHEN COMP_LOOP_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000101");
        state_var_NS <= COMP_LOOP_C_46;
      WHEN COMP_LOOP_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000110");
        state_var_NS <= COMP_LOOP_C_47;
      WHEN COMP_LOOP_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000111");
        state_var_NS <= COMP_LOOP_C_48;
      WHEN COMP_LOOP_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001000");
        state_var_NS <= COMP_LOOP_C_49;
      WHEN COMP_LOOP_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001001");
        state_var_NS <= COMP_LOOP_C_50;
      WHEN COMP_LOOP_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001010");
        state_var_NS <= COMP_LOOP_C_51;
      WHEN COMP_LOOP_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001011");
        state_var_NS <= COMP_LOOP_C_52;
      WHEN COMP_LOOP_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001100");
        state_var_NS <= COMP_LOOP_C_53;
      WHEN COMP_LOOP_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001101");
        state_var_NS <= COMP_LOOP_C_54;
      WHEN COMP_LOOP_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001110");
        state_var_NS <= COMP_LOOP_C_55;
      WHEN COMP_LOOP_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001111");
        state_var_NS <= COMP_LOOP_C_56;
      WHEN COMP_LOOP_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010000");
        state_var_NS <= COMP_LOOP_C_57;
      WHEN COMP_LOOP_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010001");
        state_var_NS <= COMP_LOOP_C_58;
      WHEN COMP_LOOP_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010010");
        state_var_NS <= COMP_LOOP_C_59;
      WHEN COMP_LOOP_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010011");
        state_var_NS <= COMP_LOOP_C_60;
      WHEN COMP_LOOP_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010100");
        state_var_NS <= COMP_LOOP_C_61;
      WHEN COMP_LOOP_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010101");
        state_var_NS <= COMP_LOOP_C_62;
      WHEN COMP_LOOP_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010110");
        IF ( COMP_LOOP_C_62_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_63;
        END IF;
      WHEN COMP_LOOP_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_0;
      WHEN COMP_LOOP_2_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_1;
      WHEN COMP_LOOP_2_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_2;
      WHEN COMP_LOOP_2_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_3;
      WHEN COMP_LOOP_2_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_4;
      WHEN COMP_LOOP_2_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_5;
      WHEN COMP_LOOP_2_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_6;
      WHEN COMP_LOOP_2_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_7;
      WHEN COMP_LOOP_2_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_8;
      WHEN COMP_LOOP_2_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_9;
      WHEN COMP_LOOP_2_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_10;
      WHEN COMP_LOOP_2_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_11;
      WHEN COMP_LOOP_2_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_12;
      WHEN COMP_LOOP_2_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_13;
      WHEN COMP_LOOP_2_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_14;
      WHEN COMP_LOOP_2_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_15;
      WHEN COMP_LOOP_2_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_16;
      WHEN COMP_LOOP_2_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_17;
      WHEN COMP_LOOP_2_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_18;
      WHEN COMP_LOOP_2_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_19;
      WHEN COMP_LOOP_2_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_20;
      WHEN COMP_LOOP_2_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_21;
      WHEN COMP_LOOP_2_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_22;
      WHEN COMP_LOOP_2_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_23;
      WHEN COMP_LOOP_2_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_24;
      WHEN COMP_LOOP_2_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_25;
      WHEN COMP_LOOP_2_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_26;
      WHEN COMP_LOOP_2_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_27;
      WHEN COMP_LOOP_2_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_28;
      WHEN COMP_LOOP_2_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_29;
      WHEN COMP_LOOP_2_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_30;
      WHEN COMP_LOOP_2_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110110");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_31;
      WHEN COMP_LOOP_2_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110111");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_32;
      WHEN COMP_LOOP_2_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111000");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_33;
      WHEN COMP_LOOP_2_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111001");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_34;
      WHEN COMP_LOOP_2_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111010");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_35;
      WHEN COMP_LOOP_2_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111011");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_36;
      WHEN COMP_LOOP_2_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111100");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_37;
      WHEN COMP_LOOP_2_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111101");
        state_var_NS <= COMP_LOOP_2_modExp_1_while_C_38;
      WHEN COMP_LOOP_2_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111110");
        IF ( COMP_LOOP_2_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_64;
        ELSE
          state_var_NS <= COMP_LOOP_2_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111111");
        state_var_NS <= COMP_LOOP_C_65;
      WHEN COMP_LOOP_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000000");
        state_var_NS <= COMP_LOOP_C_66;
      WHEN COMP_LOOP_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000001");
        state_var_NS <= COMP_LOOP_C_67;
      WHEN COMP_LOOP_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000010");
        state_var_NS <= COMP_LOOP_C_68;
      WHEN COMP_LOOP_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000011");
        state_var_NS <= COMP_LOOP_C_69;
      WHEN COMP_LOOP_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000100");
        state_var_NS <= COMP_LOOP_C_70;
      WHEN COMP_LOOP_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000101");
        state_var_NS <= COMP_LOOP_C_71;
      WHEN COMP_LOOP_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000110");
        state_var_NS <= COMP_LOOP_C_72;
      WHEN COMP_LOOP_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000111");
        state_var_NS <= COMP_LOOP_C_73;
      WHEN COMP_LOOP_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001000");
        state_var_NS <= COMP_LOOP_C_74;
      WHEN COMP_LOOP_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001001");
        state_var_NS <= COMP_LOOP_C_75;
      WHEN COMP_LOOP_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001010");
        state_var_NS <= COMP_LOOP_C_76;
      WHEN COMP_LOOP_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001011");
        state_var_NS <= COMP_LOOP_C_77;
      WHEN COMP_LOOP_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001100");
        state_var_NS <= COMP_LOOP_C_78;
      WHEN COMP_LOOP_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001101");
        state_var_NS <= COMP_LOOP_C_79;
      WHEN COMP_LOOP_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001110");
        state_var_NS <= COMP_LOOP_C_80;
      WHEN COMP_LOOP_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001111");
        state_var_NS <= COMP_LOOP_C_81;
      WHEN COMP_LOOP_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010000");
        state_var_NS <= COMP_LOOP_C_82;
      WHEN COMP_LOOP_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010001");
        state_var_NS <= COMP_LOOP_C_83;
      WHEN COMP_LOOP_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010010");
        state_var_NS <= COMP_LOOP_C_84;
      WHEN COMP_LOOP_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010011");
        state_var_NS <= COMP_LOOP_C_85;
      WHEN COMP_LOOP_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010100");
        state_var_NS <= COMP_LOOP_C_86;
      WHEN COMP_LOOP_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010101");
        state_var_NS <= COMP_LOOP_C_87;
      WHEN COMP_LOOP_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010110");
        state_var_NS <= COMP_LOOP_C_88;
      WHEN COMP_LOOP_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010111");
        state_var_NS <= COMP_LOOP_C_89;
      WHEN COMP_LOOP_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011000");
        state_var_NS <= COMP_LOOP_C_90;
      WHEN COMP_LOOP_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011001");
        state_var_NS <= COMP_LOOP_C_91;
      WHEN COMP_LOOP_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011010");
        state_var_NS <= COMP_LOOP_C_92;
      WHEN COMP_LOOP_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011011");
        state_var_NS <= COMP_LOOP_C_93;
      WHEN COMP_LOOP_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011100");
        state_var_NS <= COMP_LOOP_C_94;
      WHEN COMP_LOOP_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011101");
        state_var_NS <= COMP_LOOP_C_95;
      WHEN COMP_LOOP_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011110");
        state_var_NS <= COMP_LOOP_C_96;
      WHEN COMP_LOOP_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011111");
        state_var_NS <= COMP_LOOP_C_97;
      WHEN COMP_LOOP_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100000");
        state_var_NS <= COMP_LOOP_C_98;
      WHEN COMP_LOOP_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100001");
        state_var_NS <= COMP_LOOP_C_99;
      WHEN COMP_LOOP_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100010");
        state_var_NS <= COMP_LOOP_C_100;
      WHEN COMP_LOOP_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100011");
        state_var_NS <= COMP_LOOP_C_101;
      WHEN COMP_LOOP_C_101 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100100");
        state_var_NS <= COMP_LOOP_C_102;
      WHEN COMP_LOOP_C_102 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100101");
        state_var_NS <= COMP_LOOP_C_103;
      WHEN COMP_LOOP_C_103 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100110");
        state_var_NS <= COMP_LOOP_C_104;
      WHEN COMP_LOOP_C_104 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100111");
        state_var_NS <= COMP_LOOP_C_105;
      WHEN COMP_LOOP_C_105 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101000");
        state_var_NS <= COMP_LOOP_C_106;
      WHEN COMP_LOOP_C_106 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101001");
        state_var_NS <= COMP_LOOP_C_107;
      WHEN COMP_LOOP_C_107 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101010");
        state_var_NS <= COMP_LOOP_C_108;
      WHEN COMP_LOOP_C_108 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101011");
        state_var_NS <= COMP_LOOP_C_109;
      WHEN COMP_LOOP_C_109 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101100");
        state_var_NS <= COMP_LOOP_C_110;
      WHEN COMP_LOOP_C_110 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101101");
        state_var_NS <= COMP_LOOP_C_111;
      WHEN COMP_LOOP_C_111 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101110");
        state_var_NS <= COMP_LOOP_C_112;
      WHEN COMP_LOOP_C_112 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101111");
        state_var_NS <= COMP_LOOP_C_113;
      WHEN COMP_LOOP_C_113 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110000");
        state_var_NS <= COMP_LOOP_C_114;
      WHEN COMP_LOOP_C_114 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110001");
        state_var_NS <= COMP_LOOP_C_115;
      WHEN COMP_LOOP_C_115 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110010");
        state_var_NS <= COMP_LOOP_C_116;
      WHEN COMP_LOOP_C_116 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110011");
        state_var_NS <= COMP_LOOP_C_117;
      WHEN COMP_LOOP_C_117 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110100");
        state_var_NS <= COMP_LOOP_C_118;
      WHEN COMP_LOOP_C_118 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110101");
        state_var_NS <= COMP_LOOP_C_119;
      WHEN COMP_LOOP_C_119 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110110");
        state_var_NS <= COMP_LOOP_C_120;
      WHEN COMP_LOOP_C_120 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110111");
        state_var_NS <= COMP_LOOP_C_121;
      WHEN COMP_LOOP_C_121 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111000");
        state_var_NS <= COMP_LOOP_C_122;
      WHEN COMP_LOOP_C_122 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111001");
        state_var_NS <= COMP_LOOP_C_123;
      WHEN COMP_LOOP_C_123 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111010");
        state_var_NS <= COMP_LOOP_C_124;
      WHEN COMP_LOOP_C_124 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111011");
        IF ( COMP_LOOP_C_124_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_125;
        END IF;
      WHEN COMP_LOOP_C_125 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_0;
      WHEN COMP_LOOP_3_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_1;
      WHEN COMP_LOOP_3_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_2;
      WHEN COMP_LOOP_3_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_3;
      WHEN COMP_LOOP_3_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_4;
      WHEN COMP_LOOP_3_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_5;
      WHEN COMP_LOOP_3_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_6;
      WHEN COMP_LOOP_3_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_7;
      WHEN COMP_LOOP_3_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_8;
      WHEN COMP_LOOP_3_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_9;
      WHEN COMP_LOOP_3_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_10;
      WHEN COMP_LOOP_3_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_11;
      WHEN COMP_LOOP_3_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_12;
      WHEN COMP_LOOP_3_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_13;
      WHEN COMP_LOOP_3_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_14;
      WHEN COMP_LOOP_3_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_15;
      WHEN COMP_LOOP_3_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_16;
      WHEN COMP_LOOP_3_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_17;
      WHEN COMP_LOOP_3_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_18;
      WHEN COMP_LOOP_3_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_19;
      WHEN COMP_LOOP_3_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_20;
      WHEN COMP_LOOP_3_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_21;
      WHEN COMP_LOOP_3_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_22;
      WHEN COMP_LOOP_3_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_23;
      WHEN COMP_LOOP_3_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_24;
      WHEN COMP_LOOP_3_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_25;
      WHEN COMP_LOOP_3_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_26;
      WHEN COMP_LOOP_3_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_27;
      WHEN COMP_LOOP_3_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_28;
      WHEN COMP_LOOP_3_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_29;
      WHEN COMP_LOOP_3_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_30;
      WHEN COMP_LOOP_3_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011011");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_31;
      WHEN COMP_LOOP_3_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011100");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_32;
      WHEN COMP_LOOP_3_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011101");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_33;
      WHEN COMP_LOOP_3_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011110");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_34;
      WHEN COMP_LOOP_3_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011111");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_35;
      WHEN COMP_LOOP_3_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100000");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_36;
      WHEN COMP_LOOP_3_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100001");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_37;
      WHEN COMP_LOOP_3_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100010");
        state_var_NS <= COMP_LOOP_3_modExp_1_while_C_38;
      WHEN COMP_LOOP_3_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100011");
        IF ( COMP_LOOP_3_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_126;
        ELSE
          state_var_NS <= COMP_LOOP_3_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_126 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100100");
        state_var_NS <= COMP_LOOP_C_127;
      WHEN COMP_LOOP_C_127 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100101");
        state_var_NS <= COMP_LOOP_C_128;
      WHEN COMP_LOOP_C_128 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100110");
        state_var_NS <= COMP_LOOP_C_129;
      WHEN COMP_LOOP_C_129 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100111");
        state_var_NS <= COMP_LOOP_C_130;
      WHEN COMP_LOOP_C_130 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101000");
        state_var_NS <= COMP_LOOP_C_131;
      WHEN COMP_LOOP_C_131 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101001");
        state_var_NS <= COMP_LOOP_C_132;
      WHEN COMP_LOOP_C_132 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101010");
        state_var_NS <= COMP_LOOP_C_133;
      WHEN COMP_LOOP_C_133 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101011");
        state_var_NS <= COMP_LOOP_C_134;
      WHEN COMP_LOOP_C_134 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101100");
        state_var_NS <= COMP_LOOP_C_135;
      WHEN COMP_LOOP_C_135 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101101");
        state_var_NS <= COMP_LOOP_C_136;
      WHEN COMP_LOOP_C_136 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101110");
        state_var_NS <= COMP_LOOP_C_137;
      WHEN COMP_LOOP_C_137 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101111");
        state_var_NS <= COMP_LOOP_C_138;
      WHEN COMP_LOOP_C_138 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110000");
        state_var_NS <= COMP_LOOP_C_139;
      WHEN COMP_LOOP_C_139 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110001");
        state_var_NS <= COMP_LOOP_C_140;
      WHEN COMP_LOOP_C_140 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110010");
        state_var_NS <= COMP_LOOP_C_141;
      WHEN COMP_LOOP_C_141 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110011");
        state_var_NS <= COMP_LOOP_C_142;
      WHEN COMP_LOOP_C_142 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110100");
        state_var_NS <= COMP_LOOP_C_143;
      WHEN COMP_LOOP_C_143 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110101");
        state_var_NS <= COMP_LOOP_C_144;
      WHEN COMP_LOOP_C_144 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110110");
        state_var_NS <= COMP_LOOP_C_145;
      WHEN COMP_LOOP_C_145 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110111");
        state_var_NS <= COMP_LOOP_C_146;
      WHEN COMP_LOOP_C_146 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111000");
        state_var_NS <= COMP_LOOP_C_147;
      WHEN COMP_LOOP_C_147 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111001");
        state_var_NS <= COMP_LOOP_C_148;
      WHEN COMP_LOOP_C_148 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111010");
        state_var_NS <= COMP_LOOP_C_149;
      WHEN COMP_LOOP_C_149 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111011");
        state_var_NS <= COMP_LOOP_C_150;
      WHEN COMP_LOOP_C_150 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111100");
        state_var_NS <= COMP_LOOP_C_151;
      WHEN COMP_LOOP_C_151 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111101");
        state_var_NS <= COMP_LOOP_C_152;
      WHEN COMP_LOOP_C_152 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111110");
        state_var_NS <= COMP_LOOP_C_153;
      WHEN COMP_LOOP_C_153 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111111");
        state_var_NS <= COMP_LOOP_C_154;
      WHEN COMP_LOOP_C_154 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000000");
        state_var_NS <= COMP_LOOP_C_155;
      WHEN COMP_LOOP_C_155 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000001");
        state_var_NS <= COMP_LOOP_C_156;
      WHEN COMP_LOOP_C_156 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000010");
        state_var_NS <= COMP_LOOP_C_157;
      WHEN COMP_LOOP_C_157 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000011");
        state_var_NS <= COMP_LOOP_C_158;
      WHEN COMP_LOOP_C_158 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000100");
        state_var_NS <= COMP_LOOP_C_159;
      WHEN COMP_LOOP_C_159 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000101");
        state_var_NS <= COMP_LOOP_C_160;
      WHEN COMP_LOOP_C_160 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000110");
        state_var_NS <= COMP_LOOP_C_161;
      WHEN COMP_LOOP_C_161 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000111");
        state_var_NS <= COMP_LOOP_C_162;
      WHEN COMP_LOOP_C_162 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001000");
        state_var_NS <= COMP_LOOP_C_163;
      WHEN COMP_LOOP_C_163 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001001");
        state_var_NS <= COMP_LOOP_C_164;
      WHEN COMP_LOOP_C_164 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001010");
        state_var_NS <= COMP_LOOP_C_165;
      WHEN COMP_LOOP_C_165 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001011");
        state_var_NS <= COMP_LOOP_C_166;
      WHEN COMP_LOOP_C_166 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001100");
        state_var_NS <= COMP_LOOP_C_167;
      WHEN COMP_LOOP_C_167 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001101");
        state_var_NS <= COMP_LOOP_C_168;
      WHEN COMP_LOOP_C_168 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001110");
        state_var_NS <= COMP_LOOP_C_169;
      WHEN COMP_LOOP_C_169 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001111");
        state_var_NS <= COMP_LOOP_C_170;
      WHEN COMP_LOOP_C_170 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010000");
        state_var_NS <= COMP_LOOP_C_171;
      WHEN COMP_LOOP_C_171 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010001");
        state_var_NS <= COMP_LOOP_C_172;
      WHEN COMP_LOOP_C_172 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010010");
        state_var_NS <= COMP_LOOP_C_173;
      WHEN COMP_LOOP_C_173 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010011");
        state_var_NS <= COMP_LOOP_C_174;
      WHEN COMP_LOOP_C_174 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010100");
        state_var_NS <= COMP_LOOP_C_175;
      WHEN COMP_LOOP_C_175 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010101");
        state_var_NS <= COMP_LOOP_C_176;
      WHEN COMP_LOOP_C_176 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010110");
        state_var_NS <= COMP_LOOP_C_177;
      WHEN COMP_LOOP_C_177 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010111");
        state_var_NS <= COMP_LOOP_C_178;
      WHEN COMP_LOOP_C_178 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011000");
        state_var_NS <= COMP_LOOP_C_179;
      WHEN COMP_LOOP_C_179 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011001");
        state_var_NS <= COMP_LOOP_C_180;
      WHEN COMP_LOOP_C_180 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011010");
        state_var_NS <= COMP_LOOP_C_181;
      WHEN COMP_LOOP_C_181 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011011");
        state_var_NS <= COMP_LOOP_C_182;
      WHEN COMP_LOOP_C_182 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011100");
        state_var_NS <= COMP_LOOP_C_183;
      WHEN COMP_LOOP_C_183 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011101");
        state_var_NS <= COMP_LOOP_C_184;
      WHEN COMP_LOOP_C_184 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011110");
        state_var_NS <= COMP_LOOP_C_185;
      WHEN COMP_LOOP_C_185 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011111");
        state_var_NS <= COMP_LOOP_C_186;
      WHEN COMP_LOOP_C_186 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100000");
        IF ( COMP_LOOP_C_186_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_187;
        END IF;
      WHEN COMP_LOOP_C_187 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_0;
      WHEN COMP_LOOP_4_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_1;
      WHEN COMP_LOOP_4_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_2;
      WHEN COMP_LOOP_4_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_3;
      WHEN COMP_LOOP_4_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_4;
      WHEN COMP_LOOP_4_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_5;
      WHEN COMP_LOOP_4_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_6;
      WHEN COMP_LOOP_4_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_7;
      WHEN COMP_LOOP_4_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_8;
      WHEN COMP_LOOP_4_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_9;
      WHEN COMP_LOOP_4_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_10;
      WHEN COMP_LOOP_4_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_11;
      WHEN COMP_LOOP_4_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_12;
      WHEN COMP_LOOP_4_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_13;
      WHEN COMP_LOOP_4_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_14;
      WHEN COMP_LOOP_4_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_15;
      WHEN COMP_LOOP_4_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_16;
      WHEN COMP_LOOP_4_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_17;
      WHEN COMP_LOOP_4_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_18;
      WHEN COMP_LOOP_4_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_19;
      WHEN COMP_LOOP_4_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_20;
      WHEN COMP_LOOP_4_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_21;
      WHEN COMP_LOOP_4_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_22;
      WHEN COMP_LOOP_4_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_23;
      WHEN COMP_LOOP_4_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_24;
      WHEN COMP_LOOP_4_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_25;
      WHEN COMP_LOOP_4_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_26;
      WHEN COMP_LOOP_4_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_27;
      WHEN COMP_LOOP_4_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_28;
      WHEN COMP_LOOP_4_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_29;
      WHEN COMP_LOOP_4_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_30;
      WHEN COMP_LOOP_4_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000000");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_31;
      WHEN COMP_LOOP_4_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000001");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_32;
      WHEN COMP_LOOP_4_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000010");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_33;
      WHEN COMP_LOOP_4_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000011");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_34;
      WHEN COMP_LOOP_4_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000100");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_35;
      WHEN COMP_LOOP_4_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000101");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_36;
      WHEN COMP_LOOP_4_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000110");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_37;
      WHEN COMP_LOOP_4_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000111");
        state_var_NS <= COMP_LOOP_4_modExp_1_while_C_38;
      WHEN COMP_LOOP_4_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001000");
        IF ( COMP_LOOP_4_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_188;
        ELSE
          state_var_NS <= COMP_LOOP_4_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_188 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001001");
        state_var_NS <= COMP_LOOP_C_189;
      WHEN COMP_LOOP_C_189 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001010");
        state_var_NS <= COMP_LOOP_C_190;
      WHEN COMP_LOOP_C_190 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001011");
        state_var_NS <= COMP_LOOP_C_191;
      WHEN COMP_LOOP_C_191 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001100");
        state_var_NS <= COMP_LOOP_C_192;
      WHEN COMP_LOOP_C_192 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001101");
        state_var_NS <= COMP_LOOP_C_193;
      WHEN COMP_LOOP_C_193 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001110");
        state_var_NS <= COMP_LOOP_C_194;
      WHEN COMP_LOOP_C_194 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001111");
        state_var_NS <= COMP_LOOP_C_195;
      WHEN COMP_LOOP_C_195 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010000");
        state_var_NS <= COMP_LOOP_C_196;
      WHEN COMP_LOOP_C_196 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010001");
        state_var_NS <= COMP_LOOP_C_197;
      WHEN COMP_LOOP_C_197 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010010");
        state_var_NS <= COMP_LOOP_C_198;
      WHEN COMP_LOOP_C_198 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010011");
        state_var_NS <= COMP_LOOP_C_199;
      WHEN COMP_LOOP_C_199 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010100");
        state_var_NS <= COMP_LOOP_C_200;
      WHEN COMP_LOOP_C_200 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010101");
        state_var_NS <= COMP_LOOP_C_201;
      WHEN COMP_LOOP_C_201 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010110");
        state_var_NS <= COMP_LOOP_C_202;
      WHEN COMP_LOOP_C_202 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010111");
        state_var_NS <= COMP_LOOP_C_203;
      WHEN COMP_LOOP_C_203 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011000");
        state_var_NS <= COMP_LOOP_C_204;
      WHEN COMP_LOOP_C_204 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011001");
        state_var_NS <= COMP_LOOP_C_205;
      WHEN COMP_LOOP_C_205 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011010");
        state_var_NS <= COMP_LOOP_C_206;
      WHEN COMP_LOOP_C_206 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011011");
        state_var_NS <= COMP_LOOP_C_207;
      WHEN COMP_LOOP_C_207 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011100");
        state_var_NS <= COMP_LOOP_C_208;
      WHEN COMP_LOOP_C_208 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011101");
        state_var_NS <= COMP_LOOP_C_209;
      WHEN COMP_LOOP_C_209 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011110");
        state_var_NS <= COMP_LOOP_C_210;
      WHEN COMP_LOOP_C_210 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011111");
        state_var_NS <= COMP_LOOP_C_211;
      WHEN COMP_LOOP_C_211 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100000");
        state_var_NS <= COMP_LOOP_C_212;
      WHEN COMP_LOOP_C_212 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100001");
        state_var_NS <= COMP_LOOP_C_213;
      WHEN COMP_LOOP_C_213 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100010");
        state_var_NS <= COMP_LOOP_C_214;
      WHEN COMP_LOOP_C_214 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100011");
        state_var_NS <= COMP_LOOP_C_215;
      WHEN COMP_LOOP_C_215 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100100");
        state_var_NS <= COMP_LOOP_C_216;
      WHEN COMP_LOOP_C_216 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100101");
        state_var_NS <= COMP_LOOP_C_217;
      WHEN COMP_LOOP_C_217 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100110");
        state_var_NS <= COMP_LOOP_C_218;
      WHEN COMP_LOOP_C_218 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100111");
        state_var_NS <= COMP_LOOP_C_219;
      WHEN COMP_LOOP_C_219 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101000");
        state_var_NS <= COMP_LOOP_C_220;
      WHEN COMP_LOOP_C_220 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101001");
        state_var_NS <= COMP_LOOP_C_221;
      WHEN COMP_LOOP_C_221 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101010");
        state_var_NS <= COMP_LOOP_C_222;
      WHEN COMP_LOOP_C_222 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101011");
        state_var_NS <= COMP_LOOP_C_223;
      WHEN COMP_LOOP_C_223 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101100");
        state_var_NS <= COMP_LOOP_C_224;
      WHEN COMP_LOOP_C_224 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101101");
        state_var_NS <= COMP_LOOP_C_225;
      WHEN COMP_LOOP_C_225 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101110");
        state_var_NS <= COMP_LOOP_C_226;
      WHEN COMP_LOOP_C_226 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101111");
        state_var_NS <= COMP_LOOP_C_227;
      WHEN COMP_LOOP_C_227 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110000");
        state_var_NS <= COMP_LOOP_C_228;
      WHEN COMP_LOOP_C_228 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110001");
        state_var_NS <= COMP_LOOP_C_229;
      WHEN COMP_LOOP_C_229 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110010");
        state_var_NS <= COMP_LOOP_C_230;
      WHEN COMP_LOOP_C_230 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110011");
        state_var_NS <= COMP_LOOP_C_231;
      WHEN COMP_LOOP_C_231 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110100");
        state_var_NS <= COMP_LOOP_C_232;
      WHEN COMP_LOOP_C_232 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110101");
        state_var_NS <= COMP_LOOP_C_233;
      WHEN COMP_LOOP_C_233 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110110");
        state_var_NS <= COMP_LOOP_C_234;
      WHEN COMP_LOOP_C_234 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110111");
        state_var_NS <= COMP_LOOP_C_235;
      WHEN COMP_LOOP_C_235 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111000");
        state_var_NS <= COMP_LOOP_C_236;
      WHEN COMP_LOOP_C_236 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111001");
        state_var_NS <= COMP_LOOP_C_237;
      WHEN COMP_LOOP_C_237 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111010");
        state_var_NS <= COMP_LOOP_C_238;
      WHEN COMP_LOOP_C_238 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111011");
        state_var_NS <= COMP_LOOP_C_239;
      WHEN COMP_LOOP_C_239 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111100");
        state_var_NS <= COMP_LOOP_C_240;
      WHEN COMP_LOOP_C_240 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111101");
        state_var_NS <= COMP_LOOP_C_241;
      WHEN COMP_LOOP_C_241 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111110");
        state_var_NS <= COMP_LOOP_C_242;
      WHEN COMP_LOOP_C_242 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111111");
        state_var_NS <= COMP_LOOP_C_243;
      WHEN COMP_LOOP_C_243 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000000");
        state_var_NS <= COMP_LOOP_C_244;
      WHEN COMP_LOOP_C_244 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000001");
        state_var_NS <= COMP_LOOP_C_245;
      WHEN COMP_LOOP_C_245 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000010");
        state_var_NS <= COMP_LOOP_C_246;
      WHEN COMP_LOOP_C_246 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000011");
        state_var_NS <= COMP_LOOP_C_247;
      WHEN COMP_LOOP_C_247 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000100");
        state_var_NS <= COMP_LOOP_C_248;
      WHEN COMP_LOOP_C_248 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000101");
        IF ( COMP_LOOP_C_248_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_249;
        END IF;
      WHEN COMP_LOOP_C_249 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_0;
      WHEN COMP_LOOP_5_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_1;
      WHEN COMP_LOOP_5_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_2;
      WHEN COMP_LOOP_5_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_3;
      WHEN COMP_LOOP_5_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_4;
      WHEN COMP_LOOP_5_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_5;
      WHEN COMP_LOOP_5_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_6;
      WHEN COMP_LOOP_5_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_7;
      WHEN COMP_LOOP_5_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_8;
      WHEN COMP_LOOP_5_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_9;
      WHEN COMP_LOOP_5_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_10;
      WHEN COMP_LOOP_5_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_11;
      WHEN COMP_LOOP_5_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_12;
      WHEN COMP_LOOP_5_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_13;
      WHEN COMP_LOOP_5_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_14;
      WHEN COMP_LOOP_5_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_15;
      WHEN COMP_LOOP_5_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_16;
      WHEN COMP_LOOP_5_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_17;
      WHEN COMP_LOOP_5_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_18;
      WHEN COMP_LOOP_5_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_19;
      WHEN COMP_LOOP_5_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_20;
      WHEN COMP_LOOP_5_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_21;
      WHEN COMP_LOOP_5_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_22;
      WHEN COMP_LOOP_5_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_23;
      WHEN COMP_LOOP_5_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_24;
      WHEN COMP_LOOP_5_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_25;
      WHEN COMP_LOOP_5_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_26;
      WHEN COMP_LOOP_5_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_27;
      WHEN COMP_LOOP_5_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_28;
      WHEN COMP_LOOP_5_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_29;
      WHEN COMP_LOOP_5_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_30;
      WHEN COMP_LOOP_5_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100101");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_31;
      WHEN COMP_LOOP_5_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100110");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_32;
      WHEN COMP_LOOP_5_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100111");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_33;
      WHEN COMP_LOOP_5_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101000");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_34;
      WHEN COMP_LOOP_5_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101001");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_35;
      WHEN COMP_LOOP_5_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101010");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_36;
      WHEN COMP_LOOP_5_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101011");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_37;
      WHEN COMP_LOOP_5_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101100");
        state_var_NS <= COMP_LOOP_5_modExp_1_while_C_38;
      WHEN COMP_LOOP_5_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101101");
        IF ( COMP_LOOP_5_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_250;
        ELSE
          state_var_NS <= COMP_LOOP_5_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_250 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101110");
        state_var_NS <= COMP_LOOP_C_251;
      WHEN COMP_LOOP_C_251 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101111");
        state_var_NS <= COMP_LOOP_C_252;
      WHEN COMP_LOOP_C_252 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110000");
        state_var_NS <= COMP_LOOP_C_253;
      WHEN COMP_LOOP_C_253 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110001");
        state_var_NS <= COMP_LOOP_C_254;
      WHEN COMP_LOOP_C_254 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110010");
        state_var_NS <= COMP_LOOP_C_255;
      WHEN COMP_LOOP_C_255 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110011");
        state_var_NS <= COMP_LOOP_C_256;
      WHEN COMP_LOOP_C_256 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110100");
        state_var_NS <= COMP_LOOP_C_257;
      WHEN COMP_LOOP_C_257 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110101");
        state_var_NS <= COMP_LOOP_C_258;
      WHEN COMP_LOOP_C_258 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110110");
        state_var_NS <= COMP_LOOP_C_259;
      WHEN COMP_LOOP_C_259 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110111");
        state_var_NS <= COMP_LOOP_C_260;
      WHEN COMP_LOOP_C_260 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111000");
        state_var_NS <= COMP_LOOP_C_261;
      WHEN COMP_LOOP_C_261 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111001");
        state_var_NS <= COMP_LOOP_C_262;
      WHEN COMP_LOOP_C_262 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111010");
        state_var_NS <= COMP_LOOP_C_263;
      WHEN COMP_LOOP_C_263 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111011");
        state_var_NS <= COMP_LOOP_C_264;
      WHEN COMP_LOOP_C_264 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111100");
        state_var_NS <= COMP_LOOP_C_265;
      WHEN COMP_LOOP_C_265 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111101");
        state_var_NS <= COMP_LOOP_C_266;
      WHEN COMP_LOOP_C_266 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111110");
        state_var_NS <= COMP_LOOP_C_267;
      WHEN COMP_LOOP_C_267 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111111");
        state_var_NS <= COMP_LOOP_C_268;
      WHEN COMP_LOOP_C_268 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000000");
        state_var_NS <= COMP_LOOP_C_269;
      WHEN COMP_LOOP_C_269 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000001");
        state_var_NS <= COMP_LOOP_C_270;
      WHEN COMP_LOOP_C_270 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000010");
        state_var_NS <= COMP_LOOP_C_271;
      WHEN COMP_LOOP_C_271 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000011");
        state_var_NS <= COMP_LOOP_C_272;
      WHEN COMP_LOOP_C_272 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000100");
        state_var_NS <= COMP_LOOP_C_273;
      WHEN COMP_LOOP_C_273 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000101");
        state_var_NS <= COMP_LOOP_C_274;
      WHEN COMP_LOOP_C_274 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000110");
        state_var_NS <= COMP_LOOP_C_275;
      WHEN COMP_LOOP_C_275 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000111");
        state_var_NS <= COMP_LOOP_C_276;
      WHEN COMP_LOOP_C_276 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001000");
        state_var_NS <= COMP_LOOP_C_277;
      WHEN COMP_LOOP_C_277 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001001");
        state_var_NS <= COMP_LOOP_C_278;
      WHEN COMP_LOOP_C_278 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001010");
        state_var_NS <= COMP_LOOP_C_279;
      WHEN COMP_LOOP_C_279 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001011");
        state_var_NS <= COMP_LOOP_C_280;
      WHEN COMP_LOOP_C_280 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001100");
        state_var_NS <= COMP_LOOP_C_281;
      WHEN COMP_LOOP_C_281 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001101");
        state_var_NS <= COMP_LOOP_C_282;
      WHEN COMP_LOOP_C_282 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001110");
        state_var_NS <= COMP_LOOP_C_283;
      WHEN COMP_LOOP_C_283 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001111");
        state_var_NS <= COMP_LOOP_C_284;
      WHEN COMP_LOOP_C_284 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010000");
        state_var_NS <= COMP_LOOP_C_285;
      WHEN COMP_LOOP_C_285 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010001");
        state_var_NS <= COMP_LOOP_C_286;
      WHEN COMP_LOOP_C_286 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010010");
        state_var_NS <= COMP_LOOP_C_287;
      WHEN COMP_LOOP_C_287 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010011");
        state_var_NS <= COMP_LOOP_C_288;
      WHEN COMP_LOOP_C_288 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010100");
        state_var_NS <= COMP_LOOP_C_289;
      WHEN COMP_LOOP_C_289 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010101");
        state_var_NS <= COMP_LOOP_C_290;
      WHEN COMP_LOOP_C_290 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010110");
        state_var_NS <= COMP_LOOP_C_291;
      WHEN COMP_LOOP_C_291 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010111");
        state_var_NS <= COMP_LOOP_C_292;
      WHEN COMP_LOOP_C_292 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011000");
        state_var_NS <= COMP_LOOP_C_293;
      WHEN COMP_LOOP_C_293 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011001");
        state_var_NS <= COMP_LOOP_C_294;
      WHEN COMP_LOOP_C_294 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011010");
        state_var_NS <= COMP_LOOP_C_295;
      WHEN COMP_LOOP_C_295 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011011");
        state_var_NS <= COMP_LOOP_C_296;
      WHEN COMP_LOOP_C_296 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011100");
        state_var_NS <= COMP_LOOP_C_297;
      WHEN COMP_LOOP_C_297 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011101");
        state_var_NS <= COMP_LOOP_C_298;
      WHEN COMP_LOOP_C_298 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011110");
        state_var_NS <= COMP_LOOP_C_299;
      WHEN COMP_LOOP_C_299 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011111");
        state_var_NS <= COMP_LOOP_C_300;
      WHEN COMP_LOOP_C_300 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100000");
        state_var_NS <= COMP_LOOP_C_301;
      WHEN COMP_LOOP_C_301 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100001");
        state_var_NS <= COMP_LOOP_C_302;
      WHEN COMP_LOOP_C_302 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100010");
        state_var_NS <= COMP_LOOP_C_303;
      WHEN COMP_LOOP_C_303 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100011");
        state_var_NS <= COMP_LOOP_C_304;
      WHEN COMP_LOOP_C_304 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100100");
        state_var_NS <= COMP_LOOP_C_305;
      WHEN COMP_LOOP_C_305 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100101");
        state_var_NS <= COMP_LOOP_C_306;
      WHEN COMP_LOOP_C_306 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100110");
        state_var_NS <= COMP_LOOP_C_307;
      WHEN COMP_LOOP_C_307 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100111");
        state_var_NS <= COMP_LOOP_C_308;
      WHEN COMP_LOOP_C_308 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101000");
        state_var_NS <= COMP_LOOP_C_309;
      WHEN COMP_LOOP_C_309 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101001");
        state_var_NS <= COMP_LOOP_C_310;
      WHEN COMP_LOOP_C_310 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101010");
        IF ( COMP_LOOP_C_310_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_311;
        END IF;
      WHEN COMP_LOOP_C_311 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_0;
      WHEN COMP_LOOP_6_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_1;
      WHEN COMP_LOOP_6_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_2;
      WHEN COMP_LOOP_6_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_3;
      WHEN COMP_LOOP_6_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_4;
      WHEN COMP_LOOP_6_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_5;
      WHEN COMP_LOOP_6_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_6;
      WHEN COMP_LOOP_6_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_7;
      WHEN COMP_LOOP_6_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_8;
      WHEN COMP_LOOP_6_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_9;
      WHEN COMP_LOOP_6_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_10;
      WHEN COMP_LOOP_6_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_11;
      WHEN COMP_LOOP_6_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_12;
      WHEN COMP_LOOP_6_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_13;
      WHEN COMP_LOOP_6_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_14;
      WHEN COMP_LOOP_6_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_15;
      WHEN COMP_LOOP_6_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_16;
      WHEN COMP_LOOP_6_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_17;
      WHEN COMP_LOOP_6_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_18;
      WHEN COMP_LOOP_6_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_19;
      WHEN COMP_LOOP_6_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_20;
      WHEN COMP_LOOP_6_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_21;
      WHEN COMP_LOOP_6_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_22;
      WHEN COMP_LOOP_6_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_23;
      WHEN COMP_LOOP_6_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_24;
      WHEN COMP_LOOP_6_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_25;
      WHEN COMP_LOOP_6_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_26;
      WHEN COMP_LOOP_6_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_27;
      WHEN COMP_LOOP_6_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_28;
      WHEN COMP_LOOP_6_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_29;
      WHEN COMP_LOOP_6_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_30;
      WHEN COMP_LOOP_6_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001010");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_31;
      WHEN COMP_LOOP_6_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001011");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_32;
      WHEN COMP_LOOP_6_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001100");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_33;
      WHEN COMP_LOOP_6_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001101");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_34;
      WHEN COMP_LOOP_6_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001110");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_35;
      WHEN COMP_LOOP_6_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001111");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_36;
      WHEN COMP_LOOP_6_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010000");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_37;
      WHEN COMP_LOOP_6_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010001");
        state_var_NS <= COMP_LOOP_6_modExp_1_while_C_38;
      WHEN COMP_LOOP_6_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010010");
        IF ( COMP_LOOP_6_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_312;
        ELSE
          state_var_NS <= COMP_LOOP_6_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_312 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010011");
        state_var_NS <= COMP_LOOP_C_313;
      WHEN COMP_LOOP_C_313 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010100");
        state_var_NS <= COMP_LOOP_C_314;
      WHEN COMP_LOOP_C_314 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010101");
        state_var_NS <= COMP_LOOP_C_315;
      WHEN COMP_LOOP_C_315 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010110");
        state_var_NS <= COMP_LOOP_C_316;
      WHEN COMP_LOOP_C_316 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010111");
        state_var_NS <= COMP_LOOP_C_317;
      WHEN COMP_LOOP_C_317 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011000");
        state_var_NS <= COMP_LOOP_C_318;
      WHEN COMP_LOOP_C_318 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011001");
        state_var_NS <= COMP_LOOP_C_319;
      WHEN COMP_LOOP_C_319 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011010");
        state_var_NS <= COMP_LOOP_C_320;
      WHEN COMP_LOOP_C_320 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011011");
        state_var_NS <= COMP_LOOP_C_321;
      WHEN COMP_LOOP_C_321 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011100");
        state_var_NS <= COMP_LOOP_C_322;
      WHEN COMP_LOOP_C_322 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011101");
        state_var_NS <= COMP_LOOP_C_323;
      WHEN COMP_LOOP_C_323 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011110");
        state_var_NS <= COMP_LOOP_C_324;
      WHEN COMP_LOOP_C_324 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011111");
        state_var_NS <= COMP_LOOP_C_325;
      WHEN COMP_LOOP_C_325 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100000");
        state_var_NS <= COMP_LOOP_C_326;
      WHEN COMP_LOOP_C_326 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100001");
        state_var_NS <= COMP_LOOP_C_327;
      WHEN COMP_LOOP_C_327 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100010");
        state_var_NS <= COMP_LOOP_C_328;
      WHEN COMP_LOOP_C_328 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100011");
        state_var_NS <= COMP_LOOP_C_329;
      WHEN COMP_LOOP_C_329 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100100");
        state_var_NS <= COMP_LOOP_C_330;
      WHEN COMP_LOOP_C_330 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100101");
        state_var_NS <= COMP_LOOP_C_331;
      WHEN COMP_LOOP_C_331 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100110");
        state_var_NS <= COMP_LOOP_C_332;
      WHEN COMP_LOOP_C_332 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100111");
        state_var_NS <= COMP_LOOP_C_333;
      WHEN COMP_LOOP_C_333 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101000");
        state_var_NS <= COMP_LOOP_C_334;
      WHEN COMP_LOOP_C_334 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101001");
        state_var_NS <= COMP_LOOP_C_335;
      WHEN COMP_LOOP_C_335 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101010");
        state_var_NS <= COMP_LOOP_C_336;
      WHEN COMP_LOOP_C_336 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101011");
        state_var_NS <= COMP_LOOP_C_337;
      WHEN COMP_LOOP_C_337 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101100");
        state_var_NS <= COMP_LOOP_C_338;
      WHEN COMP_LOOP_C_338 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101101");
        state_var_NS <= COMP_LOOP_C_339;
      WHEN COMP_LOOP_C_339 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101110");
        state_var_NS <= COMP_LOOP_C_340;
      WHEN COMP_LOOP_C_340 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101111");
        state_var_NS <= COMP_LOOP_C_341;
      WHEN COMP_LOOP_C_341 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110000");
        state_var_NS <= COMP_LOOP_C_342;
      WHEN COMP_LOOP_C_342 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110001");
        state_var_NS <= COMP_LOOP_C_343;
      WHEN COMP_LOOP_C_343 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110010");
        state_var_NS <= COMP_LOOP_C_344;
      WHEN COMP_LOOP_C_344 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110011");
        state_var_NS <= COMP_LOOP_C_345;
      WHEN COMP_LOOP_C_345 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110100");
        state_var_NS <= COMP_LOOP_C_346;
      WHEN COMP_LOOP_C_346 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110101");
        state_var_NS <= COMP_LOOP_C_347;
      WHEN COMP_LOOP_C_347 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110110");
        state_var_NS <= COMP_LOOP_C_348;
      WHEN COMP_LOOP_C_348 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110111");
        state_var_NS <= COMP_LOOP_C_349;
      WHEN COMP_LOOP_C_349 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111000");
        state_var_NS <= COMP_LOOP_C_350;
      WHEN COMP_LOOP_C_350 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111001");
        state_var_NS <= COMP_LOOP_C_351;
      WHEN COMP_LOOP_C_351 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111010");
        state_var_NS <= COMP_LOOP_C_352;
      WHEN COMP_LOOP_C_352 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111011");
        state_var_NS <= COMP_LOOP_C_353;
      WHEN COMP_LOOP_C_353 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111100");
        state_var_NS <= COMP_LOOP_C_354;
      WHEN COMP_LOOP_C_354 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111101");
        state_var_NS <= COMP_LOOP_C_355;
      WHEN COMP_LOOP_C_355 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111110");
        state_var_NS <= COMP_LOOP_C_356;
      WHEN COMP_LOOP_C_356 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111111");
        state_var_NS <= COMP_LOOP_C_357;
      WHEN COMP_LOOP_C_357 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000000");
        state_var_NS <= COMP_LOOP_C_358;
      WHEN COMP_LOOP_C_358 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000001");
        state_var_NS <= COMP_LOOP_C_359;
      WHEN COMP_LOOP_C_359 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000010");
        state_var_NS <= COMP_LOOP_C_360;
      WHEN COMP_LOOP_C_360 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000011");
        state_var_NS <= COMP_LOOP_C_361;
      WHEN COMP_LOOP_C_361 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000100");
        state_var_NS <= COMP_LOOP_C_362;
      WHEN COMP_LOOP_C_362 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000101");
        state_var_NS <= COMP_LOOP_C_363;
      WHEN COMP_LOOP_C_363 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000110");
        state_var_NS <= COMP_LOOP_C_364;
      WHEN COMP_LOOP_C_364 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000111");
        state_var_NS <= COMP_LOOP_C_365;
      WHEN COMP_LOOP_C_365 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001000");
        state_var_NS <= COMP_LOOP_C_366;
      WHEN COMP_LOOP_C_366 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001001");
        state_var_NS <= COMP_LOOP_C_367;
      WHEN COMP_LOOP_C_367 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001010");
        state_var_NS <= COMP_LOOP_C_368;
      WHEN COMP_LOOP_C_368 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001011");
        state_var_NS <= COMP_LOOP_C_369;
      WHEN COMP_LOOP_C_369 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001100");
        state_var_NS <= COMP_LOOP_C_370;
      WHEN COMP_LOOP_C_370 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001101");
        state_var_NS <= COMP_LOOP_C_371;
      WHEN COMP_LOOP_C_371 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001110");
        state_var_NS <= COMP_LOOP_C_372;
      WHEN COMP_LOOP_C_372 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001111");
        IF ( COMP_LOOP_C_372_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_373;
        END IF;
      WHEN COMP_LOOP_C_373 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_0;
      WHEN COMP_LOOP_7_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_1;
      WHEN COMP_LOOP_7_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_2;
      WHEN COMP_LOOP_7_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_3;
      WHEN COMP_LOOP_7_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_4;
      WHEN COMP_LOOP_7_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_5;
      WHEN COMP_LOOP_7_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_6;
      WHEN COMP_LOOP_7_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_7;
      WHEN COMP_LOOP_7_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_8;
      WHEN COMP_LOOP_7_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_9;
      WHEN COMP_LOOP_7_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_10;
      WHEN COMP_LOOP_7_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_11;
      WHEN COMP_LOOP_7_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_12;
      WHEN COMP_LOOP_7_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_13;
      WHEN COMP_LOOP_7_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_14;
      WHEN COMP_LOOP_7_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_15;
      WHEN COMP_LOOP_7_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_16;
      WHEN COMP_LOOP_7_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_17;
      WHEN COMP_LOOP_7_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_18;
      WHEN COMP_LOOP_7_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_19;
      WHEN COMP_LOOP_7_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_20;
      WHEN COMP_LOOP_7_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_21;
      WHEN COMP_LOOP_7_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_22;
      WHEN COMP_LOOP_7_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_23;
      WHEN COMP_LOOP_7_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_24;
      WHEN COMP_LOOP_7_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_25;
      WHEN COMP_LOOP_7_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_26;
      WHEN COMP_LOOP_7_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_27;
      WHEN COMP_LOOP_7_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_28;
      WHEN COMP_LOOP_7_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_29;
      WHEN COMP_LOOP_7_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_30;
      WHEN COMP_LOOP_7_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101111");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_31;
      WHEN COMP_LOOP_7_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110000");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_32;
      WHEN COMP_LOOP_7_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110001");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_33;
      WHEN COMP_LOOP_7_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110010");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_34;
      WHEN COMP_LOOP_7_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110011");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_35;
      WHEN COMP_LOOP_7_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110100");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_36;
      WHEN COMP_LOOP_7_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110101");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_37;
      WHEN COMP_LOOP_7_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110110");
        state_var_NS <= COMP_LOOP_7_modExp_1_while_C_38;
      WHEN COMP_LOOP_7_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110111");
        IF ( COMP_LOOP_7_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_374;
        ELSE
          state_var_NS <= COMP_LOOP_7_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_374 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111000");
        state_var_NS <= COMP_LOOP_C_375;
      WHEN COMP_LOOP_C_375 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111001");
        state_var_NS <= COMP_LOOP_C_376;
      WHEN COMP_LOOP_C_376 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111010");
        state_var_NS <= COMP_LOOP_C_377;
      WHEN COMP_LOOP_C_377 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111011");
        state_var_NS <= COMP_LOOP_C_378;
      WHEN COMP_LOOP_C_378 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111100");
        state_var_NS <= COMP_LOOP_C_379;
      WHEN COMP_LOOP_C_379 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111101");
        state_var_NS <= COMP_LOOP_C_380;
      WHEN COMP_LOOP_C_380 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111110");
        state_var_NS <= COMP_LOOP_C_381;
      WHEN COMP_LOOP_C_381 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111111");
        state_var_NS <= COMP_LOOP_C_382;
      WHEN COMP_LOOP_C_382 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000000");
        state_var_NS <= COMP_LOOP_C_383;
      WHEN COMP_LOOP_C_383 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000001");
        state_var_NS <= COMP_LOOP_C_384;
      WHEN COMP_LOOP_C_384 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000010");
        state_var_NS <= COMP_LOOP_C_385;
      WHEN COMP_LOOP_C_385 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000011");
        state_var_NS <= COMP_LOOP_C_386;
      WHEN COMP_LOOP_C_386 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000100");
        state_var_NS <= COMP_LOOP_C_387;
      WHEN COMP_LOOP_C_387 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000101");
        state_var_NS <= COMP_LOOP_C_388;
      WHEN COMP_LOOP_C_388 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000110");
        state_var_NS <= COMP_LOOP_C_389;
      WHEN COMP_LOOP_C_389 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000111");
        state_var_NS <= COMP_LOOP_C_390;
      WHEN COMP_LOOP_C_390 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001000");
        state_var_NS <= COMP_LOOP_C_391;
      WHEN COMP_LOOP_C_391 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001001");
        state_var_NS <= COMP_LOOP_C_392;
      WHEN COMP_LOOP_C_392 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001010");
        state_var_NS <= COMP_LOOP_C_393;
      WHEN COMP_LOOP_C_393 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001011");
        state_var_NS <= COMP_LOOP_C_394;
      WHEN COMP_LOOP_C_394 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001100");
        state_var_NS <= COMP_LOOP_C_395;
      WHEN COMP_LOOP_C_395 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001101");
        state_var_NS <= COMP_LOOP_C_396;
      WHEN COMP_LOOP_C_396 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001110");
        state_var_NS <= COMP_LOOP_C_397;
      WHEN COMP_LOOP_C_397 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001111");
        state_var_NS <= COMP_LOOP_C_398;
      WHEN COMP_LOOP_C_398 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010000");
        state_var_NS <= COMP_LOOP_C_399;
      WHEN COMP_LOOP_C_399 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010001");
        state_var_NS <= COMP_LOOP_C_400;
      WHEN COMP_LOOP_C_400 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010010");
        state_var_NS <= COMP_LOOP_C_401;
      WHEN COMP_LOOP_C_401 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010011");
        state_var_NS <= COMP_LOOP_C_402;
      WHEN COMP_LOOP_C_402 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010100");
        state_var_NS <= COMP_LOOP_C_403;
      WHEN COMP_LOOP_C_403 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010101");
        state_var_NS <= COMP_LOOP_C_404;
      WHEN COMP_LOOP_C_404 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010110");
        state_var_NS <= COMP_LOOP_C_405;
      WHEN COMP_LOOP_C_405 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010111");
        state_var_NS <= COMP_LOOP_C_406;
      WHEN COMP_LOOP_C_406 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011000");
        state_var_NS <= COMP_LOOP_C_407;
      WHEN COMP_LOOP_C_407 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011001");
        state_var_NS <= COMP_LOOP_C_408;
      WHEN COMP_LOOP_C_408 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011010");
        state_var_NS <= COMP_LOOP_C_409;
      WHEN COMP_LOOP_C_409 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011011");
        state_var_NS <= COMP_LOOP_C_410;
      WHEN COMP_LOOP_C_410 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011100");
        state_var_NS <= COMP_LOOP_C_411;
      WHEN COMP_LOOP_C_411 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011101");
        state_var_NS <= COMP_LOOP_C_412;
      WHEN COMP_LOOP_C_412 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011110");
        state_var_NS <= COMP_LOOP_C_413;
      WHEN COMP_LOOP_C_413 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011111");
        state_var_NS <= COMP_LOOP_C_414;
      WHEN COMP_LOOP_C_414 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100000");
        state_var_NS <= COMP_LOOP_C_415;
      WHEN COMP_LOOP_C_415 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100001");
        state_var_NS <= COMP_LOOP_C_416;
      WHEN COMP_LOOP_C_416 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100010");
        state_var_NS <= COMP_LOOP_C_417;
      WHEN COMP_LOOP_C_417 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100011");
        state_var_NS <= COMP_LOOP_C_418;
      WHEN COMP_LOOP_C_418 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100100");
        state_var_NS <= COMP_LOOP_C_419;
      WHEN COMP_LOOP_C_419 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100101");
        state_var_NS <= COMP_LOOP_C_420;
      WHEN COMP_LOOP_C_420 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100110");
        state_var_NS <= COMP_LOOP_C_421;
      WHEN COMP_LOOP_C_421 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100111");
        state_var_NS <= COMP_LOOP_C_422;
      WHEN COMP_LOOP_C_422 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101000");
        state_var_NS <= COMP_LOOP_C_423;
      WHEN COMP_LOOP_C_423 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101001");
        state_var_NS <= COMP_LOOP_C_424;
      WHEN COMP_LOOP_C_424 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101010");
        state_var_NS <= COMP_LOOP_C_425;
      WHEN COMP_LOOP_C_425 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101011");
        state_var_NS <= COMP_LOOP_C_426;
      WHEN COMP_LOOP_C_426 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101100");
        state_var_NS <= COMP_LOOP_C_427;
      WHEN COMP_LOOP_C_427 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101101");
        state_var_NS <= COMP_LOOP_C_428;
      WHEN COMP_LOOP_C_428 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101110");
        state_var_NS <= COMP_LOOP_C_429;
      WHEN COMP_LOOP_C_429 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101111");
        state_var_NS <= COMP_LOOP_C_430;
      WHEN COMP_LOOP_C_430 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110000");
        state_var_NS <= COMP_LOOP_C_431;
      WHEN COMP_LOOP_C_431 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110001");
        state_var_NS <= COMP_LOOP_C_432;
      WHEN COMP_LOOP_C_432 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110010");
        state_var_NS <= COMP_LOOP_C_433;
      WHEN COMP_LOOP_C_433 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110011");
        state_var_NS <= COMP_LOOP_C_434;
      WHEN COMP_LOOP_C_434 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110100");
        IF ( COMP_LOOP_C_434_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_435;
        END IF;
      WHEN COMP_LOOP_C_435 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_0;
      WHEN COMP_LOOP_8_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_1;
      WHEN COMP_LOOP_8_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_2;
      WHEN COMP_LOOP_8_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_3;
      WHEN COMP_LOOP_8_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_4;
      WHEN COMP_LOOP_8_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_5;
      WHEN COMP_LOOP_8_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_6;
      WHEN COMP_LOOP_8_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_7;
      WHEN COMP_LOOP_8_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_8;
      WHEN COMP_LOOP_8_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_9;
      WHEN COMP_LOOP_8_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_10;
      WHEN COMP_LOOP_8_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_11;
      WHEN COMP_LOOP_8_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_12;
      WHEN COMP_LOOP_8_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_13;
      WHEN COMP_LOOP_8_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_14;
      WHEN COMP_LOOP_8_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_15;
      WHEN COMP_LOOP_8_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_16;
      WHEN COMP_LOOP_8_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_17;
      WHEN COMP_LOOP_8_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_18;
      WHEN COMP_LOOP_8_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_19;
      WHEN COMP_LOOP_8_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_20;
      WHEN COMP_LOOP_8_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_21;
      WHEN COMP_LOOP_8_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_22;
      WHEN COMP_LOOP_8_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_23;
      WHEN COMP_LOOP_8_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_24;
      WHEN COMP_LOOP_8_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_25;
      WHEN COMP_LOOP_8_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_26;
      WHEN COMP_LOOP_8_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_27;
      WHEN COMP_LOOP_8_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_28;
      WHEN COMP_LOOP_8_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_29;
      WHEN COMP_LOOP_8_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_30;
      WHEN COMP_LOOP_8_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010100");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_31;
      WHEN COMP_LOOP_8_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010101");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_32;
      WHEN COMP_LOOP_8_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010110");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_33;
      WHEN COMP_LOOP_8_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010111");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_34;
      WHEN COMP_LOOP_8_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011000");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_35;
      WHEN COMP_LOOP_8_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011001");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_36;
      WHEN COMP_LOOP_8_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011010");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_37;
      WHEN COMP_LOOP_8_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011011");
        state_var_NS <= COMP_LOOP_8_modExp_1_while_C_38;
      WHEN COMP_LOOP_8_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011100");
        IF ( COMP_LOOP_8_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_436;
        ELSE
          state_var_NS <= COMP_LOOP_8_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_436 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011101");
        state_var_NS <= COMP_LOOP_C_437;
      WHEN COMP_LOOP_C_437 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011110");
        state_var_NS <= COMP_LOOP_C_438;
      WHEN COMP_LOOP_C_438 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011111");
        state_var_NS <= COMP_LOOP_C_439;
      WHEN COMP_LOOP_C_439 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100000");
        state_var_NS <= COMP_LOOP_C_440;
      WHEN COMP_LOOP_C_440 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100001");
        state_var_NS <= COMP_LOOP_C_441;
      WHEN COMP_LOOP_C_441 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100010");
        state_var_NS <= COMP_LOOP_C_442;
      WHEN COMP_LOOP_C_442 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100011");
        state_var_NS <= COMP_LOOP_C_443;
      WHEN COMP_LOOP_C_443 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100100");
        state_var_NS <= COMP_LOOP_C_444;
      WHEN COMP_LOOP_C_444 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100101");
        state_var_NS <= COMP_LOOP_C_445;
      WHEN COMP_LOOP_C_445 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100110");
        state_var_NS <= COMP_LOOP_C_446;
      WHEN COMP_LOOP_C_446 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100111");
        state_var_NS <= COMP_LOOP_C_447;
      WHEN COMP_LOOP_C_447 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101000");
        state_var_NS <= COMP_LOOP_C_448;
      WHEN COMP_LOOP_C_448 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101001");
        state_var_NS <= COMP_LOOP_C_449;
      WHEN COMP_LOOP_C_449 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101010");
        state_var_NS <= COMP_LOOP_C_450;
      WHEN COMP_LOOP_C_450 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101011");
        state_var_NS <= COMP_LOOP_C_451;
      WHEN COMP_LOOP_C_451 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101100");
        state_var_NS <= COMP_LOOP_C_452;
      WHEN COMP_LOOP_C_452 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101101");
        state_var_NS <= COMP_LOOP_C_453;
      WHEN COMP_LOOP_C_453 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101110");
        state_var_NS <= COMP_LOOP_C_454;
      WHEN COMP_LOOP_C_454 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101111");
        state_var_NS <= COMP_LOOP_C_455;
      WHEN COMP_LOOP_C_455 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110000");
        state_var_NS <= COMP_LOOP_C_456;
      WHEN COMP_LOOP_C_456 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110001");
        state_var_NS <= COMP_LOOP_C_457;
      WHEN COMP_LOOP_C_457 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110010");
        state_var_NS <= COMP_LOOP_C_458;
      WHEN COMP_LOOP_C_458 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110011");
        state_var_NS <= COMP_LOOP_C_459;
      WHEN COMP_LOOP_C_459 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110100");
        state_var_NS <= COMP_LOOP_C_460;
      WHEN COMP_LOOP_C_460 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110101");
        state_var_NS <= COMP_LOOP_C_461;
      WHEN COMP_LOOP_C_461 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110110");
        state_var_NS <= COMP_LOOP_C_462;
      WHEN COMP_LOOP_C_462 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110111");
        state_var_NS <= COMP_LOOP_C_463;
      WHEN COMP_LOOP_C_463 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111000");
        state_var_NS <= COMP_LOOP_C_464;
      WHEN COMP_LOOP_C_464 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111001");
        state_var_NS <= COMP_LOOP_C_465;
      WHEN COMP_LOOP_C_465 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111010");
        state_var_NS <= COMP_LOOP_C_466;
      WHEN COMP_LOOP_C_466 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111011");
        state_var_NS <= COMP_LOOP_C_467;
      WHEN COMP_LOOP_C_467 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111100");
        state_var_NS <= COMP_LOOP_C_468;
      WHEN COMP_LOOP_C_468 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111101");
        state_var_NS <= COMP_LOOP_C_469;
      WHEN COMP_LOOP_C_469 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111110");
        state_var_NS <= COMP_LOOP_C_470;
      WHEN COMP_LOOP_C_470 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111111");
        state_var_NS <= COMP_LOOP_C_471;
      WHEN COMP_LOOP_C_471 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000000");
        state_var_NS <= COMP_LOOP_C_472;
      WHEN COMP_LOOP_C_472 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000001");
        state_var_NS <= COMP_LOOP_C_473;
      WHEN COMP_LOOP_C_473 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000010");
        state_var_NS <= COMP_LOOP_C_474;
      WHEN COMP_LOOP_C_474 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000011");
        state_var_NS <= COMP_LOOP_C_475;
      WHEN COMP_LOOP_C_475 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000100");
        state_var_NS <= COMP_LOOP_C_476;
      WHEN COMP_LOOP_C_476 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000101");
        state_var_NS <= COMP_LOOP_C_477;
      WHEN COMP_LOOP_C_477 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000110");
        state_var_NS <= COMP_LOOP_C_478;
      WHEN COMP_LOOP_C_478 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000111");
        state_var_NS <= COMP_LOOP_C_479;
      WHEN COMP_LOOP_C_479 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001000");
        state_var_NS <= COMP_LOOP_C_480;
      WHEN COMP_LOOP_C_480 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001001");
        state_var_NS <= COMP_LOOP_C_481;
      WHEN COMP_LOOP_C_481 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001010");
        state_var_NS <= COMP_LOOP_C_482;
      WHEN COMP_LOOP_C_482 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001011");
        state_var_NS <= COMP_LOOP_C_483;
      WHEN COMP_LOOP_C_483 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001100");
        state_var_NS <= COMP_LOOP_C_484;
      WHEN COMP_LOOP_C_484 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001101");
        state_var_NS <= COMP_LOOP_C_485;
      WHEN COMP_LOOP_C_485 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001110");
        state_var_NS <= COMP_LOOP_C_486;
      WHEN COMP_LOOP_C_486 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001111");
        state_var_NS <= COMP_LOOP_C_487;
      WHEN COMP_LOOP_C_487 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010000");
        state_var_NS <= COMP_LOOP_C_488;
      WHEN COMP_LOOP_C_488 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010001");
        state_var_NS <= COMP_LOOP_C_489;
      WHEN COMP_LOOP_C_489 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010010");
        state_var_NS <= COMP_LOOP_C_490;
      WHEN COMP_LOOP_C_490 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010011");
        state_var_NS <= COMP_LOOP_C_491;
      WHEN COMP_LOOP_C_491 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010100");
        state_var_NS <= COMP_LOOP_C_492;
      WHEN COMP_LOOP_C_492 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010101");
        state_var_NS <= COMP_LOOP_C_493;
      WHEN COMP_LOOP_C_493 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010110");
        state_var_NS <= COMP_LOOP_C_494;
      WHEN COMP_LOOP_C_494 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010111");
        state_var_NS <= COMP_LOOP_C_495;
      WHEN COMP_LOOP_C_495 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011000");
        state_var_NS <= COMP_LOOP_C_496;
      WHEN COMP_LOOP_C_496 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011001");
        IF ( COMP_LOOP_C_496_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_497;
        END IF;
      WHEN COMP_LOOP_C_497 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_0;
      WHEN COMP_LOOP_9_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_1;
      WHEN COMP_LOOP_9_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_2;
      WHEN COMP_LOOP_9_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_3;
      WHEN COMP_LOOP_9_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_4;
      WHEN COMP_LOOP_9_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_5;
      WHEN COMP_LOOP_9_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_6;
      WHEN COMP_LOOP_9_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100001");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_7;
      WHEN COMP_LOOP_9_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_8;
      WHEN COMP_LOOP_9_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_9;
      WHEN COMP_LOOP_9_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_10;
      WHEN COMP_LOOP_9_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_11;
      WHEN COMP_LOOP_9_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_12;
      WHEN COMP_LOOP_9_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_13;
      WHEN COMP_LOOP_9_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_14;
      WHEN COMP_LOOP_9_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101001");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_15;
      WHEN COMP_LOOP_9_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_16;
      WHEN COMP_LOOP_9_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_17;
      WHEN COMP_LOOP_9_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_18;
      WHEN COMP_LOOP_9_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_19;
      WHEN COMP_LOOP_9_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_20;
      WHEN COMP_LOOP_9_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_21;
      WHEN COMP_LOOP_9_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_22;
      WHEN COMP_LOOP_9_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110001");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_23;
      WHEN COMP_LOOP_9_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_24;
      WHEN COMP_LOOP_9_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_25;
      WHEN COMP_LOOP_9_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_26;
      WHEN COMP_LOOP_9_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_27;
      WHEN COMP_LOOP_9_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_28;
      WHEN COMP_LOOP_9_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_29;
      WHEN COMP_LOOP_9_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_30;
      WHEN COMP_LOOP_9_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111001");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_31;
      WHEN COMP_LOOP_9_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111010");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_32;
      WHEN COMP_LOOP_9_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111011");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_33;
      WHEN COMP_LOOP_9_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111100");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_34;
      WHEN COMP_LOOP_9_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111101");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_35;
      WHEN COMP_LOOP_9_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111110");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_36;
      WHEN COMP_LOOP_9_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111111");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_37;
      WHEN COMP_LOOP_9_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000000");
        state_var_NS <= COMP_LOOP_9_modExp_1_while_C_38;
      WHEN COMP_LOOP_9_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000001");
        IF ( COMP_LOOP_9_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_498;
        ELSE
          state_var_NS <= COMP_LOOP_9_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_498 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000010");
        state_var_NS <= COMP_LOOP_C_499;
      WHEN COMP_LOOP_C_499 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000011");
        state_var_NS <= COMP_LOOP_C_500;
      WHEN COMP_LOOP_C_500 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000100");
        state_var_NS <= COMP_LOOP_C_501;
      WHEN COMP_LOOP_C_501 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000101");
        state_var_NS <= COMP_LOOP_C_502;
      WHEN COMP_LOOP_C_502 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000110");
        state_var_NS <= COMP_LOOP_C_503;
      WHEN COMP_LOOP_C_503 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000111");
        state_var_NS <= COMP_LOOP_C_504;
      WHEN COMP_LOOP_C_504 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001000");
        state_var_NS <= COMP_LOOP_C_505;
      WHEN COMP_LOOP_C_505 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001001");
        state_var_NS <= COMP_LOOP_C_506;
      WHEN COMP_LOOP_C_506 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001010");
        state_var_NS <= COMP_LOOP_C_507;
      WHEN COMP_LOOP_C_507 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001011");
        state_var_NS <= COMP_LOOP_C_508;
      WHEN COMP_LOOP_C_508 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001100");
        state_var_NS <= COMP_LOOP_C_509;
      WHEN COMP_LOOP_C_509 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001101");
        state_var_NS <= COMP_LOOP_C_510;
      WHEN COMP_LOOP_C_510 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001110");
        state_var_NS <= COMP_LOOP_C_511;
      WHEN COMP_LOOP_C_511 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001111");
        state_var_NS <= COMP_LOOP_C_512;
      WHEN COMP_LOOP_C_512 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010000");
        state_var_NS <= COMP_LOOP_C_513;
      WHEN COMP_LOOP_C_513 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010001");
        state_var_NS <= COMP_LOOP_C_514;
      WHEN COMP_LOOP_C_514 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010010");
        state_var_NS <= COMP_LOOP_C_515;
      WHEN COMP_LOOP_C_515 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010011");
        state_var_NS <= COMP_LOOP_C_516;
      WHEN COMP_LOOP_C_516 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010100");
        state_var_NS <= COMP_LOOP_C_517;
      WHEN COMP_LOOP_C_517 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010101");
        state_var_NS <= COMP_LOOP_C_518;
      WHEN COMP_LOOP_C_518 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010110");
        state_var_NS <= COMP_LOOP_C_519;
      WHEN COMP_LOOP_C_519 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010111");
        state_var_NS <= COMP_LOOP_C_520;
      WHEN COMP_LOOP_C_520 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011000");
        state_var_NS <= COMP_LOOP_C_521;
      WHEN COMP_LOOP_C_521 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011001");
        state_var_NS <= COMP_LOOP_C_522;
      WHEN COMP_LOOP_C_522 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011010");
        state_var_NS <= COMP_LOOP_C_523;
      WHEN COMP_LOOP_C_523 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011011");
        state_var_NS <= COMP_LOOP_C_524;
      WHEN COMP_LOOP_C_524 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011100");
        state_var_NS <= COMP_LOOP_C_525;
      WHEN COMP_LOOP_C_525 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011101");
        state_var_NS <= COMP_LOOP_C_526;
      WHEN COMP_LOOP_C_526 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011110");
        state_var_NS <= COMP_LOOP_C_527;
      WHEN COMP_LOOP_C_527 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011111");
        state_var_NS <= COMP_LOOP_C_528;
      WHEN COMP_LOOP_C_528 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100000");
        state_var_NS <= COMP_LOOP_C_529;
      WHEN COMP_LOOP_C_529 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100001");
        state_var_NS <= COMP_LOOP_C_530;
      WHEN COMP_LOOP_C_530 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100010");
        state_var_NS <= COMP_LOOP_C_531;
      WHEN COMP_LOOP_C_531 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100011");
        state_var_NS <= COMP_LOOP_C_532;
      WHEN COMP_LOOP_C_532 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100100");
        state_var_NS <= COMP_LOOP_C_533;
      WHEN COMP_LOOP_C_533 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100101");
        state_var_NS <= COMP_LOOP_C_534;
      WHEN COMP_LOOP_C_534 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100110");
        state_var_NS <= COMP_LOOP_C_535;
      WHEN COMP_LOOP_C_535 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100111");
        state_var_NS <= COMP_LOOP_C_536;
      WHEN COMP_LOOP_C_536 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101000");
        state_var_NS <= COMP_LOOP_C_537;
      WHEN COMP_LOOP_C_537 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101001");
        state_var_NS <= COMP_LOOP_C_538;
      WHEN COMP_LOOP_C_538 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101010");
        state_var_NS <= COMP_LOOP_C_539;
      WHEN COMP_LOOP_C_539 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101011");
        state_var_NS <= COMP_LOOP_C_540;
      WHEN COMP_LOOP_C_540 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101100");
        state_var_NS <= COMP_LOOP_C_541;
      WHEN COMP_LOOP_C_541 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101101");
        state_var_NS <= COMP_LOOP_C_542;
      WHEN COMP_LOOP_C_542 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101110");
        state_var_NS <= COMP_LOOP_C_543;
      WHEN COMP_LOOP_C_543 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101111");
        state_var_NS <= COMP_LOOP_C_544;
      WHEN COMP_LOOP_C_544 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110000");
        state_var_NS <= COMP_LOOP_C_545;
      WHEN COMP_LOOP_C_545 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110001");
        state_var_NS <= COMP_LOOP_C_546;
      WHEN COMP_LOOP_C_546 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110010");
        state_var_NS <= COMP_LOOP_C_547;
      WHEN COMP_LOOP_C_547 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110011");
        state_var_NS <= COMP_LOOP_C_548;
      WHEN COMP_LOOP_C_548 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110100");
        state_var_NS <= COMP_LOOP_C_549;
      WHEN COMP_LOOP_C_549 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110101");
        state_var_NS <= COMP_LOOP_C_550;
      WHEN COMP_LOOP_C_550 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110110");
        state_var_NS <= COMP_LOOP_C_551;
      WHEN COMP_LOOP_C_551 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110111");
        state_var_NS <= COMP_LOOP_C_552;
      WHEN COMP_LOOP_C_552 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111000");
        state_var_NS <= COMP_LOOP_C_553;
      WHEN COMP_LOOP_C_553 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111001");
        state_var_NS <= COMP_LOOP_C_554;
      WHEN COMP_LOOP_C_554 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111010");
        state_var_NS <= COMP_LOOP_C_555;
      WHEN COMP_LOOP_C_555 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111011");
        state_var_NS <= COMP_LOOP_C_556;
      WHEN COMP_LOOP_C_556 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111100");
        state_var_NS <= COMP_LOOP_C_557;
      WHEN COMP_LOOP_C_557 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111101");
        state_var_NS <= COMP_LOOP_C_558;
      WHEN COMP_LOOP_C_558 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111110");
        IF ( COMP_LOOP_C_558_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_559;
        END IF;
      WHEN COMP_LOOP_C_559 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_0;
      WHEN COMP_LOOP_10_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_1;
      WHEN COMP_LOOP_10_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_2;
      WHEN COMP_LOOP_10_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_3;
      WHEN COMP_LOOP_10_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_4;
      WHEN COMP_LOOP_10_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_5;
      WHEN COMP_LOOP_10_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_6;
      WHEN COMP_LOOP_10_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_7;
      WHEN COMP_LOOP_10_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_8;
      WHEN COMP_LOOP_10_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_9;
      WHEN COMP_LOOP_10_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_10;
      WHEN COMP_LOOP_10_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_11;
      WHEN COMP_LOOP_10_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_12;
      WHEN COMP_LOOP_10_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_13;
      WHEN COMP_LOOP_10_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_14;
      WHEN COMP_LOOP_10_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_15;
      WHEN COMP_LOOP_10_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_16;
      WHEN COMP_LOOP_10_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_17;
      WHEN COMP_LOOP_10_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_18;
      WHEN COMP_LOOP_10_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_19;
      WHEN COMP_LOOP_10_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_20;
      WHEN COMP_LOOP_10_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_21;
      WHEN COMP_LOOP_10_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_22;
      WHEN COMP_LOOP_10_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_23;
      WHEN COMP_LOOP_10_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_24;
      WHEN COMP_LOOP_10_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_25;
      WHEN COMP_LOOP_10_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_26;
      WHEN COMP_LOOP_10_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_27;
      WHEN COMP_LOOP_10_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_28;
      WHEN COMP_LOOP_10_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_29;
      WHEN COMP_LOOP_10_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_30;
      WHEN COMP_LOOP_10_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011110");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_31;
      WHEN COMP_LOOP_10_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011111");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_32;
      WHEN COMP_LOOP_10_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100000");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_33;
      WHEN COMP_LOOP_10_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100001");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_34;
      WHEN COMP_LOOP_10_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100010");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_35;
      WHEN COMP_LOOP_10_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100011");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_36;
      WHEN COMP_LOOP_10_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100100");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_37;
      WHEN COMP_LOOP_10_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100101");
        state_var_NS <= COMP_LOOP_10_modExp_1_while_C_38;
      WHEN COMP_LOOP_10_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100110");
        IF ( COMP_LOOP_10_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_560;
        ELSE
          state_var_NS <= COMP_LOOP_10_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_560 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100111");
        state_var_NS <= COMP_LOOP_C_561;
      WHEN COMP_LOOP_C_561 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101000");
        state_var_NS <= COMP_LOOP_C_562;
      WHEN COMP_LOOP_C_562 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101001");
        state_var_NS <= COMP_LOOP_C_563;
      WHEN COMP_LOOP_C_563 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101010");
        state_var_NS <= COMP_LOOP_C_564;
      WHEN COMP_LOOP_C_564 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101011");
        state_var_NS <= COMP_LOOP_C_565;
      WHEN COMP_LOOP_C_565 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101100");
        state_var_NS <= COMP_LOOP_C_566;
      WHEN COMP_LOOP_C_566 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101101");
        state_var_NS <= COMP_LOOP_C_567;
      WHEN COMP_LOOP_C_567 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101110");
        state_var_NS <= COMP_LOOP_C_568;
      WHEN COMP_LOOP_C_568 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101111");
        state_var_NS <= COMP_LOOP_C_569;
      WHEN COMP_LOOP_C_569 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110000");
        state_var_NS <= COMP_LOOP_C_570;
      WHEN COMP_LOOP_C_570 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110001");
        state_var_NS <= COMP_LOOP_C_571;
      WHEN COMP_LOOP_C_571 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110010");
        state_var_NS <= COMP_LOOP_C_572;
      WHEN COMP_LOOP_C_572 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110011");
        state_var_NS <= COMP_LOOP_C_573;
      WHEN COMP_LOOP_C_573 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110100");
        state_var_NS <= COMP_LOOP_C_574;
      WHEN COMP_LOOP_C_574 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110101");
        state_var_NS <= COMP_LOOP_C_575;
      WHEN COMP_LOOP_C_575 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110110");
        state_var_NS <= COMP_LOOP_C_576;
      WHEN COMP_LOOP_C_576 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110111");
        state_var_NS <= COMP_LOOP_C_577;
      WHEN COMP_LOOP_C_577 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111000");
        state_var_NS <= COMP_LOOP_C_578;
      WHEN COMP_LOOP_C_578 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111001");
        state_var_NS <= COMP_LOOP_C_579;
      WHEN COMP_LOOP_C_579 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111010");
        state_var_NS <= COMP_LOOP_C_580;
      WHEN COMP_LOOP_C_580 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111011");
        state_var_NS <= COMP_LOOP_C_581;
      WHEN COMP_LOOP_C_581 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111100");
        state_var_NS <= COMP_LOOP_C_582;
      WHEN COMP_LOOP_C_582 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111101");
        state_var_NS <= COMP_LOOP_C_583;
      WHEN COMP_LOOP_C_583 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111110");
        state_var_NS <= COMP_LOOP_C_584;
      WHEN COMP_LOOP_C_584 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111111");
        state_var_NS <= COMP_LOOP_C_585;
      WHEN COMP_LOOP_C_585 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000000");
        state_var_NS <= COMP_LOOP_C_586;
      WHEN COMP_LOOP_C_586 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000001");
        state_var_NS <= COMP_LOOP_C_587;
      WHEN COMP_LOOP_C_587 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000010");
        state_var_NS <= COMP_LOOP_C_588;
      WHEN COMP_LOOP_C_588 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000011");
        state_var_NS <= COMP_LOOP_C_589;
      WHEN COMP_LOOP_C_589 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000100");
        state_var_NS <= COMP_LOOP_C_590;
      WHEN COMP_LOOP_C_590 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000101");
        state_var_NS <= COMP_LOOP_C_591;
      WHEN COMP_LOOP_C_591 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000110");
        state_var_NS <= COMP_LOOP_C_592;
      WHEN COMP_LOOP_C_592 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000111");
        state_var_NS <= COMP_LOOP_C_593;
      WHEN COMP_LOOP_C_593 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001000");
        state_var_NS <= COMP_LOOP_C_594;
      WHEN COMP_LOOP_C_594 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001001");
        state_var_NS <= COMP_LOOP_C_595;
      WHEN COMP_LOOP_C_595 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001010");
        state_var_NS <= COMP_LOOP_C_596;
      WHEN COMP_LOOP_C_596 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001011");
        state_var_NS <= COMP_LOOP_C_597;
      WHEN COMP_LOOP_C_597 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001100");
        state_var_NS <= COMP_LOOP_C_598;
      WHEN COMP_LOOP_C_598 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001101");
        state_var_NS <= COMP_LOOP_C_599;
      WHEN COMP_LOOP_C_599 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001110");
        state_var_NS <= COMP_LOOP_C_600;
      WHEN COMP_LOOP_C_600 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001111");
        state_var_NS <= COMP_LOOP_C_601;
      WHEN COMP_LOOP_C_601 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010000");
        state_var_NS <= COMP_LOOP_C_602;
      WHEN COMP_LOOP_C_602 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010001");
        state_var_NS <= COMP_LOOP_C_603;
      WHEN COMP_LOOP_C_603 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010010");
        state_var_NS <= COMP_LOOP_C_604;
      WHEN COMP_LOOP_C_604 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010011");
        state_var_NS <= COMP_LOOP_C_605;
      WHEN COMP_LOOP_C_605 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010100");
        state_var_NS <= COMP_LOOP_C_606;
      WHEN COMP_LOOP_C_606 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010101");
        state_var_NS <= COMP_LOOP_C_607;
      WHEN COMP_LOOP_C_607 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010110");
        state_var_NS <= COMP_LOOP_C_608;
      WHEN COMP_LOOP_C_608 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010111");
        state_var_NS <= COMP_LOOP_C_609;
      WHEN COMP_LOOP_C_609 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011000");
        state_var_NS <= COMP_LOOP_C_610;
      WHEN COMP_LOOP_C_610 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011001");
        state_var_NS <= COMP_LOOP_C_611;
      WHEN COMP_LOOP_C_611 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011010");
        state_var_NS <= COMP_LOOP_C_612;
      WHEN COMP_LOOP_C_612 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011011");
        state_var_NS <= COMP_LOOP_C_613;
      WHEN COMP_LOOP_C_613 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011100");
        state_var_NS <= COMP_LOOP_C_614;
      WHEN COMP_LOOP_C_614 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011101");
        state_var_NS <= COMP_LOOP_C_615;
      WHEN COMP_LOOP_C_615 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011110");
        state_var_NS <= COMP_LOOP_C_616;
      WHEN COMP_LOOP_C_616 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011111");
        state_var_NS <= COMP_LOOP_C_617;
      WHEN COMP_LOOP_C_617 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100000");
        state_var_NS <= COMP_LOOP_C_618;
      WHEN COMP_LOOP_C_618 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100001");
        state_var_NS <= COMP_LOOP_C_619;
      WHEN COMP_LOOP_C_619 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100010");
        state_var_NS <= COMP_LOOP_C_620;
      WHEN COMP_LOOP_C_620 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100011");
        IF ( COMP_LOOP_C_620_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_621;
        END IF;
      WHEN COMP_LOOP_C_621 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_0;
      WHEN COMP_LOOP_11_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_1;
      WHEN COMP_LOOP_11_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_2;
      WHEN COMP_LOOP_11_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_3;
      WHEN COMP_LOOP_11_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_4;
      WHEN COMP_LOOP_11_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_5;
      WHEN COMP_LOOP_11_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_6;
      WHEN COMP_LOOP_11_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_7;
      WHEN COMP_LOOP_11_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_8;
      WHEN COMP_LOOP_11_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_9;
      WHEN COMP_LOOP_11_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_10;
      WHEN COMP_LOOP_11_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_11;
      WHEN COMP_LOOP_11_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_12;
      WHEN COMP_LOOP_11_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_13;
      WHEN COMP_LOOP_11_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_14;
      WHEN COMP_LOOP_11_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_15;
      WHEN COMP_LOOP_11_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_16;
      WHEN COMP_LOOP_11_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_17;
      WHEN COMP_LOOP_11_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_18;
      WHEN COMP_LOOP_11_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_19;
      WHEN COMP_LOOP_11_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_20;
      WHEN COMP_LOOP_11_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_21;
      WHEN COMP_LOOP_11_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_22;
      WHEN COMP_LOOP_11_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_23;
      WHEN COMP_LOOP_11_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_24;
      WHEN COMP_LOOP_11_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_25;
      WHEN COMP_LOOP_11_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_26;
      WHEN COMP_LOOP_11_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_27;
      WHEN COMP_LOOP_11_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_28;
      WHEN COMP_LOOP_11_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_29;
      WHEN COMP_LOOP_11_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_30;
      WHEN COMP_LOOP_11_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000011");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_31;
      WHEN COMP_LOOP_11_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000100");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_32;
      WHEN COMP_LOOP_11_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000101");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_33;
      WHEN COMP_LOOP_11_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000110");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_34;
      WHEN COMP_LOOP_11_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000111");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_35;
      WHEN COMP_LOOP_11_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001000");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_36;
      WHEN COMP_LOOP_11_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001001");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_37;
      WHEN COMP_LOOP_11_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001010");
        state_var_NS <= COMP_LOOP_11_modExp_1_while_C_38;
      WHEN COMP_LOOP_11_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001011");
        IF ( COMP_LOOP_11_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_622;
        ELSE
          state_var_NS <= COMP_LOOP_11_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_622 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001100");
        state_var_NS <= COMP_LOOP_C_623;
      WHEN COMP_LOOP_C_623 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001101");
        state_var_NS <= COMP_LOOP_C_624;
      WHEN COMP_LOOP_C_624 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001110");
        state_var_NS <= COMP_LOOP_C_625;
      WHEN COMP_LOOP_C_625 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001111");
        state_var_NS <= COMP_LOOP_C_626;
      WHEN COMP_LOOP_C_626 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010000");
        state_var_NS <= COMP_LOOP_C_627;
      WHEN COMP_LOOP_C_627 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010001");
        state_var_NS <= COMP_LOOP_C_628;
      WHEN COMP_LOOP_C_628 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010010");
        state_var_NS <= COMP_LOOP_C_629;
      WHEN COMP_LOOP_C_629 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010011");
        state_var_NS <= COMP_LOOP_C_630;
      WHEN COMP_LOOP_C_630 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010100");
        state_var_NS <= COMP_LOOP_C_631;
      WHEN COMP_LOOP_C_631 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010101");
        state_var_NS <= COMP_LOOP_C_632;
      WHEN COMP_LOOP_C_632 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010110");
        state_var_NS <= COMP_LOOP_C_633;
      WHEN COMP_LOOP_C_633 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010111");
        state_var_NS <= COMP_LOOP_C_634;
      WHEN COMP_LOOP_C_634 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011000");
        state_var_NS <= COMP_LOOP_C_635;
      WHEN COMP_LOOP_C_635 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011001");
        state_var_NS <= COMP_LOOP_C_636;
      WHEN COMP_LOOP_C_636 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011010");
        state_var_NS <= COMP_LOOP_C_637;
      WHEN COMP_LOOP_C_637 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011011");
        state_var_NS <= COMP_LOOP_C_638;
      WHEN COMP_LOOP_C_638 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011100");
        state_var_NS <= COMP_LOOP_C_639;
      WHEN COMP_LOOP_C_639 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011101");
        state_var_NS <= COMP_LOOP_C_640;
      WHEN COMP_LOOP_C_640 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011110");
        state_var_NS <= COMP_LOOP_C_641;
      WHEN COMP_LOOP_C_641 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011111");
        state_var_NS <= COMP_LOOP_C_642;
      WHEN COMP_LOOP_C_642 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100000");
        state_var_NS <= COMP_LOOP_C_643;
      WHEN COMP_LOOP_C_643 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100001");
        state_var_NS <= COMP_LOOP_C_644;
      WHEN COMP_LOOP_C_644 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100010");
        state_var_NS <= COMP_LOOP_C_645;
      WHEN COMP_LOOP_C_645 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100011");
        state_var_NS <= COMP_LOOP_C_646;
      WHEN COMP_LOOP_C_646 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100100");
        state_var_NS <= COMP_LOOP_C_647;
      WHEN COMP_LOOP_C_647 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100101");
        state_var_NS <= COMP_LOOP_C_648;
      WHEN COMP_LOOP_C_648 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100110");
        state_var_NS <= COMP_LOOP_C_649;
      WHEN COMP_LOOP_C_649 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100111");
        state_var_NS <= COMP_LOOP_C_650;
      WHEN COMP_LOOP_C_650 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101000");
        state_var_NS <= COMP_LOOP_C_651;
      WHEN COMP_LOOP_C_651 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101001");
        state_var_NS <= COMP_LOOP_C_652;
      WHEN COMP_LOOP_C_652 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101010");
        state_var_NS <= COMP_LOOP_C_653;
      WHEN COMP_LOOP_C_653 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101011");
        state_var_NS <= COMP_LOOP_C_654;
      WHEN COMP_LOOP_C_654 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101100");
        state_var_NS <= COMP_LOOP_C_655;
      WHEN COMP_LOOP_C_655 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101101");
        state_var_NS <= COMP_LOOP_C_656;
      WHEN COMP_LOOP_C_656 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101110");
        state_var_NS <= COMP_LOOP_C_657;
      WHEN COMP_LOOP_C_657 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101111");
        state_var_NS <= COMP_LOOP_C_658;
      WHEN COMP_LOOP_C_658 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110000");
        state_var_NS <= COMP_LOOP_C_659;
      WHEN COMP_LOOP_C_659 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110001");
        state_var_NS <= COMP_LOOP_C_660;
      WHEN COMP_LOOP_C_660 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110010");
        state_var_NS <= COMP_LOOP_C_661;
      WHEN COMP_LOOP_C_661 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110011");
        state_var_NS <= COMP_LOOP_C_662;
      WHEN COMP_LOOP_C_662 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110100");
        state_var_NS <= COMP_LOOP_C_663;
      WHEN COMP_LOOP_C_663 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110101");
        state_var_NS <= COMP_LOOP_C_664;
      WHEN COMP_LOOP_C_664 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110110");
        state_var_NS <= COMP_LOOP_C_665;
      WHEN COMP_LOOP_C_665 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110111");
        state_var_NS <= COMP_LOOP_C_666;
      WHEN COMP_LOOP_C_666 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111000");
        state_var_NS <= COMP_LOOP_C_667;
      WHEN COMP_LOOP_C_667 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111001");
        state_var_NS <= COMP_LOOP_C_668;
      WHEN COMP_LOOP_C_668 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111010");
        state_var_NS <= COMP_LOOP_C_669;
      WHEN COMP_LOOP_C_669 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111011");
        state_var_NS <= COMP_LOOP_C_670;
      WHEN COMP_LOOP_C_670 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111100");
        state_var_NS <= COMP_LOOP_C_671;
      WHEN COMP_LOOP_C_671 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111101");
        state_var_NS <= COMP_LOOP_C_672;
      WHEN COMP_LOOP_C_672 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111110");
        state_var_NS <= COMP_LOOP_C_673;
      WHEN COMP_LOOP_C_673 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111111");
        state_var_NS <= COMP_LOOP_C_674;
      WHEN COMP_LOOP_C_674 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000000");
        state_var_NS <= COMP_LOOP_C_675;
      WHEN COMP_LOOP_C_675 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000001");
        state_var_NS <= COMP_LOOP_C_676;
      WHEN COMP_LOOP_C_676 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000010");
        state_var_NS <= COMP_LOOP_C_677;
      WHEN COMP_LOOP_C_677 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000011");
        state_var_NS <= COMP_LOOP_C_678;
      WHEN COMP_LOOP_C_678 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000100");
        state_var_NS <= COMP_LOOP_C_679;
      WHEN COMP_LOOP_C_679 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000101");
        state_var_NS <= COMP_LOOP_C_680;
      WHEN COMP_LOOP_C_680 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000110");
        state_var_NS <= COMP_LOOP_C_681;
      WHEN COMP_LOOP_C_681 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000111");
        state_var_NS <= COMP_LOOP_C_682;
      WHEN COMP_LOOP_C_682 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001000");
        IF ( COMP_LOOP_C_682_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_683;
        END IF;
      WHEN COMP_LOOP_C_683 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_0;
      WHEN COMP_LOOP_12_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_1;
      WHEN COMP_LOOP_12_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_2;
      WHEN COMP_LOOP_12_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_3;
      WHEN COMP_LOOP_12_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_4;
      WHEN COMP_LOOP_12_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_5;
      WHEN COMP_LOOP_12_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_6;
      WHEN COMP_LOOP_12_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_7;
      WHEN COMP_LOOP_12_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_8;
      WHEN COMP_LOOP_12_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_9;
      WHEN COMP_LOOP_12_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_10;
      WHEN COMP_LOOP_12_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_11;
      WHEN COMP_LOOP_12_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_12;
      WHEN COMP_LOOP_12_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_13;
      WHEN COMP_LOOP_12_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_14;
      WHEN COMP_LOOP_12_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_15;
      WHEN COMP_LOOP_12_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_16;
      WHEN COMP_LOOP_12_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_17;
      WHEN COMP_LOOP_12_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_18;
      WHEN COMP_LOOP_12_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_19;
      WHEN COMP_LOOP_12_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_20;
      WHEN COMP_LOOP_12_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_21;
      WHEN COMP_LOOP_12_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_22;
      WHEN COMP_LOOP_12_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_23;
      WHEN COMP_LOOP_12_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_24;
      WHEN COMP_LOOP_12_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_25;
      WHEN COMP_LOOP_12_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_26;
      WHEN COMP_LOOP_12_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_27;
      WHEN COMP_LOOP_12_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_28;
      WHEN COMP_LOOP_12_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_29;
      WHEN COMP_LOOP_12_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_30;
      WHEN COMP_LOOP_12_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101000");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_31;
      WHEN COMP_LOOP_12_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101001");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_32;
      WHEN COMP_LOOP_12_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101010");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_33;
      WHEN COMP_LOOP_12_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101011");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_34;
      WHEN COMP_LOOP_12_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101100");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_35;
      WHEN COMP_LOOP_12_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101101");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_36;
      WHEN COMP_LOOP_12_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101110");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_37;
      WHEN COMP_LOOP_12_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101111");
        state_var_NS <= COMP_LOOP_12_modExp_1_while_C_38;
      WHEN COMP_LOOP_12_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110000");
        IF ( COMP_LOOP_12_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_684;
        ELSE
          state_var_NS <= COMP_LOOP_12_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_684 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110001");
        state_var_NS <= COMP_LOOP_C_685;
      WHEN COMP_LOOP_C_685 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110010");
        state_var_NS <= COMP_LOOP_C_686;
      WHEN COMP_LOOP_C_686 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110011");
        state_var_NS <= COMP_LOOP_C_687;
      WHEN COMP_LOOP_C_687 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110100");
        state_var_NS <= COMP_LOOP_C_688;
      WHEN COMP_LOOP_C_688 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110101");
        state_var_NS <= COMP_LOOP_C_689;
      WHEN COMP_LOOP_C_689 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110110");
        state_var_NS <= COMP_LOOP_C_690;
      WHEN COMP_LOOP_C_690 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110111");
        state_var_NS <= COMP_LOOP_C_691;
      WHEN COMP_LOOP_C_691 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111000");
        state_var_NS <= COMP_LOOP_C_692;
      WHEN COMP_LOOP_C_692 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111001");
        state_var_NS <= COMP_LOOP_C_693;
      WHEN COMP_LOOP_C_693 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111010");
        state_var_NS <= COMP_LOOP_C_694;
      WHEN COMP_LOOP_C_694 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111011");
        state_var_NS <= COMP_LOOP_C_695;
      WHEN COMP_LOOP_C_695 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111100");
        state_var_NS <= COMP_LOOP_C_696;
      WHEN COMP_LOOP_C_696 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111101");
        state_var_NS <= COMP_LOOP_C_697;
      WHEN COMP_LOOP_C_697 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111110");
        state_var_NS <= COMP_LOOP_C_698;
      WHEN COMP_LOOP_C_698 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111111");
        state_var_NS <= COMP_LOOP_C_699;
      WHEN COMP_LOOP_C_699 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000000");
        state_var_NS <= COMP_LOOP_C_700;
      WHEN COMP_LOOP_C_700 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000001");
        state_var_NS <= COMP_LOOP_C_701;
      WHEN COMP_LOOP_C_701 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000010");
        state_var_NS <= COMP_LOOP_C_702;
      WHEN COMP_LOOP_C_702 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000011");
        state_var_NS <= COMP_LOOP_C_703;
      WHEN COMP_LOOP_C_703 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000100");
        state_var_NS <= COMP_LOOP_C_704;
      WHEN COMP_LOOP_C_704 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000101");
        state_var_NS <= COMP_LOOP_C_705;
      WHEN COMP_LOOP_C_705 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000110");
        state_var_NS <= COMP_LOOP_C_706;
      WHEN COMP_LOOP_C_706 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000111");
        state_var_NS <= COMP_LOOP_C_707;
      WHEN COMP_LOOP_C_707 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001000");
        state_var_NS <= COMP_LOOP_C_708;
      WHEN COMP_LOOP_C_708 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001001");
        state_var_NS <= COMP_LOOP_C_709;
      WHEN COMP_LOOP_C_709 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001010");
        state_var_NS <= COMP_LOOP_C_710;
      WHEN COMP_LOOP_C_710 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001011");
        state_var_NS <= COMP_LOOP_C_711;
      WHEN COMP_LOOP_C_711 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001100");
        state_var_NS <= COMP_LOOP_C_712;
      WHEN COMP_LOOP_C_712 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001101");
        state_var_NS <= COMP_LOOP_C_713;
      WHEN COMP_LOOP_C_713 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001110");
        state_var_NS <= COMP_LOOP_C_714;
      WHEN COMP_LOOP_C_714 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001111");
        state_var_NS <= COMP_LOOP_C_715;
      WHEN COMP_LOOP_C_715 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010000");
        state_var_NS <= COMP_LOOP_C_716;
      WHEN COMP_LOOP_C_716 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010001");
        state_var_NS <= COMP_LOOP_C_717;
      WHEN COMP_LOOP_C_717 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010010");
        state_var_NS <= COMP_LOOP_C_718;
      WHEN COMP_LOOP_C_718 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010011");
        state_var_NS <= COMP_LOOP_C_719;
      WHEN COMP_LOOP_C_719 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010100");
        state_var_NS <= COMP_LOOP_C_720;
      WHEN COMP_LOOP_C_720 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010101");
        state_var_NS <= COMP_LOOP_C_721;
      WHEN COMP_LOOP_C_721 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010110");
        state_var_NS <= COMP_LOOP_C_722;
      WHEN COMP_LOOP_C_722 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010111");
        state_var_NS <= COMP_LOOP_C_723;
      WHEN COMP_LOOP_C_723 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011000");
        state_var_NS <= COMP_LOOP_C_724;
      WHEN COMP_LOOP_C_724 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011001");
        state_var_NS <= COMP_LOOP_C_725;
      WHEN COMP_LOOP_C_725 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011010");
        state_var_NS <= COMP_LOOP_C_726;
      WHEN COMP_LOOP_C_726 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011011");
        state_var_NS <= COMP_LOOP_C_727;
      WHEN COMP_LOOP_C_727 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011100");
        state_var_NS <= COMP_LOOP_C_728;
      WHEN COMP_LOOP_C_728 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011101");
        state_var_NS <= COMP_LOOP_C_729;
      WHEN COMP_LOOP_C_729 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011110");
        state_var_NS <= COMP_LOOP_C_730;
      WHEN COMP_LOOP_C_730 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011111");
        state_var_NS <= COMP_LOOP_C_731;
      WHEN COMP_LOOP_C_731 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100000");
        state_var_NS <= COMP_LOOP_C_732;
      WHEN COMP_LOOP_C_732 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100001");
        state_var_NS <= COMP_LOOP_C_733;
      WHEN COMP_LOOP_C_733 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100010");
        state_var_NS <= COMP_LOOP_C_734;
      WHEN COMP_LOOP_C_734 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100011");
        state_var_NS <= COMP_LOOP_C_735;
      WHEN COMP_LOOP_C_735 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100100");
        state_var_NS <= COMP_LOOP_C_736;
      WHEN COMP_LOOP_C_736 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100101");
        state_var_NS <= COMP_LOOP_C_737;
      WHEN COMP_LOOP_C_737 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100110");
        state_var_NS <= COMP_LOOP_C_738;
      WHEN COMP_LOOP_C_738 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100111");
        state_var_NS <= COMP_LOOP_C_739;
      WHEN COMP_LOOP_C_739 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101000");
        state_var_NS <= COMP_LOOP_C_740;
      WHEN COMP_LOOP_C_740 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101001");
        state_var_NS <= COMP_LOOP_C_741;
      WHEN COMP_LOOP_C_741 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101010");
        state_var_NS <= COMP_LOOP_C_742;
      WHEN COMP_LOOP_C_742 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101011");
        state_var_NS <= COMP_LOOP_C_743;
      WHEN COMP_LOOP_C_743 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101100");
        state_var_NS <= COMP_LOOP_C_744;
      WHEN COMP_LOOP_C_744 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101101");
        IF ( COMP_LOOP_C_744_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_745;
        END IF;
      WHEN COMP_LOOP_C_745 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_0;
      WHEN COMP_LOOP_13_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_1;
      WHEN COMP_LOOP_13_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_2;
      WHEN COMP_LOOP_13_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_3;
      WHEN COMP_LOOP_13_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_4;
      WHEN COMP_LOOP_13_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_5;
      WHEN COMP_LOOP_13_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_6;
      WHEN COMP_LOOP_13_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110101");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_7;
      WHEN COMP_LOOP_13_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_8;
      WHEN COMP_LOOP_13_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_9;
      WHEN COMP_LOOP_13_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_10;
      WHEN COMP_LOOP_13_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_11;
      WHEN COMP_LOOP_13_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_12;
      WHEN COMP_LOOP_13_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_13;
      WHEN COMP_LOOP_13_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_14;
      WHEN COMP_LOOP_13_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111101");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_15;
      WHEN COMP_LOOP_13_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_16;
      WHEN COMP_LOOP_13_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_17;
      WHEN COMP_LOOP_13_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_18;
      WHEN COMP_LOOP_13_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_19;
      WHEN COMP_LOOP_13_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_20;
      WHEN COMP_LOOP_13_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_21;
      WHEN COMP_LOOP_13_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_22;
      WHEN COMP_LOOP_13_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000101");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_23;
      WHEN COMP_LOOP_13_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_24;
      WHEN COMP_LOOP_13_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_25;
      WHEN COMP_LOOP_13_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_26;
      WHEN COMP_LOOP_13_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_27;
      WHEN COMP_LOOP_13_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_28;
      WHEN COMP_LOOP_13_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_29;
      WHEN COMP_LOOP_13_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_30;
      WHEN COMP_LOOP_13_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001101");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_31;
      WHEN COMP_LOOP_13_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001110");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_32;
      WHEN COMP_LOOP_13_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001111");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_33;
      WHEN COMP_LOOP_13_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010000");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_34;
      WHEN COMP_LOOP_13_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010001");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_35;
      WHEN COMP_LOOP_13_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010010");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_36;
      WHEN COMP_LOOP_13_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010011");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_37;
      WHEN COMP_LOOP_13_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010100");
        state_var_NS <= COMP_LOOP_13_modExp_1_while_C_38;
      WHEN COMP_LOOP_13_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010101");
        IF ( COMP_LOOP_13_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_746;
        ELSE
          state_var_NS <= COMP_LOOP_13_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_746 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010110");
        state_var_NS <= COMP_LOOP_C_747;
      WHEN COMP_LOOP_C_747 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010111");
        state_var_NS <= COMP_LOOP_C_748;
      WHEN COMP_LOOP_C_748 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011000");
        state_var_NS <= COMP_LOOP_C_749;
      WHEN COMP_LOOP_C_749 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011001");
        state_var_NS <= COMP_LOOP_C_750;
      WHEN COMP_LOOP_C_750 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011010");
        state_var_NS <= COMP_LOOP_C_751;
      WHEN COMP_LOOP_C_751 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011011");
        state_var_NS <= COMP_LOOP_C_752;
      WHEN COMP_LOOP_C_752 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011100");
        state_var_NS <= COMP_LOOP_C_753;
      WHEN COMP_LOOP_C_753 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011101");
        state_var_NS <= COMP_LOOP_C_754;
      WHEN COMP_LOOP_C_754 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011110");
        state_var_NS <= COMP_LOOP_C_755;
      WHEN COMP_LOOP_C_755 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011111");
        state_var_NS <= COMP_LOOP_C_756;
      WHEN COMP_LOOP_C_756 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100000");
        state_var_NS <= COMP_LOOP_C_757;
      WHEN COMP_LOOP_C_757 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100001");
        state_var_NS <= COMP_LOOP_C_758;
      WHEN COMP_LOOP_C_758 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100010");
        state_var_NS <= COMP_LOOP_C_759;
      WHEN COMP_LOOP_C_759 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100011");
        state_var_NS <= COMP_LOOP_C_760;
      WHEN COMP_LOOP_C_760 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100100");
        state_var_NS <= COMP_LOOP_C_761;
      WHEN COMP_LOOP_C_761 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100101");
        state_var_NS <= COMP_LOOP_C_762;
      WHEN COMP_LOOP_C_762 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100110");
        state_var_NS <= COMP_LOOP_C_763;
      WHEN COMP_LOOP_C_763 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100111");
        state_var_NS <= COMP_LOOP_C_764;
      WHEN COMP_LOOP_C_764 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101000");
        state_var_NS <= COMP_LOOP_C_765;
      WHEN COMP_LOOP_C_765 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101001");
        state_var_NS <= COMP_LOOP_C_766;
      WHEN COMP_LOOP_C_766 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101010");
        state_var_NS <= COMP_LOOP_C_767;
      WHEN COMP_LOOP_C_767 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101011");
        state_var_NS <= COMP_LOOP_C_768;
      WHEN COMP_LOOP_C_768 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101100");
        state_var_NS <= COMP_LOOP_C_769;
      WHEN COMP_LOOP_C_769 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101101");
        state_var_NS <= COMP_LOOP_C_770;
      WHEN COMP_LOOP_C_770 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101110");
        state_var_NS <= COMP_LOOP_C_771;
      WHEN COMP_LOOP_C_771 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101111");
        state_var_NS <= COMP_LOOP_C_772;
      WHEN COMP_LOOP_C_772 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110000");
        state_var_NS <= COMP_LOOP_C_773;
      WHEN COMP_LOOP_C_773 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110001");
        state_var_NS <= COMP_LOOP_C_774;
      WHEN COMP_LOOP_C_774 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110010");
        state_var_NS <= COMP_LOOP_C_775;
      WHEN COMP_LOOP_C_775 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110011");
        state_var_NS <= COMP_LOOP_C_776;
      WHEN COMP_LOOP_C_776 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110100");
        state_var_NS <= COMP_LOOP_C_777;
      WHEN COMP_LOOP_C_777 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110101");
        state_var_NS <= COMP_LOOP_C_778;
      WHEN COMP_LOOP_C_778 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110110");
        state_var_NS <= COMP_LOOP_C_779;
      WHEN COMP_LOOP_C_779 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110111");
        state_var_NS <= COMP_LOOP_C_780;
      WHEN COMP_LOOP_C_780 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111000");
        state_var_NS <= COMP_LOOP_C_781;
      WHEN COMP_LOOP_C_781 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111001");
        state_var_NS <= COMP_LOOP_C_782;
      WHEN COMP_LOOP_C_782 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111010");
        state_var_NS <= COMP_LOOP_C_783;
      WHEN COMP_LOOP_C_783 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111011");
        state_var_NS <= COMP_LOOP_C_784;
      WHEN COMP_LOOP_C_784 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111100");
        state_var_NS <= COMP_LOOP_C_785;
      WHEN COMP_LOOP_C_785 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111101");
        state_var_NS <= COMP_LOOP_C_786;
      WHEN COMP_LOOP_C_786 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111110");
        state_var_NS <= COMP_LOOP_C_787;
      WHEN COMP_LOOP_C_787 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111111");
        state_var_NS <= COMP_LOOP_C_788;
      WHEN COMP_LOOP_C_788 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000000");
        state_var_NS <= COMP_LOOP_C_789;
      WHEN COMP_LOOP_C_789 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000001");
        state_var_NS <= COMP_LOOP_C_790;
      WHEN COMP_LOOP_C_790 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000010");
        state_var_NS <= COMP_LOOP_C_791;
      WHEN COMP_LOOP_C_791 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000011");
        state_var_NS <= COMP_LOOP_C_792;
      WHEN COMP_LOOP_C_792 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000100");
        state_var_NS <= COMP_LOOP_C_793;
      WHEN COMP_LOOP_C_793 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000101");
        state_var_NS <= COMP_LOOP_C_794;
      WHEN COMP_LOOP_C_794 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000110");
        state_var_NS <= COMP_LOOP_C_795;
      WHEN COMP_LOOP_C_795 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000111");
        state_var_NS <= COMP_LOOP_C_796;
      WHEN COMP_LOOP_C_796 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001000");
        state_var_NS <= COMP_LOOP_C_797;
      WHEN COMP_LOOP_C_797 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001001");
        state_var_NS <= COMP_LOOP_C_798;
      WHEN COMP_LOOP_C_798 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001010");
        state_var_NS <= COMP_LOOP_C_799;
      WHEN COMP_LOOP_C_799 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001011");
        state_var_NS <= COMP_LOOP_C_800;
      WHEN COMP_LOOP_C_800 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001100");
        state_var_NS <= COMP_LOOP_C_801;
      WHEN COMP_LOOP_C_801 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001101");
        state_var_NS <= COMP_LOOP_C_802;
      WHEN COMP_LOOP_C_802 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001110");
        state_var_NS <= COMP_LOOP_C_803;
      WHEN COMP_LOOP_C_803 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001111");
        state_var_NS <= COMP_LOOP_C_804;
      WHEN COMP_LOOP_C_804 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010000");
        state_var_NS <= COMP_LOOP_C_805;
      WHEN COMP_LOOP_C_805 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010001");
        state_var_NS <= COMP_LOOP_C_806;
      WHEN COMP_LOOP_C_806 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010010");
        IF ( COMP_LOOP_C_806_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_807;
        END IF;
      WHEN COMP_LOOP_C_807 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_0;
      WHEN COMP_LOOP_14_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_1;
      WHEN COMP_LOOP_14_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_2;
      WHEN COMP_LOOP_14_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_3;
      WHEN COMP_LOOP_14_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_4;
      WHEN COMP_LOOP_14_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_5;
      WHEN COMP_LOOP_14_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_6;
      WHEN COMP_LOOP_14_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_7;
      WHEN COMP_LOOP_14_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_8;
      WHEN COMP_LOOP_14_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_9;
      WHEN COMP_LOOP_14_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_10;
      WHEN COMP_LOOP_14_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_11;
      WHEN COMP_LOOP_14_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_12;
      WHEN COMP_LOOP_14_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_13;
      WHEN COMP_LOOP_14_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_14;
      WHEN COMP_LOOP_14_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_15;
      WHEN COMP_LOOP_14_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_16;
      WHEN COMP_LOOP_14_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_17;
      WHEN COMP_LOOP_14_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_18;
      WHEN COMP_LOOP_14_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_19;
      WHEN COMP_LOOP_14_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_20;
      WHEN COMP_LOOP_14_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_21;
      WHEN COMP_LOOP_14_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_22;
      WHEN COMP_LOOP_14_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_23;
      WHEN COMP_LOOP_14_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_24;
      WHEN COMP_LOOP_14_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_25;
      WHEN COMP_LOOP_14_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_26;
      WHEN COMP_LOOP_14_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_27;
      WHEN COMP_LOOP_14_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_28;
      WHEN COMP_LOOP_14_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_29;
      WHEN COMP_LOOP_14_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_30;
      WHEN COMP_LOOP_14_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110010");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_31;
      WHEN COMP_LOOP_14_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110011");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_32;
      WHEN COMP_LOOP_14_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110100");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_33;
      WHEN COMP_LOOP_14_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110101");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_34;
      WHEN COMP_LOOP_14_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110110");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_35;
      WHEN COMP_LOOP_14_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110111");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_36;
      WHEN COMP_LOOP_14_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111000");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_37;
      WHEN COMP_LOOP_14_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111001");
        state_var_NS <= COMP_LOOP_14_modExp_1_while_C_38;
      WHEN COMP_LOOP_14_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111010");
        IF ( COMP_LOOP_14_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_808;
        ELSE
          state_var_NS <= COMP_LOOP_14_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_808 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111011");
        state_var_NS <= COMP_LOOP_C_809;
      WHEN COMP_LOOP_C_809 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111100");
        state_var_NS <= COMP_LOOP_C_810;
      WHEN COMP_LOOP_C_810 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111101");
        state_var_NS <= COMP_LOOP_C_811;
      WHEN COMP_LOOP_C_811 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111110");
        state_var_NS <= COMP_LOOP_C_812;
      WHEN COMP_LOOP_C_812 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111111");
        state_var_NS <= COMP_LOOP_C_813;
      WHEN COMP_LOOP_C_813 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000000");
        state_var_NS <= COMP_LOOP_C_814;
      WHEN COMP_LOOP_C_814 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000001");
        state_var_NS <= COMP_LOOP_C_815;
      WHEN COMP_LOOP_C_815 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000010");
        state_var_NS <= COMP_LOOP_C_816;
      WHEN COMP_LOOP_C_816 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000011");
        state_var_NS <= COMP_LOOP_C_817;
      WHEN COMP_LOOP_C_817 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000100");
        state_var_NS <= COMP_LOOP_C_818;
      WHEN COMP_LOOP_C_818 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000101");
        state_var_NS <= COMP_LOOP_C_819;
      WHEN COMP_LOOP_C_819 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000110");
        state_var_NS <= COMP_LOOP_C_820;
      WHEN COMP_LOOP_C_820 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000111");
        state_var_NS <= COMP_LOOP_C_821;
      WHEN COMP_LOOP_C_821 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001000");
        state_var_NS <= COMP_LOOP_C_822;
      WHEN COMP_LOOP_C_822 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001001");
        state_var_NS <= COMP_LOOP_C_823;
      WHEN COMP_LOOP_C_823 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001010");
        state_var_NS <= COMP_LOOP_C_824;
      WHEN COMP_LOOP_C_824 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001011");
        state_var_NS <= COMP_LOOP_C_825;
      WHEN COMP_LOOP_C_825 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001100");
        state_var_NS <= COMP_LOOP_C_826;
      WHEN COMP_LOOP_C_826 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001101");
        state_var_NS <= COMP_LOOP_C_827;
      WHEN COMP_LOOP_C_827 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001110");
        state_var_NS <= COMP_LOOP_C_828;
      WHEN COMP_LOOP_C_828 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001111");
        state_var_NS <= COMP_LOOP_C_829;
      WHEN COMP_LOOP_C_829 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010000");
        state_var_NS <= COMP_LOOP_C_830;
      WHEN COMP_LOOP_C_830 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010001");
        state_var_NS <= COMP_LOOP_C_831;
      WHEN COMP_LOOP_C_831 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010010");
        state_var_NS <= COMP_LOOP_C_832;
      WHEN COMP_LOOP_C_832 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010011");
        state_var_NS <= COMP_LOOP_C_833;
      WHEN COMP_LOOP_C_833 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010100");
        state_var_NS <= COMP_LOOP_C_834;
      WHEN COMP_LOOP_C_834 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010101");
        state_var_NS <= COMP_LOOP_C_835;
      WHEN COMP_LOOP_C_835 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010110");
        state_var_NS <= COMP_LOOP_C_836;
      WHEN COMP_LOOP_C_836 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010111");
        state_var_NS <= COMP_LOOP_C_837;
      WHEN COMP_LOOP_C_837 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011000");
        state_var_NS <= COMP_LOOP_C_838;
      WHEN COMP_LOOP_C_838 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011001");
        state_var_NS <= COMP_LOOP_C_839;
      WHEN COMP_LOOP_C_839 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011010");
        state_var_NS <= COMP_LOOP_C_840;
      WHEN COMP_LOOP_C_840 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011011");
        state_var_NS <= COMP_LOOP_C_841;
      WHEN COMP_LOOP_C_841 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011100");
        state_var_NS <= COMP_LOOP_C_842;
      WHEN COMP_LOOP_C_842 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011101");
        state_var_NS <= COMP_LOOP_C_843;
      WHEN COMP_LOOP_C_843 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011110");
        state_var_NS <= COMP_LOOP_C_844;
      WHEN COMP_LOOP_C_844 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011111");
        state_var_NS <= COMP_LOOP_C_845;
      WHEN COMP_LOOP_C_845 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100000");
        state_var_NS <= COMP_LOOP_C_846;
      WHEN COMP_LOOP_C_846 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100001");
        state_var_NS <= COMP_LOOP_C_847;
      WHEN COMP_LOOP_C_847 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100010");
        state_var_NS <= COMP_LOOP_C_848;
      WHEN COMP_LOOP_C_848 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100011");
        state_var_NS <= COMP_LOOP_C_849;
      WHEN COMP_LOOP_C_849 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100100");
        state_var_NS <= COMP_LOOP_C_850;
      WHEN COMP_LOOP_C_850 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100101");
        state_var_NS <= COMP_LOOP_C_851;
      WHEN COMP_LOOP_C_851 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100110");
        state_var_NS <= COMP_LOOP_C_852;
      WHEN COMP_LOOP_C_852 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100111");
        state_var_NS <= COMP_LOOP_C_853;
      WHEN COMP_LOOP_C_853 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101000");
        state_var_NS <= COMP_LOOP_C_854;
      WHEN COMP_LOOP_C_854 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101001");
        state_var_NS <= COMP_LOOP_C_855;
      WHEN COMP_LOOP_C_855 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101010");
        state_var_NS <= COMP_LOOP_C_856;
      WHEN COMP_LOOP_C_856 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101011");
        state_var_NS <= COMP_LOOP_C_857;
      WHEN COMP_LOOP_C_857 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101100");
        state_var_NS <= COMP_LOOP_C_858;
      WHEN COMP_LOOP_C_858 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101101");
        state_var_NS <= COMP_LOOP_C_859;
      WHEN COMP_LOOP_C_859 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101110");
        state_var_NS <= COMP_LOOP_C_860;
      WHEN COMP_LOOP_C_860 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101111");
        state_var_NS <= COMP_LOOP_C_861;
      WHEN COMP_LOOP_C_861 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110000");
        state_var_NS <= COMP_LOOP_C_862;
      WHEN COMP_LOOP_C_862 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110001");
        state_var_NS <= COMP_LOOP_C_863;
      WHEN COMP_LOOP_C_863 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110010");
        state_var_NS <= COMP_LOOP_C_864;
      WHEN COMP_LOOP_C_864 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110011");
        state_var_NS <= COMP_LOOP_C_865;
      WHEN COMP_LOOP_C_865 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110100");
        state_var_NS <= COMP_LOOP_C_866;
      WHEN COMP_LOOP_C_866 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110101");
        state_var_NS <= COMP_LOOP_C_867;
      WHEN COMP_LOOP_C_867 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110110");
        state_var_NS <= COMP_LOOP_C_868;
      WHEN COMP_LOOP_C_868 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110111");
        IF ( COMP_LOOP_C_868_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_869;
        END IF;
      WHEN COMP_LOOP_C_869 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_0;
      WHEN COMP_LOOP_15_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_1;
      WHEN COMP_LOOP_15_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_2;
      WHEN COMP_LOOP_15_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_3;
      WHEN COMP_LOOP_15_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_4;
      WHEN COMP_LOOP_15_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_5;
      WHEN COMP_LOOP_15_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_6;
      WHEN COMP_LOOP_15_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_7;
      WHEN COMP_LOOP_15_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_8;
      WHEN COMP_LOOP_15_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_9;
      WHEN COMP_LOOP_15_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_10;
      WHEN COMP_LOOP_15_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_11;
      WHEN COMP_LOOP_15_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_12;
      WHEN COMP_LOOP_15_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_13;
      WHEN COMP_LOOP_15_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_14;
      WHEN COMP_LOOP_15_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_15;
      WHEN COMP_LOOP_15_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_16;
      WHEN COMP_LOOP_15_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_17;
      WHEN COMP_LOOP_15_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_18;
      WHEN COMP_LOOP_15_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_19;
      WHEN COMP_LOOP_15_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_20;
      WHEN COMP_LOOP_15_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_21;
      WHEN COMP_LOOP_15_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_22;
      WHEN COMP_LOOP_15_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_23;
      WHEN COMP_LOOP_15_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_24;
      WHEN COMP_LOOP_15_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_25;
      WHEN COMP_LOOP_15_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_26;
      WHEN COMP_LOOP_15_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_27;
      WHEN COMP_LOOP_15_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_28;
      WHEN COMP_LOOP_15_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_29;
      WHEN COMP_LOOP_15_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_30;
      WHEN COMP_LOOP_15_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010111");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_31;
      WHEN COMP_LOOP_15_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011000");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_32;
      WHEN COMP_LOOP_15_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011001");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_33;
      WHEN COMP_LOOP_15_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011010");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_34;
      WHEN COMP_LOOP_15_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011011");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_35;
      WHEN COMP_LOOP_15_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011100");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_36;
      WHEN COMP_LOOP_15_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011101");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_37;
      WHEN COMP_LOOP_15_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011110");
        state_var_NS <= COMP_LOOP_15_modExp_1_while_C_38;
      WHEN COMP_LOOP_15_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011111");
        IF ( COMP_LOOP_15_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_870;
        ELSE
          state_var_NS <= COMP_LOOP_15_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_870 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100000");
        state_var_NS <= COMP_LOOP_C_871;
      WHEN COMP_LOOP_C_871 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100001");
        state_var_NS <= COMP_LOOP_C_872;
      WHEN COMP_LOOP_C_872 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100010");
        state_var_NS <= COMP_LOOP_C_873;
      WHEN COMP_LOOP_C_873 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100011");
        state_var_NS <= COMP_LOOP_C_874;
      WHEN COMP_LOOP_C_874 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100100");
        state_var_NS <= COMP_LOOP_C_875;
      WHEN COMP_LOOP_C_875 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100101");
        state_var_NS <= COMP_LOOP_C_876;
      WHEN COMP_LOOP_C_876 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100110");
        state_var_NS <= COMP_LOOP_C_877;
      WHEN COMP_LOOP_C_877 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100111");
        state_var_NS <= COMP_LOOP_C_878;
      WHEN COMP_LOOP_C_878 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101000");
        state_var_NS <= COMP_LOOP_C_879;
      WHEN COMP_LOOP_C_879 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101001");
        state_var_NS <= COMP_LOOP_C_880;
      WHEN COMP_LOOP_C_880 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101010");
        state_var_NS <= COMP_LOOP_C_881;
      WHEN COMP_LOOP_C_881 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101011");
        state_var_NS <= COMP_LOOP_C_882;
      WHEN COMP_LOOP_C_882 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101100");
        state_var_NS <= COMP_LOOP_C_883;
      WHEN COMP_LOOP_C_883 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101101");
        state_var_NS <= COMP_LOOP_C_884;
      WHEN COMP_LOOP_C_884 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101110");
        state_var_NS <= COMP_LOOP_C_885;
      WHEN COMP_LOOP_C_885 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101111");
        state_var_NS <= COMP_LOOP_C_886;
      WHEN COMP_LOOP_C_886 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110000");
        state_var_NS <= COMP_LOOP_C_887;
      WHEN COMP_LOOP_C_887 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110001");
        state_var_NS <= COMP_LOOP_C_888;
      WHEN COMP_LOOP_C_888 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110010");
        state_var_NS <= COMP_LOOP_C_889;
      WHEN COMP_LOOP_C_889 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110011");
        state_var_NS <= COMP_LOOP_C_890;
      WHEN COMP_LOOP_C_890 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110100");
        state_var_NS <= COMP_LOOP_C_891;
      WHEN COMP_LOOP_C_891 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110101");
        state_var_NS <= COMP_LOOP_C_892;
      WHEN COMP_LOOP_C_892 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110110");
        state_var_NS <= COMP_LOOP_C_893;
      WHEN COMP_LOOP_C_893 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110111");
        state_var_NS <= COMP_LOOP_C_894;
      WHEN COMP_LOOP_C_894 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111000");
        state_var_NS <= COMP_LOOP_C_895;
      WHEN COMP_LOOP_C_895 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111001");
        state_var_NS <= COMP_LOOP_C_896;
      WHEN COMP_LOOP_C_896 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111010");
        state_var_NS <= COMP_LOOP_C_897;
      WHEN COMP_LOOP_C_897 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111011");
        state_var_NS <= COMP_LOOP_C_898;
      WHEN COMP_LOOP_C_898 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111100");
        state_var_NS <= COMP_LOOP_C_899;
      WHEN COMP_LOOP_C_899 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111101");
        state_var_NS <= COMP_LOOP_C_900;
      WHEN COMP_LOOP_C_900 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111110");
        state_var_NS <= COMP_LOOP_C_901;
      WHEN COMP_LOOP_C_901 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111111");
        state_var_NS <= COMP_LOOP_C_902;
      WHEN COMP_LOOP_C_902 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000000");
        state_var_NS <= COMP_LOOP_C_903;
      WHEN COMP_LOOP_C_903 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000001");
        state_var_NS <= COMP_LOOP_C_904;
      WHEN COMP_LOOP_C_904 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000010");
        state_var_NS <= COMP_LOOP_C_905;
      WHEN COMP_LOOP_C_905 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000011");
        state_var_NS <= COMP_LOOP_C_906;
      WHEN COMP_LOOP_C_906 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000100");
        state_var_NS <= COMP_LOOP_C_907;
      WHEN COMP_LOOP_C_907 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000101");
        state_var_NS <= COMP_LOOP_C_908;
      WHEN COMP_LOOP_C_908 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000110");
        state_var_NS <= COMP_LOOP_C_909;
      WHEN COMP_LOOP_C_909 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000111");
        state_var_NS <= COMP_LOOP_C_910;
      WHEN COMP_LOOP_C_910 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001000");
        state_var_NS <= COMP_LOOP_C_911;
      WHEN COMP_LOOP_C_911 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001001");
        state_var_NS <= COMP_LOOP_C_912;
      WHEN COMP_LOOP_C_912 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001010");
        state_var_NS <= COMP_LOOP_C_913;
      WHEN COMP_LOOP_C_913 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001011");
        state_var_NS <= COMP_LOOP_C_914;
      WHEN COMP_LOOP_C_914 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001100");
        state_var_NS <= COMP_LOOP_C_915;
      WHEN COMP_LOOP_C_915 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001101");
        state_var_NS <= COMP_LOOP_C_916;
      WHEN COMP_LOOP_C_916 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001110");
        state_var_NS <= COMP_LOOP_C_917;
      WHEN COMP_LOOP_C_917 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001111");
        state_var_NS <= COMP_LOOP_C_918;
      WHEN COMP_LOOP_C_918 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010000");
        state_var_NS <= COMP_LOOP_C_919;
      WHEN COMP_LOOP_C_919 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010001");
        state_var_NS <= COMP_LOOP_C_920;
      WHEN COMP_LOOP_C_920 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010010");
        state_var_NS <= COMP_LOOP_C_921;
      WHEN COMP_LOOP_C_921 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010011");
        state_var_NS <= COMP_LOOP_C_922;
      WHEN COMP_LOOP_C_922 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010100");
        state_var_NS <= COMP_LOOP_C_923;
      WHEN COMP_LOOP_C_923 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010101");
        state_var_NS <= COMP_LOOP_C_924;
      WHEN COMP_LOOP_C_924 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010110");
        state_var_NS <= COMP_LOOP_C_925;
      WHEN COMP_LOOP_C_925 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010111");
        state_var_NS <= COMP_LOOP_C_926;
      WHEN COMP_LOOP_C_926 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011000");
        state_var_NS <= COMP_LOOP_C_927;
      WHEN COMP_LOOP_C_927 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011001");
        state_var_NS <= COMP_LOOP_C_928;
      WHEN COMP_LOOP_C_928 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011010");
        state_var_NS <= COMP_LOOP_C_929;
      WHEN COMP_LOOP_C_929 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011011");
        state_var_NS <= COMP_LOOP_C_930;
      WHEN COMP_LOOP_C_930 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011100");
        IF ( COMP_LOOP_C_930_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_931;
        END IF;
      WHEN COMP_LOOP_C_931 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_0;
      WHEN COMP_LOOP_16_modExp_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_1;
      WHEN COMP_LOOP_16_modExp_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_2;
      WHEN COMP_LOOP_16_modExp_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_3;
      WHEN COMP_LOOP_16_modExp_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_4;
      WHEN COMP_LOOP_16_modExp_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_5;
      WHEN COMP_LOOP_16_modExp_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_6;
      WHEN COMP_LOOP_16_modExp_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_7;
      WHEN COMP_LOOP_16_modExp_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_8;
      WHEN COMP_LOOP_16_modExp_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_9;
      WHEN COMP_LOOP_16_modExp_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_10;
      WHEN COMP_LOOP_16_modExp_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_11;
      WHEN COMP_LOOP_16_modExp_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_12;
      WHEN COMP_LOOP_16_modExp_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_13;
      WHEN COMP_LOOP_16_modExp_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_14;
      WHEN COMP_LOOP_16_modExp_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_15;
      WHEN COMP_LOOP_16_modExp_1_while_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_16;
      WHEN COMP_LOOP_16_modExp_1_while_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_17;
      WHEN COMP_LOOP_16_modExp_1_while_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_18;
      WHEN COMP_LOOP_16_modExp_1_while_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_19;
      WHEN COMP_LOOP_16_modExp_1_while_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_20;
      WHEN COMP_LOOP_16_modExp_1_while_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_21;
      WHEN COMP_LOOP_16_modExp_1_while_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_22;
      WHEN COMP_LOOP_16_modExp_1_while_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_23;
      WHEN COMP_LOOP_16_modExp_1_while_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_24;
      WHEN COMP_LOOP_16_modExp_1_while_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_25;
      WHEN COMP_LOOP_16_modExp_1_while_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_26;
      WHEN COMP_LOOP_16_modExp_1_while_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_27;
      WHEN COMP_LOOP_16_modExp_1_while_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_28;
      WHEN COMP_LOOP_16_modExp_1_while_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_29;
      WHEN COMP_LOOP_16_modExp_1_while_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_30;
      WHEN COMP_LOOP_16_modExp_1_while_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111100");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_31;
      WHEN COMP_LOOP_16_modExp_1_while_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111101");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_32;
      WHEN COMP_LOOP_16_modExp_1_while_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111110");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_33;
      WHEN COMP_LOOP_16_modExp_1_while_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111111");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_34;
      WHEN COMP_LOOP_16_modExp_1_while_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000000");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_35;
      WHEN COMP_LOOP_16_modExp_1_while_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000001");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_36;
      WHEN COMP_LOOP_16_modExp_1_while_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000010");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_37;
      WHEN COMP_LOOP_16_modExp_1_while_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000011");
        state_var_NS <= COMP_LOOP_16_modExp_1_while_C_38;
      WHEN COMP_LOOP_16_modExp_1_while_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000100");
        IF ( COMP_LOOP_16_modExp_1_while_C_38_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_932;
        ELSE
          state_var_NS <= COMP_LOOP_16_modExp_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_932 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000101");
        state_var_NS <= COMP_LOOP_C_933;
      WHEN COMP_LOOP_C_933 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000110");
        state_var_NS <= COMP_LOOP_C_934;
      WHEN COMP_LOOP_C_934 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000111");
        state_var_NS <= COMP_LOOP_C_935;
      WHEN COMP_LOOP_C_935 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001000");
        state_var_NS <= COMP_LOOP_C_936;
      WHEN COMP_LOOP_C_936 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001001");
        state_var_NS <= COMP_LOOP_C_937;
      WHEN COMP_LOOP_C_937 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001010");
        state_var_NS <= COMP_LOOP_C_938;
      WHEN COMP_LOOP_C_938 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001011");
        state_var_NS <= COMP_LOOP_C_939;
      WHEN COMP_LOOP_C_939 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001100");
        state_var_NS <= COMP_LOOP_C_940;
      WHEN COMP_LOOP_C_940 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001101");
        state_var_NS <= COMP_LOOP_C_941;
      WHEN COMP_LOOP_C_941 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001110");
        state_var_NS <= COMP_LOOP_C_942;
      WHEN COMP_LOOP_C_942 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001111");
        state_var_NS <= COMP_LOOP_C_943;
      WHEN COMP_LOOP_C_943 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010000");
        state_var_NS <= COMP_LOOP_C_944;
      WHEN COMP_LOOP_C_944 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010001");
        state_var_NS <= COMP_LOOP_C_945;
      WHEN COMP_LOOP_C_945 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010010");
        state_var_NS <= COMP_LOOP_C_946;
      WHEN COMP_LOOP_C_946 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010011");
        state_var_NS <= COMP_LOOP_C_947;
      WHEN COMP_LOOP_C_947 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010100");
        state_var_NS <= COMP_LOOP_C_948;
      WHEN COMP_LOOP_C_948 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010101");
        state_var_NS <= COMP_LOOP_C_949;
      WHEN COMP_LOOP_C_949 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010110");
        state_var_NS <= COMP_LOOP_C_950;
      WHEN COMP_LOOP_C_950 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010111");
        state_var_NS <= COMP_LOOP_C_951;
      WHEN COMP_LOOP_C_951 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011000");
        state_var_NS <= COMP_LOOP_C_952;
      WHEN COMP_LOOP_C_952 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011001");
        state_var_NS <= COMP_LOOP_C_953;
      WHEN COMP_LOOP_C_953 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011010");
        state_var_NS <= COMP_LOOP_C_954;
      WHEN COMP_LOOP_C_954 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011011");
        state_var_NS <= COMP_LOOP_C_955;
      WHEN COMP_LOOP_C_955 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011100");
        state_var_NS <= COMP_LOOP_C_956;
      WHEN COMP_LOOP_C_956 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011101");
        state_var_NS <= COMP_LOOP_C_957;
      WHEN COMP_LOOP_C_957 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011110");
        state_var_NS <= COMP_LOOP_C_958;
      WHEN COMP_LOOP_C_958 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011111");
        state_var_NS <= COMP_LOOP_C_959;
      WHEN COMP_LOOP_C_959 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100000");
        state_var_NS <= COMP_LOOP_C_960;
      WHEN COMP_LOOP_C_960 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100001");
        state_var_NS <= COMP_LOOP_C_961;
      WHEN COMP_LOOP_C_961 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100010");
        state_var_NS <= COMP_LOOP_C_962;
      WHEN COMP_LOOP_C_962 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100011");
        state_var_NS <= COMP_LOOP_C_963;
      WHEN COMP_LOOP_C_963 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100100");
        state_var_NS <= COMP_LOOP_C_964;
      WHEN COMP_LOOP_C_964 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100101");
        state_var_NS <= COMP_LOOP_C_965;
      WHEN COMP_LOOP_C_965 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100110");
        state_var_NS <= COMP_LOOP_C_966;
      WHEN COMP_LOOP_C_966 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100111");
        state_var_NS <= COMP_LOOP_C_967;
      WHEN COMP_LOOP_C_967 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101000");
        state_var_NS <= COMP_LOOP_C_968;
      WHEN COMP_LOOP_C_968 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101001");
        state_var_NS <= COMP_LOOP_C_969;
      WHEN COMP_LOOP_C_969 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101010");
        state_var_NS <= COMP_LOOP_C_970;
      WHEN COMP_LOOP_C_970 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101011");
        state_var_NS <= COMP_LOOP_C_971;
      WHEN COMP_LOOP_C_971 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101100");
        state_var_NS <= COMP_LOOP_C_972;
      WHEN COMP_LOOP_C_972 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101101");
        state_var_NS <= COMP_LOOP_C_973;
      WHEN COMP_LOOP_C_973 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101110");
        state_var_NS <= COMP_LOOP_C_974;
      WHEN COMP_LOOP_C_974 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101111");
        state_var_NS <= COMP_LOOP_C_975;
      WHEN COMP_LOOP_C_975 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110000");
        state_var_NS <= COMP_LOOP_C_976;
      WHEN COMP_LOOP_C_976 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110001");
        state_var_NS <= COMP_LOOP_C_977;
      WHEN COMP_LOOP_C_977 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110010");
        state_var_NS <= COMP_LOOP_C_978;
      WHEN COMP_LOOP_C_978 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110011");
        state_var_NS <= COMP_LOOP_C_979;
      WHEN COMP_LOOP_C_979 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110100");
        state_var_NS <= COMP_LOOP_C_980;
      WHEN COMP_LOOP_C_980 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110101");
        state_var_NS <= COMP_LOOP_C_981;
      WHEN COMP_LOOP_C_981 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110110");
        state_var_NS <= COMP_LOOP_C_982;
      WHEN COMP_LOOP_C_982 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110111");
        state_var_NS <= COMP_LOOP_C_983;
      WHEN COMP_LOOP_C_983 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111000");
        state_var_NS <= COMP_LOOP_C_984;
      WHEN COMP_LOOP_C_984 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111001");
        state_var_NS <= COMP_LOOP_C_985;
      WHEN COMP_LOOP_C_985 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111010");
        state_var_NS <= COMP_LOOP_C_986;
      WHEN COMP_LOOP_C_986 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111011");
        state_var_NS <= COMP_LOOP_C_987;
      WHEN COMP_LOOP_C_987 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111100");
        state_var_NS <= COMP_LOOP_C_988;
      WHEN COMP_LOOP_C_988 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111101");
        state_var_NS <= COMP_LOOP_C_989;
      WHEN COMP_LOOP_C_989 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111110");
        state_var_NS <= COMP_LOOP_C_990;
      WHEN COMP_LOOP_C_990 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111111");
        state_var_NS <= COMP_LOOP_C_991;
      WHEN COMP_LOOP_C_991 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000000");
        state_var_NS <= COMP_LOOP_C_992;
      WHEN COMP_LOOP_C_992 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000001");
        IF ( COMP_LOOP_C_992_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000010");
        IF ( VEC_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_9;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000011");
        IF ( STAGE_LOOP_C_9_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000100");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS inPlaceNTT_DIT_core_core_fsm_1;

  inPlaceNTT_DIT_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIT_core_core_fsm_1_REG;

END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
    vec_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC
  );
END inPlaceNTT_DIT_core;

ARCHITECTURE v43 OF inPlaceNTT_DIT_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_b_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL or_tmp_3 : STD_LOGIC;
  SIGNAL or_tmp_4 : STD_LOGIC;
  SIGNAL or_tmp_8 : STD_LOGIC;
  SIGNAL or_tmp_9 : STD_LOGIC;
  SIGNAL or_tmp_14 : STD_LOGIC;
  SIGNAL nor_tmp_6 : STD_LOGIC;
  SIGNAL or_tmp_21 : STD_LOGIC;
  SIGNAL nor_tmp_9 : STD_LOGIC;
  SIGNAL not_tmp_34 : STD_LOGIC;
  SIGNAL not_tmp_45 : STD_LOGIC;
  SIGNAL or_tmp_110 : STD_LOGIC;
  SIGNAL not_tmp_51 : STD_LOGIC;
  SIGNAL or_tmp_118 : STD_LOGIC;
  SIGNAL or_tmp_141 : STD_LOGIC;
  SIGNAL mux_tmp_207 : STD_LOGIC;
  SIGNAL mux_tmp_226 : STD_LOGIC;
  SIGNAL or_tmp_150 : STD_LOGIC;
  SIGNAL or_tmp_178 : STD_LOGIC;
  SIGNAL or_tmp_179 : STD_LOGIC;
  SIGNAL or_tmp_180 : STD_LOGIC;
  SIGNAL or_tmp_181 : STD_LOGIC;
  SIGNAL mux_tmp_373 : STD_LOGIC;
  SIGNAL or_tmp_182 : STD_LOGIC;
  SIGNAL mux_tmp_374 : STD_LOGIC;
  SIGNAL mux_tmp_375 : STD_LOGIC;
  SIGNAL or_tmp_183 : STD_LOGIC;
  SIGNAL mux_tmp_378 : STD_LOGIC;
  SIGNAL mux_tmp_379 : STD_LOGIC;
  SIGNAL mux_tmp_380 : STD_LOGIC;
  SIGNAL mux_tmp_381 : STD_LOGIC;
  SIGNAL nor_tmp_46 : STD_LOGIC;
  SIGNAL nand_tmp_12 : STD_LOGIC;
  SIGNAL nand_tmp_13 : STD_LOGIC;
  SIGNAL or_tmp_187 : STD_LOGIC;
  SIGNAL mux_tmp_399 : STD_LOGIC;
  SIGNAL or_tmp_188 : STD_LOGIC;
  SIGNAL or_tmp_189 : STD_LOGIC;
  SIGNAL or_tmp_191 : STD_LOGIC;
  SIGNAL nand_tmp_14 : STD_LOGIC;
  SIGNAL or_tmp_195 : STD_LOGIC;
  SIGNAL mux_tmp_412 : STD_LOGIC;
  SIGNAL mux_tmp_413 : STD_LOGIC;
  SIGNAL and_dcpl : STD_LOGIC;
  SIGNAL and_dcpl_1 : STD_LOGIC;
  SIGNAL and_dcpl_2 : STD_LOGIC;
  SIGNAL or_tmp_237 : STD_LOGIC;
  SIGNAL nor_tmp_116 : STD_LOGIC;
  SIGNAL mux_tmp_741 : STD_LOGIC;
  SIGNAL or_tmp_434 : STD_LOGIC;
  SIGNAL mux_tmp_893 : STD_LOGIC;
  SIGNAL mux_tmp_917 : STD_LOGIC;
  SIGNAL and_dcpl_21 : STD_LOGIC;
  SIGNAL and_dcpl_22 : STD_LOGIC;
  SIGNAL and_dcpl_26 : STD_LOGIC;
  SIGNAL and_dcpl_30 : STD_LOGIC;
  SIGNAL and_dcpl_31 : STD_LOGIC;
  SIGNAL and_dcpl_32 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_46 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL not_tmp_219 : STD_LOGIC;
  SIGNAL and_dcpl_96 : STD_LOGIC;
  SIGNAL and_dcpl_97 : STD_LOGIC;
  SIGNAL and_dcpl_98 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_100 : STD_LOGIC;
  SIGNAL and_dcpl_101 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_106 : STD_LOGIC;
  SIGNAL and_dcpl_107 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_116 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_118 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL and_dcpl_121 : STD_LOGIC;
  SIGNAL and_dcpl_122 : STD_LOGIC;
  SIGNAL and_dcpl_123 : STD_LOGIC;
  SIGNAL and_dcpl_124 : STD_LOGIC;
  SIGNAL and_dcpl_125 : STD_LOGIC;
  SIGNAL and_dcpl_126 : STD_LOGIC;
  SIGNAL and_dcpl_127 : STD_LOGIC;
  SIGNAL and_dcpl_128 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL or_tmp_453 : STD_LOGIC;
  SIGNAL not_tmp_240 : STD_LOGIC;
  SIGNAL and_dcpl_139 : STD_LOGIC;
  SIGNAL and_dcpl_140 : STD_LOGIC;
  SIGNAL and_dcpl_141 : STD_LOGIC;
  SIGNAL and_dcpl_145 : STD_LOGIC;
  SIGNAL and_dcpl_146 : STD_LOGIC;
  SIGNAL and_dcpl_147 : STD_LOGIC;
  SIGNAL and_dcpl_148 : STD_LOGIC;
  SIGNAL and_dcpl_154 : STD_LOGIC;
  SIGNAL and_dcpl_156 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_162 : STD_LOGIC;
  SIGNAL and_dcpl_164 : STD_LOGIC;
  SIGNAL and_dcpl_165 : STD_LOGIC;
  SIGNAL nor_tmp_217 : STD_LOGIC;
  SIGNAL mux_tmp_1049 : STD_LOGIC;
  SIGNAL and_dcpl_172 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_182 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_198 : STD_LOGIC;
  SIGNAL and_dcpl_204 : STD_LOGIC;
  SIGNAL and_dcpl_206 : STD_LOGIC;
  SIGNAL and_dcpl_215 : STD_LOGIC;
  SIGNAL and_dcpl_217 : STD_LOGIC;
  SIGNAL and_dcpl_223 : STD_LOGIC;
  SIGNAL and_dcpl_225 : STD_LOGIC;
  SIGNAL and_dcpl_232 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_240 : STD_LOGIC;
  SIGNAL and_dcpl_242 : STD_LOGIC;
  SIGNAL and_dcpl_243 : STD_LOGIC;
  SIGNAL and_dcpl_245 : STD_LOGIC;
  SIGNAL and_dcpl_247 : STD_LOGIC;
  SIGNAL and_dcpl_255 : STD_LOGIC;
  SIGNAL or_tmp_515 : STD_LOGIC;
  SIGNAL or_tmp_518 : STD_LOGIC;
  SIGNAL mux_tmp_1062 : STD_LOGIC;
  SIGNAL mux_tmp_1067 : STD_LOGIC;
  SIGNAL mux_tmp_1068 : STD_LOGIC;
  SIGNAL not_tmp_260 : STD_LOGIC;
  SIGNAL or_tmp_626 : STD_LOGIC;
  SIGNAL or_tmp_630 : STD_LOGIC;
  SIGNAL mux_tmp_1139 : STD_LOGIC;
  SIGNAL mux_tmp_1150 : STD_LOGIC;
  SIGNAL mux_tmp_1152 : STD_LOGIC;
  SIGNAL or_tmp_728 : STD_LOGIC;
  SIGNAL or_tmp_731 : STD_LOGIC;
  SIGNAL mux_tmp_1206 : STD_LOGIC;
  SIGNAL mux_tmp_1211 : STD_LOGIC;
  SIGNAL mux_tmp_1212 : STD_LOGIC;
  SIGNAL or_tmp_839 : STD_LOGIC;
  SIGNAL or_tmp_843 : STD_LOGIC;
  SIGNAL mux_tmp_1283 : STD_LOGIC;
  SIGNAL mux_tmp_1294 : STD_LOGIC;
  SIGNAL mux_tmp_1296 : STD_LOGIC;
  SIGNAL or_tmp_941 : STD_LOGIC;
  SIGNAL or_tmp_944 : STD_LOGIC;
  SIGNAL mux_tmp_1350 : STD_LOGIC;
  SIGNAL mux_tmp_1355 : STD_LOGIC;
  SIGNAL mux_tmp_1356 : STD_LOGIC;
  SIGNAL or_tmp_1052 : STD_LOGIC;
  SIGNAL or_tmp_1056 : STD_LOGIC;
  SIGNAL mux_tmp_1427 : STD_LOGIC;
  SIGNAL mux_tmp_1438 : STD_LOGIC;
  SIGNAL mux_tmp_1440 : STD_LOGIC;
  SIGNAL or_tmp_1154 : STD_LOGIC;
  SIGNAL or_tmp_1157 : STD_LOGIC;
  SIGNAL mux_tmp_1494 : STD_LOGIC;
  SIGNAL mux_tmp_1499 : STD_LOGIC;
  SIGNAL mux_tmp_1500 : STD_LOGIC;
  SIGNAL or_tmp_1265 : STD_LOGIC;
  SIGNAL or_tmp_1269 : STD_LOGIC;
  SIGNAL mux_tmp_1571 : STD_LOGIC;
  SIGNAL mux_tmp_1582 : STD_LOGIC;
  SIGNAL mux_tmp_1584 : STD_LOGIC;
  SIGNAL or_tmp_1367 : STD_LOGIC;
  SIGNAL or_tmp_1370 : STD_LOGIC;
  SIGNAL mux_tmp_1638 : STD_LOGIC;
  SIGNAL mux_tmp_1643 : STD_LOGIC;
  SIGNAL mux_tmp_1644 : STD_LOGIC;
  SIGNAL or_tmp_1478 : STD_LOGIC;
  SIGNAL or_tmp_1482 : STD_LOGIC;
  SIGNAL mux_tmp_1715 : STD_LOGIC;
  SIGNAL mux_tmp_1726 : STD_LOGIC;
  SIGNAL mux_tmp_1728 : STD_LOGIC;
  SIGNAL or_tmp_1580 : STD_LOGIC;
  SIGNAL or_tmp_1583 : STD_LOGIC;
  SIGNAL mux_tmp_1782 : STD_LOGIC;
  SIGNAL mux_tmp_1787 : STD_LOGIC;
  SIGNAL mux_tmp_1788 : STD_LOGIC;
  SIGNAL or_tmp_1691 : STD_LOGIC;
  SIGNAL or_tmp_1695 : STD_LOGIC;
  SIGNAL mux_tmp_1859 : STD_LOGIC;
  SIGNAL mux_tmp_1870 : STD_LOGIC;
  SIGNAL mux_tmp_1872 : STD_LOGIC;
  SIGNAL or_tmp_1797 : STD_LOGIC;
  SIGNAL not_tmp_378 : STD_LOGIC;
  SIGNAL mux_tmp_1927 : STD_LOGIC;
  SIGNAL nand_tmp_74 : STD_LOGIC;
  SIGNAL or_tmp_1811 : STD_LOGIC;
  SIGNAL or_tmp_1812 : STD_LOGIC;
  SIGNAL not_tmp_381 : STD_LOGIC;
  SIGNAL or_tmp_1821 : STD_LOGIC;
  SIGNAL or_tmp_1907 : STD_LOGIC;
  SIGNAL or_tmp_1911 : STD_LOGIC;
  SIGNAL mux_tmp_2004 : STD_LOGIC;
  SIGNAL mux_tmp_2015 : STD_LOGIC;
  SIGNAL mux_tmp_2017 : STD_LOGIC;
  SIGNAL or_tmp_2009 : STD_LOGIC;
  SIGNAL or_tmp_2012 : STD_LOGIC;
  SIGNAL mux_tmp_2071 : STD_LOGIC;
  SIGNAL mux_tmp_2076 : STD_LOGIC;
  SIGNAL mux_tmp_2077 : STD_LOGIC;
  SIGNAL or_tmp_2120 : STD_LOGIC;
  SIGNAL or_tmp_2124 : STD_LOGIC;
  SIGNAL mux_tmp_2148 : STD_LOGIC;
  SIGNAL mux_tmp_2159 : STD_LOGIC;
  SIGNAL mux_tmp_2161 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL or_tmp_2220 : STD_LOGIC;
  SIGNAL or_tmp_2223 : STD_LOGIC;
  SIGNAL or_tmp_2225 : STD_LOGIC;
  SIGNAL or_tmp_2230 : STD_LOGIC;
  SIGNAL or_tmp_2233 : STD_LOGIC;
  SIGNAL mux_tmp_2218 : STD_LOGIC;
  SIGNAL mux_tmp_2220 : STD_LOGIC;
  SIGNAL mux_tmp_2223 : STD_LOGIC;
  SIGNAL or_tmp_2237 : STD_LOGIC;
  SIGNAL or_tmp_2238 : STD_LOGIC;
  SIGNAL mux_tmp_2239 : STD_LOGIC;
  SIGNAL nand_tmp_92 : STD_LOGIC;
  SIGNAL nor_tmp_286 : STD_LOGIC;
  SIGNAL or_tmp_2246 : STD_LOGIC;
  SIGNAL or_tmp_2248 : STD_LOGIC;
  SIGNAL not_tmp_426 : STD_LOGIC;
  SIGNAL nor_tmp_288 : STD_LOGIC;
  SIGNAL and_tmp_10 : STD_LOGIC;
  SIGNAL mux_tmp_2250 : STD_LOGIC;
  SIGNAL mux_tmp_2251 : STD_LOGIC;
  SIGNAL mux_tmp_2254 : STD_LOGIC;
  SIGNAL or_tmp_2253 : STD_LOGIC;
  SIGNAL or_tmp_2255 : STD_LOGIC;
  SIGNAL mux_tmp_2265 : STD_LOGIC;
  SIGNAL nor_tmp_291 : STD_LOGIC;
  SIGNAL or_tmp_2257 : STD_LOGIC;
  SIGNAL nor_tmp_295 : STD_LOGIC;
  SIGNAL mux_tmp_2285 : STD_LOGIC;
  SIGNAL mux_tmp_2290 : STD_LOGIC;
  SIGNAL or_tmp_2260 : STD_LOGIC;
  SIGNAL or_tmp_2263 : STD_LOGIC;
  SIGNAL nand_tmp_93 : STD_LOGIC;
  SIGNAL or_tmp_2266 : STD_LOGIC;
  SIGNAL mux_tmp_2309 : STD_LOGIC;
  SIGNAL or_tmp_2267 : STD_LOGIC;
  SIGNAL or_tmp_2269 : STD_LOGIC;
  SIGNAL nand_tmp_95 : STD_LOGIC;
  SIGNAL or_tmp_2271 : STD_LOGIC;
  SIGNAL nand_tmp_96 : STD_LOGIC;
  SIGNAL or_tmp_2275 : STD_LOGIC;
  SIGNAL or_tmp_2276 : STD_LOGIC;
  SIGNAL or_tmp_2277 : STD_LOGIC;
  SIGNAL mux_tmp_2327 : STD_LOGIC;
  SIGNAL or_tmp_2280 : STD_LOGIC;
  SIGNAL or_tmp_2281 : STD_LOGIC;
  SIGNAL or_tmp_2282 : STD_LOGIC;
  SIGNAL or_tmp_2289 : STD_LOGIC;
  SIGNAL not_tmp_463 : STD_LOGIC;
  SIGNAL mux_tmp_2349 : STD_LOGIC;
  SIGNAL and_tmp_16 : STD_LOGIC;
  SIGNAL or_tmp_2293 : STD_LOGIC;
  SIGNAL mux_tmp_2362 : STD_LOGIC;
  SIGNAL nor_tmp_300 : STD_LOGIC;
  SIGNAL or_tmp_2327 : STD_LOGIC;
  SIGNAL or_tmp_2329 : STD_LOGIC;
  SIGNAL or_tmp_2331 : STD_LOGIC;
  SIGNAL or_tmp_2333 : STD_LOGIC;
  SIGNAL or_tmp_2334 : STD_LOGIC;
  SIGNAL mux_tmp_2400 : STD_LOGIC;
  SIGNAL mux_tmp_2401 : STD_LOGIC;
  SIGNAL mux_tmp_2402 : STD_LOGIC;
  SIGNAL or_tmp_2335 : STD_LOGIC;
  SIGNAL mux_tmp_2406 : STD_LOGIC;
  SIGNAL or_tmp_2338 : STD_LOGIC;
  SIGNAL nand_tmp_105 : STD_LOGIC;
  SIGNAL mux_tmp_2423 : STD_LOGIC;
  SIGNAL nor_tmp_307 : STD_LOGIC;
  SIGNAL mux_tmp_2425 : STD_LOGIC;
  SIGNAL mux_tmp_2426 : STD_LOGIC;
  SIGNAL or_tmp_2342 : STD_LOGIC;
  SIGNAL or_tmp_2343 : STD_LOGIC;
  SIGNAL mux_tmp_2436 : STD_LOGIC;
  SIGNAL nand_tmp_107 : STD_LOGIC;
  SIGNAL nand_tmp_108 : STD_LOGIC;
  SIGNAL mux_tmp_2466 : STD_LOGIC;
  SIGNAL not_tmp_519 : STD_LOGIC;
  SIGNAL and_dcpl_264 : STD_LOGIC;
  SIGNAL and_dcpl_266 : STD_LOGIC;
  SIGNAL and_dcpl_268 : STD_LOGIC;
  SIGNAL and_dcpl_273 : STD_LOGIC;
  SIGNAL mux_tmp_2502 : STD_LOGIC;
  SIGNAL not_tmp_529 : STD_LOGIC;
  SIGNAL nor_tmp_330 : STD_LOGIC;
  SIGNAL mux_tmp_2508 : STD_LOGIC;
  SIGNAL or_tmp_2416 : STD_LOGIC;
  SIGNAL or_tmp_2419 : STD_LOGIC;
  SIGNAL mux_tmp_2519 : STD_LOGIC;
  SIGNAL mux_tmp_2523 : STD_LOGIC;
  SIGNAL mux_tmp_2525 : STD_LOGIC;
  SIGNAL nor_tmp_338 : STD_LOGIC;
  SIGNAL or_tmp_2429 : STD_LOGIC;
  SIGNAL nor_tmp_342 : STD_LOGIC;
  SIGNAL mux_tmp_2549 : STD_LOGIC;
  SIGNAL mux_tmp_2650 : STD_LOGIC;
  SIGNAL and_dcpl_279 : STD_LOGIC;
  SIGNAL and_dcpl_281 : STD_LOGIC;
  SIGNAL mux_tmp_2687 : STD_LOGIC;
  SIGNAL or_tmp_2474 : STD_LOGIC;
  SIGNAL mux_tmp_2696 : STD_LOGIC;
  SIGNAL mux_tmp_2698 : STD_LOGIC;
  SIGNAL mux_tmp_2701 : STD_LOGIC;
  SIGNAL or_tmp_2479 : STD_LOGIC;
  SIGNAL nand_tmp_119 : STD_LOGIC;
  SIGNAL or_tmp_2483 : STD_LOGIC;
  SIGNAL and_dcpl_283 : STD_LOGIC;
  SIGNAL and_dcpl_305 : STD_LOGIC;
  SIGNAL not_tmp_596 : STD_LOGIC;
  SIGNAL or_tmp_2516 : STD_LOGIC;
  SIGNAL mux_tmp_2758 : STD_LOGIC;
  SIGNAL mux_tmp_2788 : STD_LOGIC;
  SIGNAL mux_tmp_2790 : STD_LOGIC;
  SIGNAL mux_tmp_2796 : STD_LOGIC;
  SIGNAL mux_tmp_2800 : STD_LOGIC;
  SIGNAL mux_tmp_2813 : STD_LOGIC;
  SIGNAL or_tmp_2594 : STD_LOGIC;
  SIGNAL not_tmp_634 : STD_LOGIC;
  SIGNAL or_tmp_2631 : STD_LOGIC;
  SIGNAL not_tmp_646 : STD_LOGIC;
  SIGNAL or_tmp_2649 : STD_LOGIC;
  SIGNAL nand_tmp_136 : STD_LOGIC;
  SIGNAL mux_tmp_2905 : STD_LOGIC;
  SIGNAL nand_tmp_137 : STD_LOGIC;
  SIGNAL mux_tmp_2907 : STD_LOGIC;
  SIGNAL or_tmp_2652 : STD_LOGIC;
  SIGNAL or_tmp_2653 : STD_LOGIC;
  SIGNAL mux_tmp_2911 : STD_LOGIC;
  SIGNAL mux_tmp_2912 : STD_LOGIC;
  SIGNAL mux_tmp_2913 : STD_LOGIC;
  SIGNAL mux_tmp_2919 : STD_LOGIC;
  SIGNAL mux_tmp_2921 : STD_LOGIC;
  SIGNAL mux_tmp_2930 : STD_LOGIC;
  SIGNAL or_tmp_2659 : STD_LOGIC;
  SIGNAL or_tmp_2663 : STD_LOGIC;
  SIGNAL nand_tmp_140 : STD_LOGIC;
  SIGNAL or_tmp_2707 : STD_LOGIC;
  SIGNAL and_dcpl_332 : STD_LOGIC;
  SIGNAL nand_tmp_148 : STD_LOGIC;
  SIGNAL not_tmp_708 : STD_LOGIC;
  SIGNAL nor_tmp_445 : STD_LOGIC;
  SIGNAL mux_tmp_3219 : STD_LOGIC;
  SIGNAL mux_tmp_3236 : STD_LOGIC;
  SIGNAL or_tmp_2849 : STD_LOGIC;
  SIGNAL mux_tmp_3244 : STD_LOGIC;
  SIGNAL nor_tmp_456 : STD_LOGIC;
  SIGNAL mux_tmp_3256 : STD_LOGIC;
  SIGNAL not_tmp_728 : STD_LOGIC;
  SIGNAL or_tmp_2864 : STD_LOGIC;
  SIGNAL mux_tmp_3269 : STD_LOGIC;
  SIGNAL nor_tmp_461 : STD_LOGIC;
  SIGNAL mux_tmp_3280 : STD_LOGIC;
  SIGNAL mux_tmp_3281 : STD_LOGIC;
  SIGNAL nand_tmp_157 : STD_LOGIC;
  SIGNAL mux_tmp_3323 : STD_LOGIC;
  SIGNAL not_tmp_762 : STD_LOGIC;
  SIGNAL mux_tmp_3386 : STD_LOGIC;
  SIGNAL not_tmp_776 : STD_LOGIC;
  SIGNAL mux_tmp_3418 : STD_LOGIC;
  SIGNAL mux_tmp_3422 : STD_LOGIC;
  SIGNAL mux_tmp_3426 : STD_LOGIC;
  SIGNAL mux_tmp_3430 : STD_LOGIC;
  SIGNAL mux_tmp_3436 : STD_LOGIC;
  SIGNAL nand_tmp_167 : STD_LOGIC;
  SIGNAL mux_tmp_3449 : STD_LOGIC;
  SIGNAL mux_tmp_3450 : STD_LOGIC;
  SIGNAL mux_tmp_3452 : STD_LOGIC;
  SIGNAL mux_tmp_3456 : STD_LOGIC;
  SIGNAL mux_tmp_3458 : STD_LOGIC;
  SIGNAL mux_tmp_3459 : STD_LOGIC;
  SIGNAL mux_tmp_3467 : STD_LOGIC;
  SIGNAL mux_tmp_3468 : STD_LOGIC;
  SIGNAL mux_tmp_3471 : STD_LOGIC;
  SIGNAL and_tmp_36 : STD_LOGIC;
  SIGNAL or_tmp_3025 : STD_LOGIC;
  SIGNAL or_tmp_3107 : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_11_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_1_cse_6_sva_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL VEC_LOOP_j_sva_11_0 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_k_9_4_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_k_9_4_sva_2 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_12_1_1_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_19_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_13_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_10_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_14_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_16_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_6_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_17_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_8_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_12_sva : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_14_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_20_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL tmp_10_lpi_4_dfm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL mux_2770_m1c : STD_LOGIC;
  SIGNAL and_305_m1c : STD_LOGIC;
  SIGNAL and_307_m1c : STD_LOGIC;
  SIGNAL and_309_m1c : STD_LOGIC;
  SIGNAL and_312_m1c : STD_LOGIC;
  SIGNAL and_315_m1c : STD_LOGIC;
  SIGNAL and_317_m1c : STD_LOGIC;
  SIGNAL and_320_m1c : STD_LOGIC;
  SIGNAL and_322_m1c : STD_LOGIC;
  SIGNAL and_324_m1c : STD_LOGIC;
  SIGNAL and_327_m1c : STD_LOGIC;
  SIGNAL and_329_m1c : STD_LOGIC;
  SIGNAL and_331_m1c : STD_LOGIC;
  SIGNAL and_334_m1c : STD_LOGIC;
  SIGNAL and_336_m1c : STD_LOGIC;
  SIGNAL and_339_m1c : STD_LOGIC;
  SIGNAL and_300_m1c : STD_LOGIC;
  SIGNAL nor_223_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_0_15_obj_ld_cse : STD_LOGIC;
  SIGNAL and_574_cse : STD_LOGIC;
  SIGNAL or_2348_cse : STD_LOGIC;
  SIGNAL and_573_cse : STD_LOGIC;
  SIGNAL nand_375_cse : STD_LOGIC;
  SIGNAL or_495_cse : STD_LOGIC;
  SIGNAL nand_376_cse : STD_LOGIC;
  SIGNAL nor_412_cse : STD_LOGIC;
  SIGNAL and_563_cse : STD_LOGIC;
  SIGNAL or_2385_cse : STD_LOGIC;
  SIGNAL or_2894_cse : STD_LOGIC;
  SIGNAL and_517_cse : STD_LOGIC;
  SIGNAL and_528_cse : STD_LOGIC;
  SIGNAL and_565_cse : STD_LOGIC;
  SIGNAL and_456_cse : STD_LOGIC;
  SIGNAL and_458_cse : STD_LOGIC;
  SIGNAL or_3328_cse : STD_LOGIC;
  SIGNAL or_2520_cse : STD_LOGIC;
  SIGNAL nor_1203_cse : STD_LOGIC;
  SIGNAL or_2935_cse : STD_LOGIC;
  SIGNAL nand_398_cse : STD_LOGIC;
  SIGNAL or_2679_cse : STD_LOGIC;
  SIGNAL nor_381_cse : STD_LOGIC;
  SIGNAL nor_670_cse : STD_LOGIC;
  SIGNAL nand_237_cse : STD_LOGIC;
  SIGNAL modulo_result_mux_1_cse : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL nor_544_cse : STD_LOGIC;
  SIGNAL or_212_cse : STD_LOGIC;
  SIGNAL nor_422_cse : STD_LOGIC;
  SIGNAL and_472_cse : STD_LOGIC;
  SIGNAL and_491_cse : STD_LOGIC;
  SIGNAL and_816_cse : STD_LOGIC;
  SIGNAL mux_726_cse : STD_LOGIC;
  SIGNAL nor_601_cse : STD_LOGIC;
  SIGNAL nor_610_cse : STD_LOGIC;
  SIGNAL or_622_cse : STD_LOGIC;
  SIGNAL or_617_cse : STD_LOGIC;
  SIGNAL mux_1088_cse : STD_LOGIC;
  SIGNAL or_609_cse : STD_LOGIC;
  SIGNAL or_607_cse : STD_LOGIC;
  SIGNAL nand_25_cse : STD_LOGIC;
  SIGNAL or_601_cse : STD_LOGIC;
  SIGNAL mux_1073_cse : STD_LOGIC;
  SIGNAL or_2898_cse : STD_LOGIC;
  SIGNAL or_15_cse : STD_LOGIC;
  SIGNAL nor_784_cse : STD_LOGIC;
  SIGNAL or_2824_cse : STD_LOGIC;
  SIGNAL or_529_cse : STD_LOGIC;
  SIGNAL nand_226_cse : STD_LOGIC;
  SIGNAL or_2826_cse : STD_LOGIC;
  SIGNAL or_2839_cse : STD_LOGIC;
  SIGNAL nor_1276_cse : STD_LOGIC;
  SIGNAL nor_1279_cse : STD_LOGIC;
  SIGNAL and_459_cse : STD_LOGIC;
  SIGNAL and_440_cse : STD_LOGIC;
  SIGNAL nand_402_cse : STD_LOGIC;
  SIGNAL and_815_cse : STD_LOGIC;
  SIGNAL nor_539_cse : STD_LOGIC;
  SIGNAL mux_71_cse : STD_LOGIC;
  SIGNAL and_464_cse : STD_LOGIC;
  SIGNAL or_525_cse : STD_LOGIC;
  SIGNAL nand_240_cse : STD_LOGIC;
  SIGNAL mux_3498_cse : STD_LOGIC;
  SIGNAL or_154_cse : STD_LOGIC;
  SIGNAL or_2951_cse : STD_LOGIC;
  SIGNAL nor_1316_cse : STD_LOGIC;
  SIGNAL and_450_cse : STD_LOGIC;
  SIGNAL nor_515_cse : STD_LOGIC;
  SIGNAL mux_2746_cse : STD_LOGIC;
  SIGNAL or_3002_cse : STD_LOGIC;
  SIGNAL or_163_cse : STD_LOGIC;
  SIGNAL or_3308_cse : STD_LOGIC;
  SIGNAL or_3279_cse : STD_LOGIC;
  SIGNAL or_621_cse : STD_LOGIC;
  SIGNAL or_596_cse : STD_LOGIC;
  SIGNAL and_359_cse : STD_LOGIC;
  SIGNAL mux_3394_cse : STD_LOGIC;
  SIGNAL mux_3385_cse : STD_LOGIC;
  SIGNAL or_2729_cse : STD_LOGIC;
  SIGNAL and_754_cse : STD_LOGIC;
  SIGNAL mux_28_cse : STD_LOGIC;
  SIGNAL or_2902_cse : STD_LOGIC;
  SIGNAL or_36_cse : STD_LOGIC;
  SIGNAL or_2819_cse : STD_LOGIC;
  SIGNAL mux_3_cse : STD_LOGIC;
  SIGNAL mux_7_cse : STD_LOGIC;
  SIGNAL mux_9_cse : STD_LOGIC;
  SIGNAL mux_3143_cse : STD_LOGIC;
  SIGNAL mux_2463_cse : STD_LOGIC;
  SIGNAL mux_3603_cse : STD_LOGIC;
  SIGNAL nor_545_cse : STD_LOGIC;
  SIGNAL or_3018_cse : STD_LOGIC;
  SIGNAL or_3016_cse : STD_LOGIC;
  SIGNAL mux_3392_cse : STD_LOGIC;
  SIGNAL and_540_cse : STD_LOGIC;
  SIGNAL mux_3388_cse : STD_LOGIC;
  SIGNAL mux_384_cse : STD_LOGIC;
  SIGNAL mux_382_cse : STD_LOGIC;
  SIGNAL mux_3557_cse : STD_LOGIC;
  SIGNAL mux_3575_cse : STD_LOGIC;
  SIGNAL mux_3555_cse : STD_LOGIC;
  SIGNAL mux_3551_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_psp_sva_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL mux_2433_itm : STD_LOGIC;
  SIGNAL mux_2435_itm : STD_LOGIC;
  SIGNAL mux_2475_itm : STD_LOGIC;
  SIGNAL mux_3369_itm : STD_LOGIC;
  SIGNAL and_dcpl_348 : STD_LOGIC;
  SIGNAL and_dcpl_350 : STD_LOGIC;
  SIGNAL and_dcpl_351 : STD_LOGIC;
  SIGNAL and_dcpl_353 : STD_LOGIC;
  SIGNAL and_dcpl_354 : STD_LOGIC;
  SIGNAL and_dcpl_356 : STD_LOGIC;
  SIGNAL and_dcpl_358 : STD_LOGIC;
  SIGNAL and_dcpl_359 : STD_LOGIC;
  SIGNAL and_dcpl_361 : STD_LOGIC;
  SIGNAL and_dcpl_365 : STD_LOGIC;
  SIGNAL and_dcpl_368 : STD_LOGIC;
  SIGNAL and_dcpl_373 : STD_LOGIC;
  SIGNAL and_dcpl_374 : STD_LOGIC;
  SIGNAL and_dcpl_375 : STD_LOGIC;
  SIGNAL and_dcpl_376 : STD_LOGIC;
  SIGNAL and_dcpl_378 : STD_LOGIC;
  SIGNAL and_dcpl_380 : STD_LOGIC;
  SIGNAL and_dcpl_384 : STD_LOGIC;
  SIGNAL and_dcpl_386 : STD_LOGIC;
  SIGNAL and_dcpl_391 : STD_LOGIC;
  SIGNAL and_dcpl_392 : STD_LOGIC;
  SIGNAL and_dcpl_394 : STD_LOGIC;
  SIGNAL and_dcpl_397 : STD_LOGIC;
  SIGNAL and_dcpl_401 : STD_LOGIC;
  SIGNAL and_dcpl_404 : STD_LOGIC;
  SIGNAL and_dcpl_406 : STD_LOGIC;
  SIGNAL and_dcpl_408 : STD_LOGIC;
  SIGNAL and_dcpl_411 : STD_LOGIC;
  SIGNAL and_dcpl_415 : STD_LOGIC;
  SIGNAL z_out : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_430 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL and_dcpl_441 : STD_LOGIC;
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL and_dcpl_502 : STD_LOGIC;
  SIGNAL and_dcpl_503 : STD_LOGIC;
  SIGNAL and_dcpl_511 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_517 : STD_LOGIC;
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_555 : STD_LOGIC;
  SIGNAL not_tmp_930 : STD_LOGIC;
  SIGNAL mux_tmp : STD_LOGIC;
  SIGNAL not_tmp_933 : STD_LOGIC;
  SIGNAL and_dcpl_564 : STD_LOGIC;
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_dcpl_568 : STD_LOGIC;
  SIGNAL and_dcpl_574 : STD_LOGIC;
  SIGNAL or_tmp_3188 : STD_LOGIC;
  SIGNAL or_tmp_3189 : STD_LOGIC;
  SIGNAL mux_tmp_3724 : STD_LOGIC;
  SIGNAL or_tmp_3191 : STD_LOGIC;
  SIGNAL or_tmp_3193 : STD_LOGIC;
  SIGNAL mux_tmp_3725 : STD_LOGIC;
  SIGNAL or_tmp_3195 : STD_LOGIC;
  SIGNAL or_tmp_3196 : STD_LOGIC;
  SIGNAL mux_tmp_3728 : STD_LOGIC;
  SIGNAL or_tmp_3200 : STD_LOGIC;
  SIGNAL or_tmp_3202 : STD_LOGIC;
  SIGNAL or_tmp_3203 : STD_LOGIC;
  SIGNAL mux_tmp_3733 : STD_LOGIC;
  SIGNAL or_tmp_3204 : STD_LOGIC;
  SIGNAL or_tmp_3205 : STD_LOGIC;
  SIGNAL mux_tmp_3735 : STD_LOGIC;
  SIGNAL mux_tmp_3737 : STD_LOGIC;
  SIGNAL or_tmp_3211 : STD_LOGIC;
  SIGNAL mux_tmp_3742 : STD_LOGIC;
  SIGNAL or_tmp_3212 : STD_LOGIC;
  SIGNAL mux_tmp_3743 : STD_LOGIC;
  SIGNAL or_tmp_3213 : STD_LOGIC;
  SIGNAL or_tmp_3218 : STD_LOGIC;
  SIGNAL mux_tmp_3751 : STD_LOGIC;
  SIGNAL mux_tmp_3753 : STD_LOGIC;
  SIGNAL mux_tmp_3762 : STD_LOGIC;
  SIGNAL mux_tmp_3771 : STD_LOGIC;
  SIGNAL and_dcpl_579 : STD_LOGIC;
  SIGNAL and_dcpl_588 : STD_LOGIC;
  SIGNAL z_out_6 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL and_dcpl_591 : STD_LOGIC;
  SIGNAL and_dcpl_592 : STD_LOGIC;
  SIGNAL and_dcpl_598 : STD_LOGIC;
  SIGNAL and_dcpl_614 : STD_LOGIC;
  SIGNAL and_dcpl_615 : STD_LOGIC;
  SIGNAL and_dcpl_618 : STD_LOGIC;
  SIGNAL and_dcpl_622 : STD_LOGIC;
  SIGNAL and_dcpl_623 : STD_LOGIC;
  SIGNAL and_dcpl_624 : STD_LOGIC;
  SIGNAL and_dcpl_628 : STD_LOGIC;
  SIGNAL and_dcpl_641 : STD_LOGIC;
  SIGNAL and_dcpl_642 : STD_LOGIC;
  SIGNAL and_dcpl_646 : STD_LOGIC;
  SIGNAL and_dcpl_651 : STD_LOGIC;
  SIGNAL and_dcpl_654 : STD_LOGIC;
  SIGNAL and_dcpl_657 : STD_LOGIC;
  SIGNAL and_dcpl_659 : STD_LOGIC;
  SIGNAL and_dcpl_663 : STD_LOGIC;
  SIGNAL and_dcpl_666 : STD_LOGIC;
  SIGNAL and_dcpl_669 : STD_LOGIC;
  SIGNAL and_dcpl_672 : STD_LOGIC;
  SIGNAL and_dcpl_676 : STD_LOGIC;
  SIGNAL and_dcpl_678 : STD_LOGIC;
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL and_dcpl_688 : STD_LOGIC;
  SIGNAL and_dcpl_698 : STD_LOGIC;
  SIGNAL not_tmp_980 : STD_LOGIC;
  SIGNAL and_dcpl_707 : STD_LOGIC;
  SIGNAL and_dcpl_717 : STD_LOGIC;
  SIGNAL and_dcpl_727 : STD_LOGIC;
  SIGNAL and_dcpl_734 : STD_LOGIC;
  SIGNAL and_dcpl_741 : STD_LOGIC;
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL z_out_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL modExp_result_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_exp_1_7_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_6_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_5_1_sva : STD_LOGIC;
  SIGNAL modExp_exp_1_4_1_sva : STD_LOGIC;
  SIGNAL COMP_LOOP_10_mul_mut : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_2_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_4_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_8_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_11_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_62_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_64_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_68_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_139_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_141_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_143_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_144_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_145_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_146_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_147_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_148_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_149_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_134_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_305_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_10_acc_8_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva_mx0c1 : STD_LOGIC;
  SIGNAL STAGE_LOOP_i_3_0_sva_2 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modExp_1_while_if_mul_mut_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL VEC_LOOP_j_sva_11_0_mx0c1 : STD_LOGIC;
  SIGNAL modExp_result_sva_mx0c0 : STD_LOGIC;
  SIGNAL operator_64_false_slc_modExp_exp_63_1_3 : STD_LOGIC_VECTOR (62 DOWNTO 0);
  SIGNAL modExp_while_and_3 : STD_LOGIC;
  SIGNAL modExp_while_and_5 : STD_LOGIC;
  SIGNAL and_345_m1c : STD_LOGIC;
  SIGNAL modExp_result_and_rgt : STD_LOGIC;
  SIGNAL modExp_result_and_1_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_or_32_cse : STD_LOGIC;
  SIGNAL nor_1148_cse : STD_LOGIC;
  SIGNAL or_642_cse : STD_LOGIC;
  SIGNAL nor_1123_cse : STD_LOGIC;
  SIGNAL or_748_cse : STD_LOGIC;
  SIGNAL nor_1098_cse : STD_LOGIC;
  SIGNAL or_855_cse : STD_LOGIC;
  SIGNAL nor_1073_cse : STD_LOGIC;
  SIGNAL or_961_cse : STD_LOGIC;
  SIGNAL nor_1048_cse : STD_LOGIC;
  SIGNAL or_1068_cse : STD_LOGIC;
  SIGNAL nor_1023_cse : STD_LOGIC;
  SIGNAL or_1174_cse : STD_LOGIC;
  SIGNAL nor_998_cse : STD_LOGIC;
  SIGNAL or_1281_cse : STD_LOGIC;
  SIGNAL nor_975_cse : STD_LOGIC;
  SIGNAL or_1387_cse : STD_LOGIC;
  SIGNAL nor_950_cse : STD_LOGIC;
  SIGNAL or_1494_cse : STD_LOGIC;
  SIGNAL nor_925_cse : STD_LOGIC;
  SIGNAL or_1600_cse : STD_LOGIC;
  SIGNAL nor_900_cse : STD_LOGIC;
  SIGNAL or_1707_cse : STD_LOGIC;
  SIGNAL nor_877_cse : STD_LOGIC;
  SIGNAL or_1813_cse : STD_LOGIC;
  SIGNAL nor_850_cse : STD_LOGIC;
  SIGNAL or_1923_cse : STD_LOGIC;
  SIGNAL nor_827_cse : STD_LOGIC;
  SIGNAL or_2029_cse : STD_LOGIC;
  SIGNAL nor_804_cse : STD_LOGIC;
  SIGNAL or_2136_cse : STD_LOGIC;
  SIGNAL and_591_cse : STD_LOGIC;
  SIGNAL nand_278_cse : STD_LOGIC;
  SIGNAL nand_257_cse : STD_LOGIC;
  SIGNAL nor_738_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_55_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_or_56_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_or_57_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_or_58_ssc : STD_LOGIC;
  SIGNAL and_850_cse : STD_LOGIC;
  SIGNAL and_857_cse : STD_LOGIC;
  SIGNAL and_869_cse : STD_LOGIC;
  SIGNAL and_875_cse : STD_LOGIC;
  SIGNAL and_886_cse : STD_LOGIC;
  SIGNAL or_tmp : STD_LOGIC;
  SIGNAL nor_tmp : STD_LOGIC;
  SIGNAL mux_tmp_3818 : STD_LOGIC;
  SIGNAL not_tmp_1007 : STD_LOGIC;
  SIGNAL mux_tmp_3819 : STD_LOGIC;
  SIGNAL mux_tmp_3822 : STD_LOGIC;
  SIGNAL or_tmp_3291 : STD_LOGIC;
  SIGNAL or_tmp_3293 : STD_LOGIC;
  SIGNAL nor_tmp_535 : STD_LOGIC;
  SIGNAL nor_tmp_536 : STD_LOGIC;
  SIGNAL mux_tmp_3828 : STD_LOGIC;
  SIGNAL mux_tmp_3834 : STD_LOGIC;
  SIGNAL nor_tmp_539 : STD_LOGIC;
  SIGNAL nor_tmp_540 : STD_LOGIC;
  SIGNAL or_tmp_3303 : STD_LOGIC;
  SIGNAL or_tmp_3304 : STD_LOGIC;
  SIGNAL mux_tmp_3846 : STD_LOGIC;
  SIGNAL mux_tmp_3853 : STD_LOGIC;
  SIGNAL not_tmp_1021 : STD_LOGIC;
  SIGNAL mux_tmp_3861 : STD_LOGIC;
  SIGNAL mux_tmp_3878 : STD_LOGIC;
  SIGNAL or_tmp_3320 : STD_LOGIC;
  SIGNAL not_tmp_1034 : STD_LOGIC;
  SIGNAL or_tmp_3327 : STD_LOGIC;
  SIGNAL mux_tmp_3898 : STD_LOGIC;
  SIGNAL or_tmp_3332 : STD_LOGIC;
  SIGNAL nand_tmp : STD_LOGIC;
  SIGNAL mux_tmp_3902 : STD_LOGIC;
  SIGNAL mux_tmp_3906 : STD_LOGIC;
  SIGNAL or_tmp_3343 : STD_LOGIC;
  SIGNAL mux_tmp_3915 : STD_LOGIC;
  SIGNAL or_tmp_3369 : STD_LOGIC;
  SIGNAL operator_64_false_mux1h_2_rgt : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_64_false_acc_mut_64 : STD_LOGIC;
  SIGNAL operator_64_false_acc_mut_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_1262_cse : STD_LOGIC;
  SIGNAL nor_1450_cse : STD_LOGIC;
  SIGNAL or_2747_cse : STD_LOGIC;
  SIGNAL nand_201_cse : STD_LOGIC;
  SIGNAL or_2415_cse : STD_LOGIC;
  SIGNAL or_3280_cse : STD_LOGIC;
  SIGNAL mux_3724_itm : STD_LOGIC;
  SIGNAL mux_3788_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_60_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_24_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_67_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_680_itm : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_itm_2_1 : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_6_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_9_cse : STD_LOGIC;
  SIGNAL z_out_8_8_7 : STD_LOGIC_VECTOR (1 DOWNTO 0);

  SIGNAL mux_1092_nl : STD_LOGIC;
  SIGNAL nand_360_nl : STD_LOGIC;
  SIGNAL or_619_nl : STD_LOGIC;
  SIGNAL modulo_result_or_nl : STD_LOGIC;
  SIGNAL mux_2303_nl : STD_LOGIC;
  SIGNAL mux_2302_nl : STD_LOGIC;
  SIGNAL mux_2301_nl : STD_LOGIC;
  SIGNAL mux_2300_nl : STD_LOGIC;
  SIGNAL mux_2299_nl : STD_LOGIC;
  SIGNAL mux_2298_nl : STD_LOGIC;
  SIGNAL mux_2297_nl : STD_LOGIC;
  SIGNAL mux_2296_nl : STD_LOGIC;
  SIGNAL mux_2295_nl : STD_LOGIC;
  SIGNAL mux_2294_nl : STD_LOGIC;
  SIGNAL mux_2293_nl : STD_LOGIC;
  SIGNAL mux_2292_nl : STD_LOGIC;
  SIGNAL mux_2291_nl : STD_LOGIC;
  SIGNAL nand_264_nl : STD_LOGIC;
  SIGNAL mux_2288_nl : STD_LOGIC;
  SIGNAL mux_2287_nl : STD_LOGIC;
  SIGNAL mux_2286_nl : STD_LOGIC;
  SIGNAL mux_2284_nl : STD_LOGIC;
  SIGNAL mux_2283_nl : STD_LOGIC;
  SIGNAL mux_2282_nl : STD_LOGIC;
  SIGNAL mux_2281_nl : STD_LOGIC;
  SIGNAL mux_2280_nl : STD_LOGIC;
  SIGNAL mux_2278_nl : STD_LOGIC;
  SIGNAL mux_2277_nl : STD_LOGIC;
  SIGNAL nand_265_nl : STD_LOGIC;
  SIGNAL mux_2276_nl : STD_LOGIC;
  SIGNAL mux_2275_nl : STD_LOGIC;
  SIGNAL mux_2274_nl : STD_LOGIC;
  SIGNAL mux_2273_nl : STD_LOGIC;
  SIGNAL mux_2272_nl : STD_LOGIC;
  SIGNAL mux_2271_nl : STD_LOGIC;
  SIGNAL mux_2270_nl : STD_LOGIC;
  SIGNAL mux_2269_nl : STD_LOGIC;
  SIGNAL mux_2268_nl : STD_LOGIC;
  SIGNAL mux_2267_nl : STD_LOGIC;
  SIGNAL mux_2266_nl : STD_LOGIC;
  SIGNAL mux_2264_nl : STD_LOGIC;
  SIGNAL mux_2263_nl : STD_LOGIC;
  SIGNAL mux_2262_nl : STD_LOGIC;
  SIGNAL nor_778_nl : STD_LOGIC;
  SIGNAL mux_2261_nl : STD_LOGIC;
  SIGNAL mux_2260_nl : STD_LOGIC;
  SIGNAL mux_2259_nl : STD_LOGIC;
  SIGNAL mux_2258_nl : STD_LOGIC;
  SIGNAL mux_2257_nl : STD_LOGIC;
  SIGNAL mux_2256_nl : STD_LOGIC;
  SIGNAL nor_779_nl : STD_LOGIC;
  SIGNAL mux_2255_nl : STD_LOGIC;
  SIGNAL mux_2253_nl : STD_LOGIC;
  SIGNAL mux_2252_nl : STD_LOGIC;
  SIGNAL mux_2249_nl : STD_LOGIC;
  SIGNAL mux_2248_nl : STD_LOGIC;
  SIGNAL mux_2247_nl : STD_LOGIC;
  SIGNAL mux_2246_nl : STD_LOGIC;
  SIGNAL or_2306_nl : STD_LOGIC;
  SIGNAL mux_2245_nl : STD_LOGIC;
  SIGNAL mux_2244_nl : STD_LOGIC;
  SIGNAL mux_2243_nl : STD_LOGIC;
  SIGNAL mux_2242_nl : STD_LOGIC;
  SIGNAL mux_2241_nl : STD_LOGIC;
  SIGNAL mux_2238_nl : STD_LOGIC;
  SIGNAL mux_2237_nl : STD_LOGIC;
  SIGNAL mux_2236_nl : STD_LOGIC;
  SIGNAL mux_2235_nl : STD_LOGIC;
  SIGNAL or_2300_nl : STD_LOGIC;
  SIGNAL nand_91_nl : STD_LOGIC;
  SIGNAL mux_2234_nl : STD_LOGIC;
  SIGNAL or_2297_nl : STD_LOGIC;
  SIGNAL mux_2233_nl : STD_LOGIC;
  SIGNAL mux_2232_nl : STD_LOGIC;
  SIGNAL or_2293_nl : STD_LOGIC;
  SIGNAL mux_2231_nl : STD_LOGIC;
  SIGNAL mux_2230_nl : STD_LOGIC;
  SIGNAL mux_2229_nl : STD_LOGIC;
  SIGNAL mux_2228_nl : STD_LOGIC;
  SIGNAL mux_2227_nl : STD_LOGIC;
  SIGNAL mux_2226_nl : STD_LOGIC;
  SIGNAL mux_2225_nl : STD_LOGIC;
  SIGNAL mux_2224_nl : STD_LOGIC;
  SIGNAL mux_2222_nl : STD_LOGIC;
  SIGNAL mux_2221_nl : STD_LOGIC;
  SIGNAL mux_2219_nl : STD_LOGIC;
  SIGNAL or_2288_nl : STD_LOGIC;
  SIGNAL mux_2217_nl : STD_LOGIC;
  SIGNAL mux_2216_nl : STD_LOGIC;
  SIGNAL mux_2215_nl : STD_LOGIC;
  SIGNAL or_2285_nl : STD_LOGIC;
  SIGNAL or_2283_nl : STD_LOGIC;
  SIGNAL mux_2214_nl : STD_LOGIC;
  SIGNAL mux_2213_nl : STD_LOGIC;
  SIGNAL mux_2212_nl : STD_LOGIC;
  SIGNAL or_2279_nl : STD_LOGIC;
  SIGNAL mux_2211_nl : STD_LOGIC;
  SIGNAL nand_90_nl : STD_LOGIC;
  SIGNAL mux_2378_nl : STD_LOGIC;
  SIGNAL mux_2377_nl : STD_LOGIC;
  SIGNAL mux_2376_nl : STD_LOGIC;
  SIGNAL mux_2375_nl : STD_LOGIC;
  SIGNAL mux_2374_nl : STD_LOGIC;
  SIGNAL mux_2373_nl : STD_LOGIC;
  SIGNAL or_2355_nl : STD_LOGIC;
  SIGNAL mux_2372_nl : STD_LOGIC;
  SIGNAL mux_2371_nl : STD_LOGIC;
  SIGNAL mux_2370_nl : STD_LOGIC;
  SIGNAL mux_2369_nl : STD_LOGIC;
  SIGNAL or_2354_nl : STD_LOGIC;
  SIGNAL mux_2368_nl : STD_LOGIC;
  SIGNAL or_2351_nl : STD_LOGIC;
  SIGNAL mux_2367_nl : STD_LOGIC;
  SIGNAL mux_2366_nl : STD_LOGIC;
  SIGNAL mux_2365_nl : STD_LOGIC;
  SIGNAL mux_2364_nl : STD_LOGIC;
  SIGNAL mux_2363_nl : STD_LOGIC;
  SIGNAL nand_100_nl : STD_LOGIC;
  SIGNAL mux_2361_nl : STD_LOGIC;
  SIGNAL mux_2360_nl : STD_LOGIC;
  SIGNAL nand_99_nl : STD_LOGIC;
  SIGNAL mux_2359_nl : STD_LOGIC;
  SIGNAL nand_98_nl : STD_LOGIC;
  SIGNAL mux_2358_nl : STD_LOGIC;
  SIGNAL mux_2357_nl : STD_LOGIC;
  SIGNAL mux_2356_nl : STD_LOGIC;
  SIGNAL mux_2355_nl : STD_LOGIC;
  SIGNAL mux_2354_nl : STD_LOGIC;
  SIGNAL mux_2353_nl : STD_LOGIC;
  SIGNAL mux_2352_nl : STD_LOGIC;
  SIGNAL mux_2351_nl : STD_LOGIC;
  SIGNAL mux_2350_nl : STD_LOGIC;
  SIGNAL mux_2348_nl : STD_LOGIC;
  SIGNAL nand_261_nl : STD_LOGIC;
  SIGNAL mux_2347_nl : STD_LOGIC;
  SIGNAL and_275_nl : STD_LOGIC;
  SIGNAL mux_2346_nl : STD_LOGIC;
  SIGNAL mux_2345_nl : STD_LOGIC;
  SIGNAL mux_2344_nl : STD_LOGIC;
  SIGNAL mux_2343_nl : STD_LOGIC;
  SIGNAL or_2343_nl : STD_LOGIC;
  SIGNAL mux_2342_nl : STD_LOGIC;
  SIGNAL or_2342_nl : STD_LOGIC;
  SIGNAL mux_2341_nl : STD_LOGIC;
  SIGNAL mux_2340_nl : STD_LOGIC;
  SIGNAL nand_262_nl : STD_LOGIC;
  SIGNAL mux_2339_nl : STD_LOGIC;
  SIGNAL or_2341_nl : STD_LOGIC;
  SIGNAL mux_2338_nl : STD_LOGIC;
  SIGNAL mux_2337_nl : STD_LOGIC;
  SIGNAL mux_2336_nl : STD_LOGIC;
  SIGNAL mux_2335_nl : STD_LOGIC;
  SIGNAL mux_2334_nl : STD_LOGIC;
  SIGNAL mux_2333_nl : STD_LOGIC;
  SIGNAL mux_2332_nl : STD_LOGIC;
  SIGNAL mux_2331_nl : STD_LOGIC;
  SIGNAL mux_2330_nl : STD_LOGIC;
  SIGNAL mux_2329_nl : STD_LOGIC;
  SIGNAL mux_2328_nl : STD_LOGIC;
  SIGNAL mux_2326_nl : STD_LOGIC;
  SIGNAL mux_2325_nl : STD_LOGIC;
  SIGNAL mux_2324_nl : STD_LOGIC;
  SIGNAL mux_2323_nl : STD_LOGIC;
  SIGNAL nand_97_nl : STD_LOGIC;
  SIGNAL mux_2322_nl : STD_LOGIC;
  SIGNAL mux_2321_nl : STD_LOGIC;
  SIGNAL mux_2320_nl : STD_LOGIC;
  SIGNAL mux_2319_nl : STD_LOGIC;
  SIGNAL mux_2318_nl : STD_LOGIC;
  SIGNAL mux_2317_nl : STD_LOGIC;
  SIGNAL mux_2316_nl : STD_LOGIC;
  SIGNAL mux_2315_nl : STD_LOGIC;
  SIGNAL mux_2314_nl : STD_LOGIC;
  SIGNAL or_2330_nl : STD_LOGIC;
  SIGNAL or_2329_nl : STD_LOGIC;
  SIGNAL mux_2313_nl : STD_LOGIC;
  SIGNAL mux_2312_nl : STD_LOGIC;
  SIGNAL mux_2311_nl : STD_LOGIC;
  SIGNAL mux_2308_nl : STD_LOGIC;
  SIGNAL nand_94_nl : STD_LOGIC;
  SIGNAL mux_2307_nl : STD_LOGIC;
  SIGNAL mux_2306_nl : STD_LOGIC;
  SIGNAL mux_2305_nl : STD_LOGIC;
  SIGNAL or_2321_nl : STD_LOGIC;
  SIGNAL mux_2304_nl : STD_LOGIC;
  SIGNAL or_2319_nl : STD_LOGIC;
  SIGNAL mux_2394_nl : STD_LOGIC;
  SIGNAL mux_2393_nl : STD_LOGIC;
  SIGNAL mux_2392_nl : STD_LOGIC;
  SIGNAL mux_2391_nl : STD_LOGIC;
  SIGNAL nor_758_nl : STD_LOGIC;
  SIGNAL nor_759_nl : STD_LOGIC;
  SIGNAL and_568_nl : STD_LOGIC;
  SIGNAL mux_2390_nl : STD_LOGIC;
  SIGNAL nor_760_nl : STD_LOGIC;
  SIGNAL nor_761_nl : STD_LOGIC;
  SIGNAL mux_2389_nl : STD_LOGIC;
  SIGNAL mux_2388_nl : STD_LOGIC;
  SIGNAL nor_762_nl : STD_LOGIC;
  SIGNAL nor_763_nl : STD_LOGIC;
  SIGNAL nor_764_nl : STD_LOGIC;
  SIGNAL mux_2387_nl : STD_LOGIC;
  SIGNAL or_2372_nl : STD_LOGIC;
  SIGNAL or_2370_nl : STD_LOGIC;
  SIGNAL mux_2386_nl : STD_LOGIC;
  SIGNAL and_569_nl : STD_LOGIC;
  SIGNAL mux_2385_nl : STD_LOGIC;
  SIGNAL and_570_nl : STD_LOGIC;
  SIGNAL mux_2384_nl : STD_LOGIC;
  SIGNAL nor_765_nl : STD_LOGIC;
  SIGNAL nor_766_nl : STD_LOGIC;
  SIGNAL nor_767_nl : STD_LOGIC;
  SIGNAL mux_2383_nl : STD_LOGIC;
  SIGNAL or_2365_nl : STD_LOGIC;
  SIGNAL or_2364_nl : STD_LOGIC;
  SIGNAL mux_2382_nl : STD_LOGIC;
  SIGNAL mux_2381_nl : STD_LOGIC;
  SIGNAL nor_768_nl : STD_LOGIC;
  SIGNAL mux_2380_nl : STD_LOGIC;
  SIGNAL mux_2379_nl : STD_LOGIC;
  SIGNAL nor_769_nl : STD_LOGIC;
  SIGNAL nor_770_nl : STD_LOGIC;
  SIGNAL nor_771_nl : STD_LOGIC;
  SIGNAL nor_772_nl : STD_LOGIC;
  SIGNAL mux_2461_nl : STD_LOGIC;
  SIGNAL mux_2460_nl : STD_LOGIC;
  SIGNAL mux_2459_nl : STD_LOGIC;
  SIGNAL mux_2458_nl : STD_LOGIC;
  SIGNAL mux_2457_nl : STD_LOGIC;
  SIGNAL mux_2456_nl : STD_LOGIC;
  SIGNAL nand_109_nl : STD_LOGIC;
  SIGNAL mux_2455_nl : STD_LOGIC;
  SIGNAL mux_2454_nl : STD_LOGIC;
  SIGNAL mux_2453_nl : STD_LOGIC;
  SIGNAL mux_2452_nl : STD_LOGIC;
  SIGNAL mux_2451_nl : STD_LOGIC;
  SIGNAL mux_2450_nl : STD_LOGIC;
  SIGNAL mux_2449_nl : STD_LOGIC;
  SIGNAL mux_2448_nl : STD_LOGIC;
  SIGNAL mux_2447_nl : STD_LOGIC;
  SIGNAL mux_2446_nl : STD_LOGIC;
  SIGNAL mux_2445_nl : STD_LOGIC;
  SIGNAL mux_2444_nl : STD_LOGIC;
  SIGNAL mux_2443_nl : STD_LOGIC;
  SIGNAL mux_2442_nl : STD_LOGIC;
  SIGNAL mux_2441_nl : STD_LOGIC;
  SIGNAL mux_2440_nl : STD_LOGIC;
  SIGNAL mux_2439_nl : STD_LOGIC;
  SIGNAL mux_2438_nl : STD_LOGIC;
  SIGNAL mux_2437_nl : STD_LOGIC;
  SIGNAL mux_2434_nl : STD_LOGIC;
  SIGNAL mux_2432_nl : STD_LOGIC;
  SIGNAL mux_2431_nl : STD_LOGIC;
  SIGNAL mux_2430_nl : STD_LOGIC;
  SIGNAL mux_2429_nl : STD_LOGIC;
  SIGNAL mux_2428_nl : STD_LOGIC;
  SIGNAL mux_2424_nl : STD_LOGIC;
  SIGNAL nand_106_nl : STD_LOGIC;
  SIGNAL mux_2421_nl : STD_LOGIC;
  SIGNAL mux_2420_nl : STD_LOGIC;
  SIGNAL mux_2419_nl : STD_LOGIC;
  SIGNAL mux_2418_nl : STD_LOGIC;
  SIGNAL mux_2417_nl : STD_LOGIC;
  SIGNAL mux_2416_nl : STD_LOGIC;
  SIGNAL or_2397_nl : STD_LOGIC;
  SIGNAL mux_2415_nl : STD_LOGIC;
  SIGNAL mux_2414_nl : STD_LOGIC;
  SIGNAL mux_2413_nl : STD_LOGIC;
  SIGNAL mux_2412_nl : STD_LOGIC;
  SIGNAL mux_2411_nl : STD_LOGIC;
  SIGNAL mux_2410_nl : STD_LOGIC;
  SIGNAL mux_2409_nl : STD_LOGIC;
  SIGNAL mux_2408_nl : STD_LOGIC;
  SIGNAL mux_2407_nl : STD_LOGIC;
  SIGNAL mux_2405_nl : STD_LOGIC;
  SIGNAL mux_2404_nl : STD_LOGIC;
  SIGNAL mux_2403_nl : STD_LOGIC;
  SIGNAL mux_2399_nl : STD_LOGIC;
  SIGNAL mux_2398_nl : STD_LOGIC;
  SIGNAL mux_2397_nl : STD_LOGIC;
  SIGNAL mux_2396_nl : STD_LOGIC;
  SIGNAL nand_104_nl : STD_LOGIC;
  SIGNAL mux_2395_nl : STD_LOGIC;
  SIGNAL or_2381_nl : STD_LOGIC;
  SIGNAL mux_2495_nl : STD_LOGIC;
  SIGNAL mux_2494_nl : STD_LOGIC;
  SIGNAL mux_2493_nl : STD_LOGIC;
  SIGNAL or_3297_nl : STD_LOGIC;
  SIGNAL nand_250_nl : STD_LOGIC;
  SIGNAL or_2778_nl : STD_LOGIC;
  SIGNAL modExp_while_if_mux1h_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_353_nl : STD_LOGIC;
  SIGNAL mux_3149_nl : STD_LOGIC;
  SIGNAL mux_3148_nl : STD_LOGIC;
  SIGNAL mux_3147_nl : STD_LOGIC;
  SIGNAL mux_3146_nl : STD_LOGIC;
  SIGNAL and_466_nl : STD_LOGIC;
  SIGNAL mux_3145_nl : STD_LOGIC;
  SIGNAL nor_637_nl : STD_LOGIC;
  SIGNAL nor_638_nl : STD_LOGIC;
  SIGNAL nor_639_nl : STD_LOGIC;
  SIGNAL and_467_nl : STD_LOGIC;
  SIGNAL and_468_nl : STD_LOGIC;
  SIGNAL mux_3144_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL nor_641_nl : STD_LOGIC;
  SIGNAL mux_3142_nl : STD_LOGIC;
  SIGNAL mux_3141_nl : STD_LOGIC;
  SIGNAL mux_3140_nl : STD_LOGIC;
  SIGNAL nor_642_nl : STD_LOGIC;
  SIGNAL and_469_nl : STD_LOGIC;
  SIGNAL nor_643_nl : STD_LOGIC;
  SIGNAL mux_3139_nl : STD_LOGIC;
  SIGNAL mux_3138_nl : STD_LOGIC;
  SIGNAL or_2773_nl : STD_LOGIC;
  SIGNAL or_2772_nl : STD_LOGIC;
  SIGNAL or_2771_nl : STD_LOGIC;
  SIGNAL mux_3137_nl : STD_LOGIC;
  SIGNAL or_2770_nl : STD_LOGIC;
  SIGNAL and_470_nl : STD_LOGIC;
  SIGNAL mux_3136_nl : STD_LOGIC;
  SIGNAL nor_644_nl : STD_LOGIC;
  SIGNAL mux_3135_nl : STD_LOGIC;
  SIGNAL nor_645_nl : STD_LOGIC;
  SIGNAL modExp_while_if_and_nl : STD_LOGIC;
  SIGNAL modExp_while_if_and_1_nl : STD_LOGIC;
  SIGNAL and_284_nl : STD_LOGIC;
  SIGNAL mux_2566_nl : STD_LOGIC;
  SIGNAL mux_2565_nl : STD_LOGIC;
  SIGNAL mux_2564_nl : STD_LOGIC;
  SIGNAL mux_2563_nl : STD_LOGIC;
  SIGNAL mux_2562_nl : STD_LOGIC;
  SIGNAL mux_2561_nl : STD_LOGIC;
  SIGNAL mux_2560_nl : STD_LOGIC;
  SIGNAL mux_2559_nl : STD_LOGIC;
  SIGNAL mux_2558_nl : STD_LOGIC;
  SIGNAL and_532_nl : STD_LOGIC;
  SIGNAL and_533_nl : STD_LOGIC;
  SIGNAL mux_2557_nl : STD_LOGIC;
  SIGNAL or_2494_nl : STD_LOGIC;
  SIGNAL mux_2556_nl : STD_LOGIC;
  SIGNAL mux_2555_nl : STD_LOGIC;
  SIGNAL mux_2554_nl : STD_LOGIC;
  SIGNAL mux_2553_nl : STD_LOGIC;
  SIGNAL and_535_nl : STD_LOGIC;
  SIGNAL or_2491_nl : STD_LOGIC;
  SIGNAL mux_2552_nl : STD_LOGIC;
  SIGNAL mux_2551_nl : STD_LOGIC;
  SIGNAL mux_2550_nl : STD_LOGIC;
  SIGNAL mux_2548_nl : STD_LOGIC;
  SIGNAL nor_731_nl : STD_LOGIC;
  SIGNAL mux_2547_nl : STD_LOGIC;
  SIGNAL mux_2546_nl : STD_LOGIC;
  SIGNAL mux_2545_nl : STD_LOGIC;
  SIGNAL mux_2544_nl : STD_LOGIC;
  SIGNAL mux_2543_nl : STD_LOGIC;
  SIGNAL mux_2542_nl : STD_LOGIC;
  SIGNAL mux_2541_nl : STD_LOGIC;
  SIGNAL or_2484_nl : STD_LOGIC;
  SIGNAL mux_2540_nl : STD_LOGIC;
  SIGNAL mux_2539_nl : STD_LOGIC;
  SIGNAL mux_2538_nl : STD_LOGIC;
  SIGNAL or_2483_nl : STD_LOGIC;
  SIGNAL mux_2537_nl : STD_LOGIC;
  SIGNAL mux_2536_nl : STD_LOGIC;
  SIGNAL mux_2535_nl : STD_LOGIC;
  SIGNAL nor_732_nl : STD_LOGIC;
  SIGNAL mux_2534_nl : STD_LOGIC;
  SIGNAL or_2480_nl : STD_LOGIC;
  SIGNAL mux_2533_nl : STD_LOGIC;
  SIGNAL mux_2532_nl : STD_LOGIC;
  SIGNAL mux_2531_nl : STD_LOGIC;
  SIGNAL mux_2530_nl : STD_LOGIC;
  SIGNAL mux_2529_nl : STD_LOGIC;
  SIGNAL mux_2528_nl : STD_LOGIC;
  SIGNAL mux_2527_nl : STD_LOGIC;
  SIGNAL mux_2526_nl : STD_LOGIC;
  SIGNAL mux_2524_nl : STD_LOGIC;
  SIGNAL mux_2522_nl : STD_LOGIC;
  SIGNAL mux_2521_nl : STD_LOGIC;
  SIGNAL nor_733_nl : STD_LOGIC;
  SIGNAL mux_2520_nl : STD_LOGIC;
  SIGNAL mux_2518_nl : STD_LOGIC;
  SIGNAL mux_2517_nl : STD_LOGIC;
  SIGNAL mux_2516_nl : STD_LOGIC;
  SIGNAL mux_2515_nl : STD_LOGIC;
  SIGNAL or_2475_nl : STD_LOGIC;
  SIGNAL mux_2514_nl : STD_LOGIC;
  SIGNAL mux_2513_nl : STD_LOGIC;
  SIGNAL or_2472_nl : STD_LOGIC;
  SIGNAL mux_2512_nl : STD_LOGIC;
  SIGNAL mux_2511_nl : STD_LOGIC;
  SIGNAL mux_2510_nl : STD_LOGIC;
  SIGNAL mux_2509_nl : STD_LOGIC;
  SIGNAL mux_2507_nl : STD_LOGIC;
  SIGNAL or_2466_nl : STD_LOGIC;
  SIGNAL mux_2506_nl : STD_LOGIC;
  SIGNAL mux_2505_nl : STD_LOGIC;
  SIGNAL mux_2504_nl : STD_LOGIC;
  SIGNAL mux_2503_nl : STD_LOGIC;
  SIGNAL or_2460_nl : STD_LOGIC;
  SIGNAL mux_2500_nl : STD_LOGIC;
  SIGNAL and_544_nl : STD_LOGIC;
  SIGNAL mux_2499_nl : STD_LOGIC;
  SIGNAL mux_2498_nl : STD_LOGIC;
  SIGNAL nand_247_nl : STD_LOGIC;
  SIGNAL mux_2497_nl : STD_LOGIC;
  SIGNAL nand_248_nl : STD_LOGIC;
  SIGNAL or_2454_nl : STD_LOGIC;
  SIGNAL mux_3896_nl : STD_LOGIC;
  SIGNAL mux_3895_nl : STD_LOGIC;
  SIGNAL mux_3894_nl : STD_LOGIC;
  SIGNAL mux_3893_nl : STD_LOGIC;
  SIGNAL mux_3892_nl : STD_LOGIC;
  SIGNAL mux_3891_nl : STD_LOGIC;
  SIGNAL mux_3890_nl : STD_LOGIC;
  SIGNAL nor_1453_nl : STD_LOGIC;
  SIGNAL mux_3889_nl : STD_LOGIC;
  SIGNAL mux_3888_nl : STD_LOGIC;
  SIGNAL mux_3887_nl : STD_LOGIC;
  SIGNAL and_1258_nl : STD_LOGIC;
  SIGNAL mux_3886_nl : STD_LOGIC;
  SIGNAL or_3508_nl : STD_LOGIC;
  SIGNAL mux_3885_nl : STD_LOGIC;
  SIGNAL mux_3884_nl : STD_LOGIC;
  SIGNAL and_1259_nl : STD_LOGIC;
  SIGNAL mux_3883_nl : STD_LOGIC;
  SIGNAL mux_3882_nl : STD_LOGIC;
  SIGNAL mux_3881_nl : STD_LOGIC;
  SIGNAL and_1260_nl : STD_LOGIC;
  SIGNAL mux_3880_nl : STD_LOGIC;
  SIGNAL or_3506_nl : STD_LOGIC;
  SIGNAL mux_3878_nl : STD_LOGIC;
  SIGNAL mux_3877_nl : STD_LOGIC;
  SIGNAL mux_3876_nl : STD_LOGIC;
  SIGNAL mux_3875_nl : STD_LOGIC;
  SIGNAL or_3505_nl : STD_LOGIC;
  SIGNAL mux_3874_nl : STD_LOGIC;
  SIGNAL or_3504_nl : STD_LOGIC;
  SIGNAL mux_3873_nl : STD_LOGIC;
  SIGNAL and_1256_nl : STD_LOGIC;
  SIGNAL mux_3872_nl : STD_LOGIC;
  SIGNAL or_3502_nl : STD_LOGIC;
  SIGNAL mux_3871_nl : STD_LOGIC;
  SIGNAL mux_3870_nl : STD_LOGIC;
  SIGNAL mux_3869_nl : STD_LOGIC;
  SIGNAL mux_3868_nl : STD_LOGIC;
  SIGNAL mux_3867_nl : STD_LOGIC;
  SIGNAL mux_3866_nl : STD_LOGIC;
  SIGNAL mux_3865_nl : STD_LOGIC;
  SIGNAL mux_3864_nl : STD_LOGIC;
  SIGNAL mux_3863_nl : STD_LOGIC;
  SIGNAL mux_3861_nl : STD_LOGIC;
  SIGNAL or_3500_nl : STD_LOGIC;
  SIGNAL mux_3860_nl : STD_LOGIC;
  SIGNAL mux_3859_nl : STD_LOGIC;
  SIGNAL mux_3858_nl : STD_LOGIC;
  SIGNAL mux_3857_nl : STD_LOGIC;
  SIGNAL mux_3856_nl : STD_LOGIC;
  SIGNAL and_1255_nl : STD_LOGIC;
  SIGNAL mux_3855_nl : STD_LOGIC;
  SIGNAL mux_3853_nl : STD_LOGIC;
  SIGNAL mux_3852_nl : STD_LOGIC;
  SIGNAL mux_3851_nl : STD_LOGIC;
  SIGNAL nor_1456_nl : STD_LOGIC;
  SIGNAL mux_3850_nl : STD_LOGIC;
  SIGNAL mux_3849_nl : STD_LOGIC;
  SIGNAL mux_3848_nl : STD_LOGIC;
  SIGNAL and_1264_nl : STD_LOGIC;
  SIGNAL mux_3846_nl : STD_LOGIC;
  SIGNAL mux_3845_nl : STD_LOGIC;
  SIGNAL mux_3844_nl : STD_LOGIC;
  SIGNAL mux_3843_nl : STD_LOGIC;
  SIGNAL mux_3842_nl : STD_LOGIC;
  SIGNAL or_3493_nl : STD_LOGIC;
  SIGNAL mux_3841_nl : STD_LOGIC;
  SIGNAL nor_1457_nl : STD_LOGIC;
  SIGNAL mux_3840_nl : STD_LOGIC;
  SIGNAL or_3490_nl : STD_LOGIC;
  SIGNAL mux_3839_nl : STD_LOGIC;
  SIGNAL mux_3838_nl : STD_LOGIC;
  SIGNAL mux_3837_nl : STD_LOGIC;
  SIGNAL mux_3836_nl : STD_LOGIC;
  SIGNAL mux_3834_nl : STD_LOGIC;
  SIGNAL mux_3833_nl : STD_LOGIC;
  SIGNAL nor_1458_nl : STD_LOGIC;
  SIGNAL mux_3832_nl : STD_LOGIC;
  SIGNAL mux_3831_nl : STD_LOGIC;
  SIGNAL mux_3830_nl : STD_LOGIC;
  SIGNAL mux_3828_nl : STD_LOGIC;
  SIGNAL mux_3827_nl : STD_LOGIC;
  SIGNAL mux_3826_nl : STD_LOGIC;
  SIGNAL nor_1459_nl : STD_LOGIC;
  SIGNAL mux_3825_nl : STD_LOGIC;
  SIGNAL mux_3824_nl : STD_LOGIC;
  SIGNAL mux_3822_nl : STD_LOGIC;
  SIGNAL or_3480_nl : STD_LOGIC;
  SIGNAL mux_3821_nl : STD_LOGIC;
  SIGNAL mux_3949_nl : STD_LOGIC;
  SIGNAL mux_3948_nl : STD_LOGIC;
  SIGNAL mux_3947_nl : STD_LOGIC;
  SIGNAL mux_3946_nl : STD_LOGIC;
  SIGNAL mux_3945_nl : STD_LOGIC;
  SIGNAL or_3579_nl : STD_LOGIC;
  SIGNAL mux_3944_nl : STD_LOGIC;
  SIGNAL nand_463_nl : STD_LOGIC;
  SIGNAL mux_3943_nl : STD_LOGIC;
  SIGNAL mux_3942_nl : STD_LOGIC;
  SIGNAL or_3577_nl : STD_LOGIC;
  SIGNAL mux_3941_nl : STD_LOGIC;
  SIGNAL mux_3940_nl : STD_LOGIC;
  SIGNAL mux_3939_nl : STD_LOGIC;
  SIGNAL nand_462_nl : STD_LOGIC;
  SIGNAL mux_3938_nl : STD_LOGIC;
  SIGNAL nor_1448_nl : STD_LOGIC;
  SIGNAL nor_1449_nl : STD_LOGIC;
  SIGNAL or_3574_nl : STD_LOGIC;
  SIGNAL or_3572_nl : STD_LOGIC;
  SIGNAL mux_3937_nl : STD_LOGIC;
  SIGNAL mux_3936_nl : STD_LOGIC;
  SIGNAL mux_3935_nl : STD_LOGIC;
  SIGNAL or_3568_nl : STD_LOGIC;
  SIGNAL mux_3934_nl : STD_LOGIC;
  SIGNAL or_3567_nl : STD_LOGIC;
  SIGNAL or_3565_nl : STD_LOGIC;
  SIGNAL mux_3933_nl : STD_LOGIC;
  SIGNAL mux_3932_nl : STD_LOGIC;
  SIGNAL nand_461_nl : STD_LOGIC;
  SIGNAL mux_3931_nl : STD_LOGIC;
  SIGNAL or_3559_nl : STD_LOGIC;
  SIGNAL mux_3930_nl : STD_LOGIC;
  SIGNAL nand_465_nl : STD_LOGIC;
  SIGNAL mux_3929_nl : STD_LOGIC;
  SIGNAL or_3556_nl : STD_LOGIC;
  SIGNAL mux_3928_nl : STD_LOGIC;
  SIGNAL mux_3927_nl : STD_LOGIC;
  SIGNAL mux_3926_nl : STD_LOGIC;
  SIGNAL mux_3925_nl : STD_LOGIC;
  SIGNAL mux_3924_nl : STD_LOGIC;
  SIGNAL mux_3923_nl : STD_LOGIC;
  SIGNAL mux_3922_nl : STD_LOGIC;
  SIGNAL or_3554_nl : STD_LOGIC;
  SIGNAL nand_471_nl : STD_LOGIC;
  SIGNAL mux_3921_nl : STD_LOGIC;
  SIGNAL or_3551_nl : STD_LOGIC;
  SIGNAL or_3550_nl : STD_LOGIC;
  SIGNAL mux_3920_nl : STD_LOGIC;
  SIGNAL mux_3919_nl : STD_LOGIC;
  SIGNAL nand_460_nl : STD_LOGIC;
  SIGNAL mux_3918_nl : STD_LOGIC;
  SIGNAL mux_3917_nl : STD_LOGIC;
  SIGNAL or_3548_nl : STD_LOGIC;
  SIGNAL or_3547_nl : STD_LOGIC;
  SIGNAL mux_3915_nl : STD_LOGIC;
  SIGNAL or_3546_nl : STD_LOGIC;
  SIGNAL mux_3914_nl : STD_LOGIC;
  SIGNAL or_3544_nl : STD_LOGIC;
  SIGNAL mux_3913_nl : STD_LOGIC;
  SIGNAL mux_3912_nl : STD_LOGIC;
  SIGNAL or_3542_nl : STD_LOGIC;
  SIGNAL or_3540_nl : STD_LOGIC;
  SIGNAL nand_459_nl : STD_LOGIC;
  SIGNAL mux_3911_nl : STD_LOGIC;
  SIGNAL or_3536_nl : STD_LOGIC;
  SIGNAL mux_3910_nl : STD_LOGIC;
  SIGNAL or_3534_nl : STD_LOGIC;
  SIGNAL mux_3909_nl : STD_LOGIC;
  SIGNAL or_3533_nl : STD_LOGIC;
  SIGNAL or_3532_nl : STD_LOGIC;
  SIGNAL mux_3908_nl : STD_LOGIC;
  SIGNAL or_3527_nl : STD_LOGIC;
  SIGNAL mux_3905_nl : STD_LOGIC;
  SIGNAL mux_3904_nl : STD_LOGIC;
  SIGNAL or_3589_nl : STD_LOGIC;
  SIGNAL mux_3901_nl : STD_LOGIC;
  SIGNAL mux_3900_nl : STD_LOGIC;
  SIGNAL or_3521_nl : STD_LOGIC;
  SIGNAL mux_3897_nl : STD_LOGIC;
  SIGNAL or_3514_nl : STD_LOGIC;
  SIGNAL or_3477_nl : STD_LOGIC;
  SIGNAL mux_2649_nl : STD_LOGIC;
  SIGNAL mux_2648_nl : STD_LOGIC;
  SIGNAL or_2515_nl : STD_LOGIC;
  SIGNAL or_2514_nl : STD_LOGIC;
  SIGNAL or_2513_nl : STD_LOGIC;
  SIGNAL mux_3952_nl : STD_LOGIC;
  SIGNAL or_3587_nl : STD_LOGIC;
  SIGNAL mux_3951_nl : STD_LOGIC;
  SIGNAL or_3585_nl : STD_LOGIC;
  SIGNAL mux_3950_nl : STD_LOGIC;
  SIGNAL or_3584_nl : STD_LOGIC;
  SIGNAL or_3583_nl : STD_LOGIC;
  SIGNAL or_3581_nl : STD_LOGIC;
  SIGNAL or_3588_nl : STD_LOGIC;
  SIGNAL mux_2675_nl : STD_LOGIC;
  SIGNAL mux_2674_nl : STD_LOGIC;
  SIGNAL mux_2673_nl : STD_LOGIC;
  SIGNAL mux_2672_nl : STD_LOGIC;
  SIGNAL mux_2671_nl : STD_LOGIC;
  SIGNAL mux_2670_nl : STD_LOGIC;
  SIGNAL nor_725_nl : STD_LOGIC;
  SIGNAL mux_2669_nl : STD_LOGIC;
  SIGNAL mux_2668_nl : STD_LOGIC;
  SIGNAL mux_2667_nl : STD_LOGIC;
  SIGNAL nand_244_nl : STD_LOGIC;
  SIGNAL or_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_23_nl : STD_LOGIC;
  SIGNAL mux_2740_nl : STD_LOGIC;
  SIGNAL mux_2739_nl : STD_LOGIC;
  SIGNAL mux_2738_nl : STD_LOGIC;
  SIGNAL mux_2737_nl : STD_LOGIC;
  SIGNAL mux_2736_nl : STD_LOGIC;
  SIGNAL nor_716_nl : STD_LOGIC;
  SIGNAL mux_2735_nl : STD_LOGIC;
  SIGNAL mux_2734_nl : STD_LOGIC;
  SIGNAL mux_2733_nl : STD_LOGIC;
  SIGNAL mux_2732_nl : STD_LOGIC;
  SIGNAL or_3268_nl : STD_LOGIC;
  SIGNAL mux_2731_nl : STD_LOGIC;
  SIGNAL mux_2730_nl : STD_LOGIC;
  SIGNAL mux_2729_nl : STD_LOGIC;
  SIGNAL mux_2728_nl : STD_LOGIC;
  SIGNAL mux_2727_nl : STD_LOGIC;
  SIGNAL mux_55_nl : STD_LOGIC;
  SIGNAL mux_2725_nl : STD_LOGIC;
  SIGNAL mux_2724_nl : STD_LOGIC;
  SIGNAL mux_2723_nl : STD_LOGIC;
  SIGNAL mux_2722_nl : STD_LOGIC;
  SIGNAL mux_50_nl : STD_LOGIC;
  SIGNAL mux_2720_nl : STD_LOGIC;
  SIGNAL mux_2719_nl : STD_LOGIC;
  SIGNAL mux_2718_nl : STD_LOGIC;
  SIGNAL mux_2717_nl : STD_LOGIC;
  SIGNAL mux_2716_nl : STD_LOGIC;
  SIGNAL mux_2715_nl : STD_LOGIC;
  SIGNAL mux_2714_nl : STD_LOGIC;
  SIGNAL mux_2713_nl : STD_LOGIC;
  SIGNAL mux_2712_nl : STD_LOGIC;
  SIGNAL nand_118_nl : STD_LOGIC;
  SIGNAL mux_2711_nl : STD_LOGIC;
  SIGNAL or_3269_nl : STD_LOGIC;
  SIGNAL mux_2710_nl : STD_LOGIC;
  SIGNAL mux_2709_nl : STD_LOGIC;
  SIGNAL mux_2708_nl : STD_LOGIC;
  SIGNAL or_2540_nl : STD_LOGIC;
  SIGNAL mux_2707_nl : STD_LOGIC;
  SIGNAL mux_2706_nl : STD_LOGIC;
  SIGNAL mux_2705_nl : STD_LOGIC;
  SIGNAL mux_2704_nl : STD_LOGIC;
  SIGNAL mux_2703_nl : STD_LOGIC;
  SIGNAL mux_2702_nl : STD_LOGIC;
  SIGNAL mux_29_nl : STD_LOGIC;
  SIGNAL mux_2699_nl : STD_LOGIC;
  SIGNAL mux_2697_nl : STD_LOGIC;
  SIGNAL mux_22_nl : STD_LOGIC;
  SIGNAL or_25_nl : STD_LOGIC;
  SIGNAL or_24_nl : STD_LOGIC;
  SIGNAL mux_2694_nl : STD_LOGIC;
  SIGNAL mux_2693_nl : STD_LOGIC;
  SIGNAL mux_2692_nl : STD_LOGIC;
  SIGNAL mux_2691_nl : STD_LOGIC;
  SIGNAL nand_116_nl : STD_LOGIC;
  SIGNAL mux_17_nl : STD_LOGIC;
  SIGNAL mux_2689_nl : STD_LOGIC;
  SIGNAL mux_2688_nl : STD_LOGIC;
  SIGNAL mux_13_nl : STD_LOGIC;
  SIGNAL or_18_nl : STD_LOGIC;
  SIGNAL mux_2685_nl : STD_LOGIC;
  SIGNAL mux_11_nl : STD_LOGIC;
  SIGNAL mux_10_nl : STD_LOGIC;
  SIGNAL mux_8_nl : STD_LOGIC;
  SIGNAL mux_2679_nl : STD_LOGIC;
  SIGNAL mux_2678_nl : STD_LOGIC;
  SIGNAL mux_2677_nl : STD_LOGIC;
  SIGNAL mux_2769_nl : STD_LOGIC;
  SIGNAL nor_694_nl : STD_LOGIC;
  SIGNAL mux_2768_nl : STD_LOGIC;
  SIGNAL or_2591_nl : STD_LOGIC;
  SIGNAL or_2589_nl : STD_LOGIC;
  SIGNAL mux_2767_nl : STD_LOGIC;
  SIGNAL or_2588_nl : STD_LOGIC;
  SIGNAL and_513_nl : STD_LOGIC;
  SIGNAL mux_2766_nl : STD_LOGIC;
  SIGNAL nor_695_nl : STD_LOGIC;
  SIGNAL nor_696_nl : STD_LOGIC;
  SIGNAL mux_2764_nl : STD_LOGIC;
  SIGNAL and_514_nl : STD_LOGIC;
  SIGNAL mux_2763_nl : STD_LOGIC;
  SIGNAL nor_697_nl : STD_LOGIC;
  SIGNAL nor_698_nl : STD_LOGIC;
  SIGNAL mux_2762_nl : STD_LOGIC;
  SIGNAL or_2581_nl : STD_LOGIC;
  SIGNAL or_2579_nl : STD_LOGIC;
  SIGNAL mux_2761_nl : STD_LOGIC;
  SIGNAL mux_2760_nl : STD_LOGIC;
  SIGNAL mux_2759_nl : STD_LOGIC;
  SIGNAL and_515_nl : STD_LOGIC;
  SIGNAL nor_699_nl : STD_LOGIC;
  SIGNAL nor_700_nl : STD_LOGIC;
  SIGNAL nor_701_nl : STD_LOGIC;
  SIGNAL nor_1302_nl : STD_LOGIC;
  SIGNAL and_801_nl : STD_LOGIC;
  SIGNAL mux_2742_nl : STD_LOGIC;
  SIGNAL nor_715_nl : STD_LOGIC;
  SIGNAL and_340_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_30_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_31_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_277_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_932_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_934_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_936_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_930_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_11_nl : STD_LOGIC;
  SIGNAL mux_114_nl : STD_LOGIC;
  SIGNAL mux_113_nl : STD_LOGIC;
  SIGNAL mux_112_nl : STD_LOGIC;
  SIGNAL nor_1265_nl : STD_LOGIC;
  SIGNAL nor_1266_nl : STD_LOGIC;
  SIGNAL mux_111_nl : STD_LOGIC;
  SIGNAL nor_1267_nl : STD_LOGIC;
  SIGNAL mux_110_nl : STD_LOGIC;
  SIGNAL or_113_nl : STD_LOGIC;
  SIGNAL nand_395_nl : STD_LOGIC;
  SIGNAL mux_109_nl : STD_LOGIC;
  SIGNAL nor_1268_nl : STD_LOGIC;
  SIGNAL mux_108_nl : STD_LOGIC;
  SIGNAL nor_1269_nl : STD_LOGIC;
  SIGNAL mux_107_nl : STD_LOGIC;
  SIGNAL or_109_nl : STD_LOGIC;
  SIGNAL or_108_nl : STD_LOGIC;
  SIGNAL nor_1270_nl : STD_LOGIC;
  SIGNAL mux_106_nl : STD_LOGIC;
  SIGNAL mux_105_nl : STD_LOGIC;
  SIGNAL mux_104_nl : STD_LOGIC;
  SIGNAL nor_1271_nl : STD_LOGIC;
  SIGNAL nor_1272_nl : STD_LOGIC;
  SIGNAL mux_103_nl : STD_LOGIC;
  SIGNAL and_794_nl : STD_LOGIC;
  SIGNAL mux_102_nl : STD_LOGIC;
  SIGNAL and_795_nl : STD_LOGIC;
  SIGNAL nor_1273_nl : STD_LOGIC;
  SIGNAL nor_1274_nl : STD_LOGIC;
  SIGNAL nor_1275_nl : STD_LOGIC;
  SIGNAL mux_101_nl : STD_LOGIC;
  SIGNAL or_98_nl : STD_LOGIC;
  SIGNAL or_96_nl : STD_LOGIC;
  SIGNAL mux_100_nl : STD_LOGIC;
  SIGNAL or_95_nl : STD_LOGIC;
  SIGNAL or_93_nl : STD_LOGIC;
  SIGNAL mux_2867_nl : STD_LOGIC;
  SIGNAL mux_2866_nl : STD_LOGIC;
  SIGNAL mux_2865_nl : STD_LOGIC;
  SIGNAL mux_2864_nl : STD_LOGIC;
  SIGNAL mux_2863_nl : STD_LOGIC;
  SIGNAL mux_2862_nl : STD_LOGIC;
  SIGNAL nor_1303_nl : STD_LOGIC;
  SIGNAL mux_2861_nl : STD_LOGIC;
  SIGNAL mux_2860_nl : STD_LOGIC;
  SIGNAL mux_2859_nl : STD_LOGIC;
  SIGNAL and_506_nl : STD_LOGIC;
  SIGNAL mux_2858_nl : STD_LOGIC;
  SIGNAL and_508_nl : STD_LOGIC;
  SIGNAL mux_2857_nl : STD_LOGIC;
  SIGNAL mux_2856_nl : STD_LOGIC;
  SIGNAL or_2643_nl : STD_LOGIC;
  SIGNAL mux_2855_nl : STD_LOGIC;
  SIGNAL mux_2854_nl : STD_LOGIC;
  SIGNAL mux_2853_nl : STD_LOGIC;
  SIGNAL mux_2852_nl : STD_LOGIC;
  SIGNAL mux_2851_nl : STD_LOGIC;
  SIGNAL mux_2850_nl : STD_LOGIC;
  SIGNAL mux_2849_nl : STD_LOGIC;
  SIGNAL and_346_nl : STD_LOGIC;
  SIGNAL mux_2848_nl : STD_LOGIC;
  SIGNAL mux_2847_nl : STD_LOGIC;
  SIGNAL mux_2846_nl : STD_LOGIC;
  SIGNAL mux_2845_nl : STD_LOGIC;
  SIGNAL mux_2844_nl : STD_LOGIC;
  SIGNAL mux_2843_nl : STD_LOGIC;
  SIGNAL mux_2842_nl : STD_LOGIC;
  SIGNAL mux_2841_nl : STD_LOGIC;
  SIGNAL mux_2840_nl : STD_LOGIC;
  SIGNAL mux_2839_nl : STD_LOGIC;
  SIGNAL or_2639_nl : STD_LOGIC;
  SIGNAL or_2638_nl : STD_LOGIC;
  SIGNAL mux_2838_nl : STD_LOGIC;
  SIGNAL mux_2837_nl : STD_LOGIC;
  SIGNAL or_2637_nl : STD_LOGIC;
  SIGNAL mux_2836_nl : STD_LOGIC;
  SIGNAL mux_2835_nl : STD_LOGIC;
  SIGNAL or_2636_nl : STD_LOGIC;
  SIGNAL mux_2834_nl : STD_LOGIC;
  SIGNAL mux_2833_nl : STD_LOGIC;
  SIGNAL mux_2832_nl : STD_LOGIC;
  SIGNAL or_3347_nl : STD_LOGIC;
  SIGNAL mux_2831_nl : STD_LOGIC;
  SIGNAL mux_2830_nl : STD_LOGIC;
  SIGNAL mux_2829_nl : STD_LOGIC;
  SIGNAL mux_2828_nl : STD_LOGIC;
  SIGNAL or_2632_nl : STD_LOGIC;
  SIGNAL mux_2827_nl : STD_LOGIC;
  SIGNAL mux_2826_nl : STD_LOGIC;
  SIGNAL mux_2825_nl : STD_LOGIC;
  SIGNAL mux_2824_nl : STD_LOGIC;
  SIGNAL mux_2823_nl : STD_LOGIC;
  SIGNAL mux_2822_nl : STD_LOGIC;
  SIGNAL mux_2821_nl : STD_LOGIC;
  SIGNAL mux_2820_nl : STD_LOGIC;
  SIGNAL mux_2819_nl : STD_LOGIC;
  SIGNAL mux_2818_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL mux_2817_nl : STD_LOGIC;
  SIGNAL mux_2816_nl : STD_LOGIC;
  SIGNAL mux_2815_nl : STD_LOGIC;
  SIGNAL mux_2814_nl : STD_LOGIC;
  SIGNAL mux_2812_nl : STD_LOGIC;
  SIGNAL mux_2811_nl : STD_LOGIC;
  SIGNAL mux_2810_nl : STD_LOGIC;
  SIGNAL mux_2809_nl : STD_LOGIC;
  SIGNAL or_2629_nl : STD_LOGIC;
  SIGNAL mux_2808_nl : STD_LOGIC;
  SIGNAL nand_128_nl : STD_LOGIC;
  SIGNAL mux_2807_nl : STD_LOGIC;
  SIGNAL mux_2806_nl : STD_LOGIC;
  SIGNAL mux_2805_nl : STD_LOGIC;
  SIGNAL mux_2804_nl : STD_LOGIC;
  SIGNAL mux_2803_nl : STD_LOGIC;
  SIGNAL mux_2802_nl : STD_LOGIC;
  SIGNAL mux_2801_nl : STD_LOGIC;
  SIGNAL nand_127_nl : STD_LOGIC;
  SIGNAL or_2626_nl : STD_LOGIC;
  SIGNAL mux_2798_nl : STD_LOGIC;
  SIGNAL or_2625_nl : STD_LOGIC;
  SIGNAL or_2624_nl : STD_LOGIC;
  SIGNAL mux_2797_nl : STD_LOGIC;
  SIGNAL or_2622_nl : STD_LOGIC;
  SIGNAL mux_2795_nl : STD_LOGIC;
  SIGNAL mux_2794_nl : STD_LOGIC;
  SIGNAL or_2620_nl : STD_LOGIC;
  SIGNAL mux_2793_nl : STD_LOGIC;
  SIGNAL mux_2792_nl : STD_LOGIC;
  SIGNAL mux_2791_nl : STD_LOGIC;
  SIGNAL mux_2789_nl : STD_LOGIC;
  SIGNAL nand_126_nl : STD_LOGIC;
  SIGNAL mux_2787_nl : STD_LOGIC;
  SIGNAL mux_2786_nl : STD_LOGIC;
  SIGNAL or_199_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_428_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_274_nl : STD_LOGIC;
  SIGNAL mux_2976_nl : STD_LOGIC;
  SIGNAL mux_2975_nl : STD_LOGIC;
  SIGNAL mux_2974_nl : STD_LOGIC;
  SIGNAL mux_2973_nl : STD_LOGIC;
  SIGNAL mux_2972_nl : STD_LOGIC;
  SIGNAL mux_2971_nl : STD_LOGIC;
  SIGNAL or_2728_nl : STD_LOGIC;
  SIGNAL mux_2970_nl : STD_LOGIC;
  SIGNAL mux_2969_nl : STD_LOGIC;
  SIGNAL mux_2968_nl : STD_LOGIC;
  SIGNAL mux_2967_nl : STD_LOGIC;
  SIGNAL mux_2966_nl : STD_LOGIC;
  SIGNAL mux_2965_nl : STD_LOGIC;
  SIGNAL mux_2964_nl : STD_LOGIC;
  SIGNAL mux_2963_nl : STD_LOGIC;
  SIGNAL mux_2962_nl : STD_LOGIC;
  SIGNAL mux_2961_nl : STD_LOGIC;
  SIGNAL mux_2960_nl : STD_LOGIC;
  SIGNAL mux_427_nl : STD_LOGIC;
  SIGNAL mux_426_nl : STD_LOGIC;
  SIGNAL mux_2957_nl : STD_LOGIC;
  SIGNAL mux_2956_nl : STD_LOGIC;
  SIGNAL mux_2955_nl : STD_LOGIC;
  SIGNAL mux_2954_nl : STD_LOGIC;
  SIGNAL mux_422_nl : STD_LOGIC;
  SIGNAL mux_421_nl : STD_LOGIC;
  SIGNAL mux_2951_nl : STD_LOGIC;
  SIGNAL mux_2950_nl : STD_LOGIC;
  SIGNAL mux_2949_nl : STD_LOGIC;
  SIGNAL mux_2948_nl : STD_LOGIC;
  SIGNAL mux_2947_nl : STD_LOGIC;
  SIGNAL mux_2946_nl : STD_LOGIC;
  SIGNAL mux_414_nl : STD_LOGIC;
  SIGNAL mux_2942_nl : STD_LOGIC;
  SIGNAL mux_2941_nl : STD_LOGIC;
  SIGNAL mux_2940_nl : STD_LOGIC;
  SIGNAL mux_2939_nl : STD_LOGIC;
  SIGNAL mux_2938_nl : STD_LOGIC;
  SIGNAL mux_2936_nl : STD_LOGIC;
  SIGNAL mux_2935_nl : STD_LOGIC;
  SIGNAL mux_2934_nl : STD_LOGIC;
  SIGNAL mux_2933_nl : STD_LOGIC;
  SIGNAL mux_2932_nl : STD_LOGIC;
  SIGNAL mux_2931_nl : STD_LOGIC;
  SIGNAL mux_2929_nl : STD_LOGIC;
  SIGNAL mux_2928_nl : STD_LOGIC;
  SIGNAL mux_2927_nl : STD_LOGIC;
  SIGNAL mux_2926_nl : STD_LOGIC;
  SIGNAL mux_2925_nl : STD_LOGIC;
  SIGNAL mux_2924_nl : STD_LOGIC;
  SIGNAL or_2718_nl : STD_LOGIC;
  SIGNAL mux_2923_nl : STD_LOGIC;
  SIGNAL mux_2922_nl : STD_LOGIC;
  SIGNAL mux_2918_nl : STD_LOGIC;
  SIGNAL mux_386_nl : STD_LOGIC;
  SIGNAL mux_2916_nl : STD_LOGIC;
  SIGNAL mux_2914_nl : STD_LOGIC;
  SIGNAL mux_2909_nl : STD_LOGIC;
  SIGNAL mux_2908_nl : STD_LOGIC;
  SIGNAL mux_2888_nl : STD_LOGIC;
  SIGNAL mux_2887_nl : STD_LOGIC;
  SIGNAL or_3351_nl : STD_LOGIC;
  SIGNAL nand_421_nl : STD_LOGIC;
  SIGNAL mux_2886_nl : STD_LOGIC;
  SIGNAL nor_667_nl : STD_LOGIC;
  SIGNAL mux_2885_nl : STD_LOGIC;
  SIGNAL or_2678_nl : STD_LOGIC;
  SIGNAL nor_668_nl : STD_LOGIC;
  SIGNAL mux_2884_nl : STD_LOGIC;
  SIGNAL or_3352_nl : STD_LOGIC;
  SIGNAL mux_2883_nl : STD_LOGIC;
  SIGNAL or_2674_nl : STD_LOGIC;
  SIGNAL or_2673_nl : STD_LOGIC;
  SIGNAL nand_422_nl : STD_LOGIC;
  SIGNAL mux_2882_nl : STD_LOGIC;
  SIGNAL nor_671_nl : STD_LOGIC;
  SIGNAL mux_2983_nl : STD_LOGIC;
  SIGNAL mux_2982_nl : STD_LOGIC;
  SIGNAL mux_2981_nl : STD_LOGIC;
  SIGNAL mux_2980_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL nor_647_nl : STD_LOGIC;
  SIGNAL nor_648_nl : STD_LOGIC;
  SIGNAL nor_649_nl : STD_LOGIC;
  SIGNAL mux_2979_nl : STD_LOGIC;
  SIGNAL nor_650_nl : STD_LOGIC;
  SIGNAL and_490_nl : STD_LOGIC;
  SIGNAL mux_2978_nl : STD_LOGIC;
  SIGNAL mux_2977_nl : STD_LOGIC;
  SIGNAL nor_651_nl : STD_LOGIC;
  SIGNAL nor_652_nl : STD_LOGIC;
  SIGNAL nor_653_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_8_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_3181_nl : STD_LOGIC;
  SIGNAL mux_3180_nl : STD_LOGIC;
  SIGNAL nor_620_nl : STD_LOGIC;
  SIGNAL mux_3179_nl : STD_LOGIC;
  SIGNAL mux_3178_nl : STD_LOGIC;
  SIGNAL or_2838_nl : STD_LOGIC;
  SIGNAL mux_3177_nl : STD_LOGIC;
  SIGNAL nor_621_nl : STD_LOGIC;
  SIGNAL mux_3176_nl : STD_LOGIC;
  SIGNAL mux_3175_nl : STD_LOGIC;
  SIGNAL nor_622_nl : STD_LOGIC;
  SIGNAL nor_623_nl : STD_LOGIC;
  SIGNAL mux_3174_nl : STD_LOGIC;
  SIGNAL mux_3173_nl : STD_LOGIC;
  SIGNAL mux_3172_nl : STD_LOGIC;
  SIGNAL nor_624_nl : STD_LOGIC;
  SIGNAL nor_625_nl : STD_LOGIC;
  SIGNAL mux_3171_nl : STD_LOGIC;
  SIGNAL mux_3170_nl : STD_LOGIC;
  SIGNAL or_2828_nl : STD_LOGIC;
  SIGNAL or_2827_nl : STD_LOGIC;
  SIGNAL and_465_nl : STD_LOGIC;
  SIGNAL mux_3169_nl : STD_LOGIC;
  SIGNAL nor_626_nl : STD_LOGIC;
  SIGNAL mux_3167_nl : STD_LOGIC;
  SIGNAL or_2817_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL nor_nl : STD_LOGIC;
  SIGNAL and_1253_nl : STD_LOGIC;
  SIGNAL mux_3217_nl : STD_LOGIC;
  SIGNAL mux_3216_nl : STD_LOGIC;
  SIGNAL or_3259_nl : STD_LOGIC;
  SIGNAL mux_3215_nl : STD_LOGIC;
  SIGNAL nor_617_nl : STD_LOGIC;
  SIGNAL or_2888_nl : STD_LOGIC;
  SIGNAL mux_3224_nl : STD_LOGIC;
  SIGNAL mux_3223_nl : STD_LOGIC;
  SIGNAL mux_3222_nl : STD_LOGIC;
  SIGNAL mux_3221_nl : STD_LOGIC;
  SIGNAL mux_3220_nl : STD_LOGIC;
  SIGNAL and_452_nl : STD_LOGIC;
  SIGNAL and_454_nl : STD_LOGIC;
  SIGNAL mux_3234_nl : STD_LOGIC;
  SIGNAL mux_3233_nl : STD_LOGIC;
  SIGNAL mux_3232_nl : STD_LOGIC;
  SIGNAL mux_3231_nl : STD_LOGIC;
  SIGNAL mux_3230_nl : STD_LOGIC;
  SIGNAL mux_3229_nl : STD_LOGIC;
  SIGNAL and_363_nl : STD_LOGIC;
  SIGNAL mux_3228_nl : STD_LOGIC;
  SIGNAL mux_3227_nl : STD_LOGIC;
  SIGNAL mux_3226_nl : STD_LOGIC;
  SIGNAL nor_729_nl : STD_LOGIC;
  SIGNAL mux_3225_nl : STD_LOGIC;
  SIGNAL mux_3242_nl : STD_LOGIC;
  SIGNAL mux_3241_nl : STD_LOGIC;
  SIGNAL mux_3240_nl : STD_LOGIC;
  SIGNAL mux_3239_nl : STD_LOGIC;
  SIGNAL mux_3238_nl : STD_LOGIC;
  SIGNAL or_2906_nl : STD_LOGIC;
  SIGNAL mux_3237_nl : STD_LOGIC;
  SIGNAL mux_3243_nl : STD_LOGIC;
  SIGNAL or_3252_nl : STD_LOGIC;
  SIGNAL nand_218_nl : STD_LOGIC;
  SIGNAL mux_3249_nl : STD_LOGIC;
  SIGNAL mux_3248_nl : STD_LOGIC;
  SIGNAL mux_3247_nl : STD_LOGIC;
  SIGNAL mux_3246_nl : STD_LOGIC;
  SIGNAL mux_3245_nl : STD_LOGIC;
  SIGNAL or_2915_nl : STD_LOGIC;
  SIGNAL or_2913_nl : STD_LOGIC;
  SIGNAL mux_3251_nl : STD_LOGIC;
  SIGNAL mux_3250_nl : STD_LOGIC;
  SIGNAL nor_1317_nl : STD_LOGIC;
  SIGNAL or_3346_nl : STD_LOGIC;
  SIGNAL mux_3255_nl : STD_LOGIC;
  SIGNAL mux_3254_nl : STD_LOGIC;
  SIGNAL mux_3253_nl : STD_LOGIC;
  SIGNAL nor_611_nl : STD_LOGIC;
  SIGNAL mux_3252_nl : STD_LOGIC;
  SIGNAL and_371_nl : STD_LOGIC;
  SIGNAL or_2922_nl : STD_LOGIC;
  SIGNAL mux_3263_nl : STD_LOGIC;
  SIGNAL mux_3262_nl : STD_LOGIC;
  SIGNAL mux_3261_nl : STD_LOGIC;
  SIGNAL mux_3260_nl : STD_LOGIC;
  SIGNAL mux_3259_nl : STD_LOGIC;
  SIGNAL mux_3258_nl : STD_LOGIC;
  SIGNAL mux_3257_nl : STD_LOGIC;
  SIGNAL mux_3267_nl : STD_LOGIC;
  SIGNAL mux_3266_nl : STD_LOGIC;
  SIGNAL mux_3265_nl : STD_LOGIC;
  SIGNAL or_2933_nl : STD_LOGIC;
  SIGNAL mux_3264_nl : STD_LOGIC;
  SIGNAL or_2930_nl : STD_LOGIC;
  SIGNAL mux_3276_nl : STD_LOGIC;
  SIGNAL mux_3275_nl : STD_LOGIC;
  SIGNAL mux_3274_nl : STD_LOGIC;
  SIGNAL mux_3273_nl : STD_LOGIC;
  SIGNAL mux_3272_nl : STD_LOGIC;
  SIGNAL mux_3271_nl : STD_LOGIC;
  SIGNAL mux_3270_nl : STD_LOGIC;
  SIGNAL and_439_nl : STD_LOGIC;
  SIGNAL mux_3288_nl : STD_LOGIC;
  SIGNAL mux_3287_nl : STD_LOGIC;
  SIGNAL mux_3286_nl : STD_LOGIC;
  SIGNAL mux_3285_nl : STD_LOGIC;
  SIGNAL and_434_nl : STD_LOGIC;
  SIGNAL mux_3284_nl : STD_LOGIC;
  SIGNAL mux_3283_nl : STD_LOGIC;
  SIGNAL mux_3282_nl : STD_LOGIC;
  SIGNAL mux_3292_nl : STD_LOGIC;
  SIGNAL mux_3291_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL mux_3290_nl : STD_LOGIC;
  SIGNAL nor_605_nl : STD_LOGIC;
  SIGNAL and_431_nl : STD_LOGIC;
  SIGNAL and_433_nl : STD_LOGIC;
  SIGNAL mux_3297_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL mux_3296_nl : STD_LOGIC;
  SIGNAL or_2947_nl : STD_LOGIC;
  SIGNAL and_375_nl : STD_LOGIC;
  SIGNAL mux_3295_nl : STD_LOGIC;
  SIGNAL and_374_nl : STD_LOGIC;
  SIGNAL mux_3294_nl : STD_LOGIC;
  SIGNAL and_430_nl : STD_LOGIC;
  SIGNAL or_2945_nl : STD_LOGIC;
  SIGNAL nor_1420_nl : STD_LOGIC;
  SIGNAL mux_3299_nl : STD_LOGIC;
  SIGNAL or_2950_nl : STD_LOGIC;
  SIGNAL and_1254_nl : STD_LOGIC;
  SIGNAL mux_3304_nl : STD_LOGIC;
  SIGNAL nor_1201_nl : STD_LOGIC;
  SIGNAL mux_3303_nl : STD_LOGIC;
  SIGNAL mux_3302_nl : STD_LOGIC;
  SIGNAL mux_3301_nl : STD_LOGIC;
  SIGNAL and_29_nl : STD_LOGIC;
  SIGNAL mux_3393_nl : STD_LOGIC;
  SIGNAL or_3014_nl : STD_LOGIC;
  SIGNAL mux_3384_nl : STD_LOGIC;
  SIGNAL or_3004_nl : STD_LOGIC;
  SIGNAL or_3001_nl : STD_LOGIC;
  SIGNAL nor_581_nl : STD_LOGIC;
  SIGNAL mux_3391_nl : STD_LOGIC;
  SIGNAL nor_582_nl : STD_LOGIC;
  SIGNAL mux_3390_nl : STD_LOGIC;
  SIGNAL and_414_nl : STD_LOGIC;
  SIGNAL mux_3389_nl : STD_LOGIC;
  SIGNAL nor_583_nl : STD_LOGIC;
  SIGNAL and_415_nl : STD_LOGIC;
  SIGNAL nor_584_nl : STD_LOGIC;
  SIGNAL mux_3387_nl : STD_LOGIC;
  SIGNAL and_416_nl : STD_LOGIC;
  SIGNAL nor_585_nl : STD_LOGIC;
  SIGNAL nor_586_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_464_nl : STD_LOGIC;
  SIGNAL mux_3396_nl : STD_LOGIC;
  SIGNAL mux_3395_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL or_3241_nl : STD_LOGIC;
  SIGNAL nand_205_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_474_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_12_nl : STD_LOGIC;
  SIGNAL mux_3492_nl : STD_LOGIC;
  SIGNAL mux_3491_nl : STD_LOGIC;
  SIGNAL mux_3490_nl : STD_LOGIC;
  SIGNAL mux_3489_nl : STD_LOGIC;
  SIGNAL mux_3488_nl : STD_LOGIC;
  SIGNAL mux_3487_nl : STD_LOGIC;
  SIGNAL mux_3486_nl : STD_LOGIC;
  SIGNAL mux_3485_nl : STD_LOGIC;
  SIGNAL mux_3484_nl : STD_LOGIC;
  SIGNAL mux_3483_nl : STD_LOGIC;
  SIGNAL mux_3482_nl : STD_LOGIC;
  SIGNAL mux_3481_nl : STD_LOGIC;
  SIGNAL mux_3480_nl : STD_LOGIC;
  SIGNAL mux_3479_nl : STD_LOGIC;
  SIGNAL mux_3478_nl : STD_LOGIC;
  SIGNAL mux_3477_nl : STD_LOGIC;
  SIGNAL mux_3476_nl : STD_LOGIC;
  SIGNAL mux_3475_nl : STD_LOGIC;
  SIGNAL mux_3474_nl : STD_LOGIC;
  SIGNAL mux_3473_nl : STD_LOGIC;
  SIGNAL mux_3472_nl : STD_LOGIC;
  SIGNAL mux_3470_nl : STD_LOGIC;
  SIGNAL mux_3469_nl : STD_LOGIC;
  SIGNAL mux_3466_nl : STD_LOGIC;
  SIGNAL mux_3465_nl : STD_LOGIC;
  SIGNAL mux_3464_nl : STD_LOGIC;
  SIGNAL mux_3463_nl : STD_LOGIC;
  SIGNAL mux_3462_nl : STD_LOGIC;
  SIGNAL mux_3461_nl : STD_LOGIC;
  SIGNAL mux_3460_nl : STD_LOGIC;
  SIGNAL mux_3457_nl : STD_LOGIC;
  SIGNAL mux_3455_nl : STD_LOGIC;
  SIGNAL mux_3454_nl : STD_LOGIC;
  SIGNAL mux_3453_nl : STD_LOGIC;
  SIGNAL mux_3451_nl : STD_LOGIC;
  SIGNAL mux_3448_nl : STD_LOGIC;
  SIGNAL mux_3447_nl : STD_LOGIC;
  SIGNAL mux_3446_nl : STD_LOGIC;
  SIGNAL mux_3445_nl : STD_LOGIC;
  SIGNAL mux_3444_nl : STD_LOGIC;
  SIGNAL mux_3443_nl : STD_LOGIC;
  SIGNAL mux_3442_nl : STD_LOGIC;
  SIGNAL mux_3441_nl : STD_LOGIC;
  SIGNAL mux_3440_nl : STD_LOGIC;
  SIGNAL mux_3439_nl : STD_LOGIC;
  SIGNAL mux_3438_nl : STD_LOGIC;
  SIGNAL mux_3437_nl : STD_LOGIC;
  SIGNAL mux_3435_nl : STD_LOGIC;
  SIGNAL mux_3434_nl : STD_LOGIC;
  SIGNAL mux_3433_nl : STD_LOGIC;
  SIGNAL mux_3432_nl : STD_LOGIC;
  SIGNAL mux_3431_nl : STD_LOGIC;
  SIGNAL mux_3429_nl : STD_LOGIC;
  SIGNAL mux_3428_nl : STD_LOGIC;
  SIGNAL mux_3427_nl : STD_LOGIC;
  SIGNAL mux_3425_nl : STD_LOGIC;
  SIGNAL mux_3424_nl : STD_LOGIC;
  SIGNAL mux_3420_nl : STD_LOGIC;
  SIGNAL mux_3506_nl : STD_LOGIC;
  SIGNAL mux_3505_nl : STD_LOGIC;
  SIGNAL or_3090_nl : STD_LOGIC;
  SIGNAL mux_3502_nl : STD_LOGIC;
  SIGNAL or_3084_nl : STD_LOGIC;
  SIGNAL mux_3501_nl : STD_LOGIC;
  SIGNAL or_3083_nl : STD_LOGIC;
  SIGNAL mux_3500_nl : STD_LOGIC;
  SIGNAL mux_3499_nl : STD_LOGIC;
  SIGNAL or_3079_nl : STD_LOGIC;
  SIGNAL mux_3497_nl : STD_LOGIC;
  SIGNAL mux_3496_nl : STD_LOGIC;
  SIGNAL nand_168_nl : STD_LOGIC;
  SIGNAL or_3076_nl : STD_LOGIC;
  SIGNAL or_3071_nl : STD_LOGIC;
  SIGNAL mux_3417_nl : STD_LOGIC;
  SIGNAL nor_569_nl : STD_LOGIC;
  SIGNAL mux_3416_nl : STD_LOGIC;
  SIGNAL or_3055_nl : STD_LOGIC;
  SIGNAL mux_3415_nl : STD_LOGIC;
  SIGNAL or_3054_nl : STD_LOGIC;
  SIGNAL or_3053_nl : STD_LOGIC;
  SIGNAL mux_3414_nl : STD_LOGIC;
  SIGNAL or_3052_nl : STD_LOGIC;
  SIGNAL or_3051_nl : STD_LOGIC;
  SIGNAL and_409_nl : STD_LOGIC;
  SIGNAL mux_3413_nl : STD_LOGIC;
  SIGNAL and_410_nl : STD_LOGIC;
  SIGNAL mux_3412_nl : STD_LOGIC;
  SIGNAL nor_570_nl : STD_LOGIC;
  SIGNAL nor_571_nl : STD_LOGIC;
  SIGNAL nor_572_nl : STD_LOGIC;
  SIGNAL mux_3411_nl : STD_LOGIC;
  SIGNAL or_3044_nl : STD_LOGIC;
  SIGNAL nand_208_nl : STD_LOGIC;
  SIGNAL mux_3513_nl : STD_LOGIC;
  SIGNAL mux_3512_nl : STD_LOGIC;
  SIGNAL mux_3511_nl : STD_LOGIC;
  SIGNAL or_3348_nl : STD_LOGIC;
  SIGNAL or_3349_nl : STD_LOGIC;
  SIGNAL mux_3510_nl : STD_LOGIC;
  SIGNAL or_3099_nl : STD_LOGIC;
  SIGNAL or_3350_nl : STD_LOGIC;
  SIGNAL mux_3509_nl : STD_LOGIC;
  SIGNAL or_3097_nl : STD_LOGIC;
  SIGNAL or_3095_nl : STD_LOGIC;
  SIGNAL nand_420_nl : STD_LOGIC;
  SIGNAL mux_3508_nl : STD_LOGIC;
  SIGNAL nor_567_nl : STD_LOGIC;
  SIGNAL and_402_nl : STD_LOGIC;
  SIGNAL mux_3507_nl : STD_LOGIC;
  SIGNAL or_3091_nl : STD_LOGIC;
  SIGNAL mux_3556_nl : STD_LOGIC;
  SIGNAL mux_3574_nl : STD_LOGIC;
  SIGNAL mux_3573_nl : STD_LOGIC;
  SIGNAL mux_3572_nl : STD_LOGIC;
  SIGNAL or_3120_nl : STD_LOGIC;
  SIGNAL mux_3056_nl : STD_LOGIC;
  SIGNAL mux_3570_nl : STD_LOGIC;
  SIGNAL mux_3569_nl : STD_LOGIC;
  SIGNAL mux_433_nl : STD_LOGIC;
  SIGNAL or_3119_nl : STD_LOGIC;
  SIGNAL mux_3567_nl : STD_LOGIC;
  SIGNAL mux_3566_nl : STD_LOGIC;
  SIGNAL mux_438_nl : STD_LOGIC;
  SIGNAL mux_437_nl : STD_LOGIC;
  SIGNAL mux_431_nl : STD_LOGIC;
  SIGNAL mux_3554_nl : STD_LOGIC;
  SIGNAL mux_420_nl : STD_LOGIC;
  SIGNAL mux_419_nl : STD_LOGIC;
  SIGNAL mux_3550_nl : STD_LOGIC;
  SIGNAL mux_3549_nl : STD_LOGIC;
  SIGNAL mux_3548_nl : STD_LOGIC;
  SIGNAL mux_3547_nl : STD_LOGIC;
  SIGNAL mux_3546_nl : STD_LOGIC;
  SIGNAL mux_403_nl : STD_LOGIC;
  SIGNAL or_3115_nl : STD_LOGIC;
  SIGNAL mux_3544_nl : STD_LOGIC;
  SIGNAL mux_3543_nl : STD_LOGIC;
  SIGNAL mux_3542_nl : STD_LOGIC;
  SIGNAL mux_402_nl : STD_LOGIC;
  SIGNAL mux_401_nl : STD_LOGIC;
  SIGNAL mux_400_nl : STD_LOGIC;
  SIGNAL mux_3536_nl : STD_LOGIC;
  SIGNAL mux_3535_nl : STD_LOGIC;
  SIGNAL mux_3534_nl : STD_LOGIC;
  SIGNAL mux_3533_nl : STD_LOGIC;
  SIGNAL nand_173_nl : STD_LOGIC;
  SIGNAL mux_3532_nl : STD_LOGIC;
  SIGNAL mux_3529_nl : STD_LOGIC;
  SIGNAL mux_3528_nl : STD_LOGIC;
  SIGNAL mux_3527_nl : STD_LOGIC;
  SIGNAL mux_383_nl : STD_LOGIC;
  SIGNAL mux_377_nl : STD_LOGIC;
  SIGNAL mux_376_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_477_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_14_nl : STD_LOGIC;
  SIGNAL mux_3577_nl : STD_LOGIC;
  SIGNAL mux_3576_nl : STD_LOGIC;
  SIGNAL mux_3562_nl : STD_LOGIC;
  SIGNAL mux_3561_nl : STD_LOGIC;
  SIGNAL mux_3560_nl : STD_LOGIC;
  SIGNAL mux_3559_nl : STD_LOGIC;
  SIGNAL mux_3558_nl : STD_LOGIC;
  SIGNAL mux_3584_nl : STD_LOGIC;
  SIGNAL mux_3583_nl : STD_LOGIC;
  SIGNAL nand_452_nl : STD_LOGIC;
  SIGNAL mux_3582_nl : STD_LOGIC;
  SIGNAL nor_558_nl : STD_LOGIC;
  SIGNAL nor_559_nl : STD_LOGIC;
  SIGNAL or_3474_nl : STD_LOGIC;
  SIGNAL mux_3581_nl : STD_LOGIC;
  SIGNAL or_3475_nl : STD_LOGIC;
  SIGNAL mux_3580_nl : STD_LOGIC;
  SIGNAL mux_3579_nl : STD_LOGIC;
  SIGNAL or_3127_nl : STD_LOGIC;
  SIGNAL or_3126_nl : STD_LOGIC;
  SIGNAL or_3125_nl : STD_LOGIC;
  SIGNAL nand_453_nl : STD_LOGIC;
  SIGNAL mux_3578_nl : STD_LOGIC;
  SIGNAL nor_562_nl : STD_LOGIC;
  SIGNAL nor_563_nl : STD_LOGIC;
  SIGNAL mux_3591_nl : STD_LOGIC;
  SIGNAL and_391_nl : STD_LOGIC;
  SIGNAL mux_3590_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL mux_3589_nl : STD_LOGIC;
  SIGNAL or_3145_nl : STD_LOGIC;
  SIGNAL and_392_nl : STD_LOGIC;
  SIGNAL mux_3588_nl : STD_LOGIC;
  SIGNAL nor_554_nl : STD_LOGIC;
  SIGNAL mux_3587_nl : STD_LOGIC;
  SIGNAL mux_3586_nl : STD_LOGIC;
  SIGNAL nor_555_nl : STD_LOGIC;
  SIGNAL nor_556_nl : STD_LOGIC;
  SIGNAL mux_3585_nl : STD_LOGIC;
  SIGNAL or_3136_nl : STD_LOGIC;
  SIGNAL or_3135_nl : STD_LOGIC;
  SIGNAL nor_557_nl : STD_LOGIC;
  SIGNAL nor_540_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_479_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_17_nl : STD_LOGIC;
  SIGNAL mux_3598_nl : STD_LOGIC;
  SIGNAL or_3342_nl : STD_LOGIC;
  SIGNAL mux_3597_nl : STD_LOGIC;
  SIGNAL mux_3596_nl : STD_LOGIC;
  SIGNAL or_3158_nl : STD_LOGIC;
  SIGNAL or_3156_nl : STD_LOGIC;
  SIGNAL or_3155_nl : STD_LOGIC;
  SIGNAL mux_3595_nl : STD_LOGIC;
  SIGNAL mux_3594_nl : STD_LOGIC;
  SIGNAL or_3343_nl : STD_LOGIC;
  SIGNAL nand_419_nl : STD_LOGIC;
  SIGNAL mux_3593_nl : STD_LOGIC;
  SIGNAL nor_548_nl : STD_LOGIC;
  SIGNAL and_820_nl : STD_LOGIC;
  SIGNAL mux_3592_nl : STD_LOGIC;
  SIGNAL or_3344_nl : STD_LOGIC;
  SIGNAL or_3345_nl : STD_LOGIC;
  SIGNAL mux_3605_nl : STD_LOGIC;
  SIGNAL nor_538_nl : STD_LOGIC;
  SIGNAL mux_3604_nl : STD_LOGIC;
  SIGNAL nand_181_nl : STD_LOGIC;
  SIGNAL nand_180_nl : STD_LOGIC;
  SIGNAL mux_3602_nl : STD_LOGIC;
  SIGNAL nor_541_nl : STD_LOGIC;
  SIGNAL nor_542_nl : STD_LOGIC;
  SIGNAL mux_3601_nl : STD_LOGIC;
  SIGNAL and_389_nl : STD_LOGIC;
  SIGNAL mux_3600_nl : STD_LOGIC;
  SIGNAL mux_3599_nl : STD_LOGIC;
  SIGNAL nor_543_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_480_nl : STD_LOGIC;
  SIGNAL mux_3673_nl : STD_LOGIC;
  SIGNAL mux_3672_nl : STD_LOGIC;
  SIGNAL mux_3671_nl : STD_LOGIC;
  SIGNAL mux_3670_nl : STD_LOGIC;
  SIGNAL mux_3669_nl : STD_LOGIC;
  SIGNAL mux_3668_nl : STD_LOGIC;
  SIGNAL mux_3667_nl : STD_LOGIC;
  SIGNAL mux_3666_nl : STD_LOGIC;
  SIGNAL mux_3665_nl : STD_LOGIC;
  SIGNAL nand_195_nl : STD_LOGIC;
  SIGNAL mux_3664_nl : STD_LOGIC;
  SIGNAL and_388_nl : STD_LOGIC;
  SIGNAL mux_3663_nl : STD_LOGIC;
  SIGNAL mux_3662_nl : STD_LOGIC;
  SIGNAL mux_3661_nl : STD_LOGIC;
  SIGNAL mux_3660_nl : STD_LOGIC;
  SIGNAL mux_3659_nl : STD_LOGIC;
  SIGNAL and_386_nl : STD_LOGIC;
  SIGNAL mux_3658_nl : STD_LOGIC;
  SIGNAL mux_3657_nl : STD_LOGIC;
  SIGNAL or_3182_nl : STD_LOGIC;
  SIGNAL and_385_nl : STD_LOGIC;
  SIGNAL mux_3656_nl : STD_LOGIC;
  SIGNAL mux_3655_nl : STD_LOGIC;
  SIGNAL mux_3654_nl : STD_LOGIC;
  SIGNAL mux_3653_nl : STD_LOGIC;
  SIGNAL mux_3652_nl : STD_LOGIC;
  SIGNAL mux_3651_nl : STD_LOGIC;
  SIGNAL mux_3650_nl : STD_LOGIC;
  SIGNAL nand_196_nl : STD_LOGIC;
  SIGNAL mux_3649_nl : STD_LOGIC;
  SIGNAL mux_3648_nl : STD_LOGIC;
  SIGNAL mux_3647_nl : STD_LOGIC;
  SIGNAL mux_3646_nl : STD_LOGIC;
  SIGNAL mux_3645_nl : STD_LOGIC;
  SIGNAL mux_3644_nl : STD_LOGIC;
  SIGNAL mux_3643_nl : STD_LOGIC;
  SIGNAL mux_3642_nl : STD_LOGIC;
  SIGNAL mux_3641_nl : STD_LOGIC;
  SIGNAL mux_3640_nl : STD_LOGIC;
  SIGNAL mux_3639_nl : STD_LOGIC;
  SIGNAL nor_536_nl : STD_LOGIC;
  SIGNAL mux_3638_nl : STD_LOGIC;
  SIGNAL nand_197_nl : STD_LOGIC;
  SIGNAL mux_3637_nl : STD_LOGIC;
  SIGNAL mux_3636_nl : STD_LOGIC;
  SIGNAL mux_3635_nl : STD_LOGIC;
  SIGNAL mux_3634_nl : STD_LOGIC;
  SIGNAL mux_3633_nl : STD_LOGIC;
  SIGNAL mux_3632_nl : STD_LOGIC;
  SIGNAL mux_3631_nl : STD_LOGIC;
  SIGNAL mux_3630_nl : STD_LOGIC;
  SIGNAL mux_3629_nl : STD_LOGIC;
  SIGNAL mux_3627_nl : STD_LOGIC;
  SIGNAL mux_3626_nl : STD_LOGIC;
  SIGNAL mux_3625_nl : STD_LOGIC;
  SIGNAL mux_3624_nl : STD_LOGIC;
  SIGNAL mux_3623_nl : STD_LOGIC;
  SIGNAL mux_2589_nl : STD_LOGIC;
  SIGNAL mux_3622_nl : STD_LOGIC;
  SIGNAL or_3179_nl : STD_LOGIC;
  SIGNAL mux_3621_nl : STD_LOGIC;
  SIGNAL mux_3620_nl : STD_LOGIC;
  SIGNAL mux_3619_nl : STD_LOGIC;
  SIGNAL mux_3618_nl : STD_LOGIC;
  SIGNAL mux_3617_nl : STD_LOGIC;
  SIGNAL or_3178_nl : STD_LOGIC;
  SIGNAL mux_3616_nl : STD_LOGIC;
  SIGNAL or_3176_nl : STD_LOGIC;
  SIGNAL mux_3615_nl : STD_LOGIC;
  SIGNAL mux_3614_nl : STD_LOGIC;
  SIGNAL mux_3612_nl : STD_LOGIC;
  SIGNAL mux_3611_nl : STD_LOGIC;
  SIGNAL mux_3610_nl : STD_LOGIC;
  SIGNAL mux_3609_nl : STD_LOGIC;
  SIGNAL mux_3608_nl : STD_LOGIC;
  SIGNAL mux_3607_nl : STD_LOGIC;
  SIGNAL mux_3606_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_28_nl : STD_LOGIC;
  SIGNAL mux_371_nl : STD_LOGIC;
  SIGNAL mux_372_nl : STD_LOGIC;
  SIGNAL mux_406_nl : STD_LOGIC;
  SIGNAL mux_1027_nl : STD_LOGIC;
  SIGNAL or_3295_nl : STD_LOGIC;
  SIGNAL and_659_nl : STD_LOGIC;
  SIGNAL nor_1193_nl : STD_LOGIC;
  SIGNAL or_579_nl : STD_LOGIC;
  SIGNAL mux_1061_nl : STD_LOGIC;
  SIGNAL or_578_nl : STD_LOGIC;
  SIGNAL or_577_nl : STD_LOGIC;
  SIGNAL mux_1066_nl : STD_LOGIC;
  SIGNAL mux_1065_nl : STD_LOGIC;
  SIGNAL or_587_nl : STD_LOGIC;
  SIGNAL or_586_nl : STD_LOGIC;
  SIGNAL or_585_nl : STD_LOGIC;
  SIGNAL or_583_nl : STD_LOGIC;
  SIGNAL or_591_nl : STD_LOGIC;
  SIGNAL or_589_nl : STD_LOGIC;
  SIGNAL mux_1087_nl : STD_LOGIC;
  SIGNAL or_614_nl : STD_LOGIC;
  SIGNAL or_613_nl : STD_LOGIC;
  SIGNAL mux_1086_nl : STD_LOGIC;
  SIGNAL or_611_nl : STD_LOGIC;
  SIGNAL or_610_nl : STD_LOGIC;
  SIGNAL mux_1080_nl : STD_LOGIC;
  SIGNAL nor_1170_nl : STD_LOGIC;
  SIGNAL nor_1171_nl : STD_LOGIC;
  SIGNAL or_600_nl : STD_LOGIC;
  SIGNAL or_599_nl : STD_LOGIC;
  SIGNAL or_693_nl : STD_LOGIC;
  SIGNAL mux_1138_nl : STD_LOGIC;
  SIGNAL or_692_nl : STD_LOGIC;
  SIGNAL or_691_nl : STD_LOGIC;
  SIGNAL mux_1149_nl : STD_LOGIC;
  SIGNAL mux_1148_nl : STD_LOGIC;
  SIGNAL or_709_nl : STD_LOGIC;
  SIGNAL or_708_nl : STD_LOGIC;
  SIGNAL or_707_nl : STD_LOGIC;
  SIGNAL or_705_nl : STD_LOGIC;
  SIGNAL or_712_nl : STD_LOGIC;
  SIGNAL or_710_nl : STD_LOGIC;
  SIGNAL or_792_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL or_791_nl : STD_LOGIC;
  SIGNAL or_790_nl : STD_LOGIC;
  SIGNAL mux_1210_nl : STD_LOGIC;
  SIGNAL mux_1209_nl : STD_LOGIC;
  SIGNAL or_800_nl : STD_LOGIC;
  SIGNAL or_799_nl : STD_LOGIC;
  SIGNAL or_798_nl : STD_LOGIC;
  SIGNAL or_796_nl : STD_LOGIC;
  SIGNAL or_804_nl : STD_LOGIC;
  SIGNAL or_802_nl : STD_LOGIC;
  SIGNAL or_906_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL or_905_nl : STD_LOGIC;
  SIGNAL or_904_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL mux_1292_nl : STD_LOGIC;
  SIGNAL or_922_nl : STD_LOGIC;
  SIGNAL or_921_nl : STD_LOGIC;
  SIGNAL nand_433_nl : STD_LOGIC;
  SIGNAL or_918_nl : STD_LOGIC;
  SIGNAL or_925_nl : STD_LOGIC;
  SIGNAL or_923_nl : STD_LOGIC;
  SIGNAL or_1005_nl : STD_LOGIC;
  SIGNAL mux_1349_nl : STD_LOGIC;
  SIGNAL or_1004_nl : STD_LOGIC;
  SIGNAL or_1003_nl : STD_LOGIC;
  SIGNAL mux_1354_nl : STD_LOGIC;
  SIGNAL mux_1353_nl : STD_LOGIC;
  SIGNAL or_1013_nl : STD_LOGIC;
  SIGNAL or_1012_nl : STD_LOGIC;
  SIGNAL or_1011_nl : STD_LOGIC;
  SIGNAL or_1009_nl : STD_LOGIC;
  SIGNAL or_1017_nl : STD_LOGIC;
  SIGNAL or_1015_nl : STD_LOGIC;
  SIGNAL or_1119_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL or_1118_nl : STD_LOGIC;
  SIGNAL or_1117_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL mux_1436_nl : STD_LOGIC;
  SIGNAL or_1135_nl : STD_LOGIC;
  SIGNAL or_1134_nl : STD_LOGIC;
  SIGNAL nand_432_nl : STD_LOGIC;
  SIGNAL or_1131_nl : STD_LOGIC;
  SIGNAL or_1138_nl : STD_LOGIC;
  SIGNAL or_1136_nl : STD_LOGIC;
  SIGNAL or_1218_nl : STD_LOGIC;
  SIGNAL mux_1493_nl : STD_LOGIC;
  SIGNAL or_1217_nl : STD_LOGIC;
  SIGNAL or_1216_nl : STD_LOGIC;
  SIGNAL mux_1498_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL or_1226_nl : STD_LOGIC;
  SIGNAL or_1225_nl : STD_LOGIC;
  SIGNAL nand_431_nl : STD_LOGIC;
  SIGNAL or_1222_nl : STD_LOGIC;
  SIGNAL or_1230_nl : STD_LOGIC;
  SIGNAL or_1228_nl : STD_LOGIC;
  SIGNAL or_1332_nl : STD_LOGIC;
  SIGNAL mux_1570_nl : STD_LOGIC;
  SIGNAL or_1331_nl : STD_LOGIC;
  SIGNAL or_1330_nl : STD_LOGIC;
  SIGNAL mux_1581_nl : STD_LOGIC;
  SIGNAL mux_1580_nl : STD_LOGIC;
  SIGNAL or_1348_nl : STD_LOGIC;
  SIGNAL or_1347_nl : STD_LOGIC;
  SIGNAL nand_430_nl : STD_LOGIC;
  SIGNAL or_1344_nl : STD_LOGIC;
  SIGNAL nand_418_nl : STD_LOGIC;
  SIGNAL or_1349_nl : STD_LOGIC;
  SIGNAL or_1431_nl : STD_LOGIC;
  SIGNAL mux_1637_nl : STD_LOGIC;
  SIGNAL or_1430_nl : STD_LOGIC;
  SIGNAL or_1429_nl : STD_LOGIC;
  SIGNAL mux_1642_nl : STD_LOGIC;
  SIGNAL mux_1641_nl : STD_LOGIC;
  SIGNAL or_1439_nl : STD_LOGIC;
  SIGNAL or_1438_nl : STD_LOGIC;
  SIGNAL or_1437_nl : STD_LOGIC;
  SIGNAL or_1435_nl : STD_LOGIC;
  SIGNAL or_1443_nl : STD_LOGIC;
  SIGNAL or_1441_nl : STD_LOGIC;
  SIGNAL or_1545_nl : STD_LOGIC;
  SIGNAL mux_1714_nl : STD_LOGIC;
  SIGNAL or_1544_nl : STD_LOGIC;
  SIGNAL or_1543_nl : STD_LOGIC;
  SIGNAL mux_1725_nl : STD_LOGIC;
  SIGNAL mux_1724_nl : STD_LOGIC;
  SIGNAL or_1561_nl : STD_LOGIC;
  SIGNAL or_1560_nl : STD_LOGIC;
  SIGNAL nand_429_nl : STD_LOGIC;
  SIGNAL or_1557_nl : STD_LOGIC;
  SIGNAL or_1564_nl : STD_LOGIC;
  SIGNAL or_1562_nl : STD_LOGIC;
  SIGNAL or_1644_nl : STD_LOGIC;
  SIGNAL mux_1781_nl : STD_LOGIC;
  SIGNAL or_1643_nl : STD_LOGIC;
  SIGNAL or_1642_nl : STD_LOGIC;
  SIGNAL mux_1786_nl : STD_LOGIC;
  SIGNAL mux_1785_nl : STD_LOGIC;
  SIGNAL or_1652_nl : STD_LOGIC;
  SIGNAL or_1651_nl : STD_LOGIC;
  SIGNAL nand_428_nl : STD_LOGIC;
  SIGNAL or_1648_nl : STD_LOGIC;
  SIGNAL or_1656_nl : STD_LOGIC;
  SIGNAL or_1654_nl : STD_LOGIC;
  SIGNAL or_1758_nl : STD_LOGIC;
  SIGNAL mux_1858_nl : STD_LOGIC;
  SIGNAL or_1757_nl : STD_LOGIC;
  SIGNAL or_1756_nl : STD_LOGIC;
  SIGNAL mux_1869_nl : STD_LOGIC;
  SIGNAL mux_1868_nl : STD_LOGIC;
  SIGNAL or_1774_nl : STD_LOGIC;
  SIGNAL or_1773_nl : STD_LOGIC;
  SIGNAL nand_427_nl : STD_LOGIC;
  SIGNAL or_1770_nl : STD_LOGIC;
  SIGNAL nand_416_nl : STD_LOGIC;
  SIGNAL or_1775_nl : STD_LOGIC;
  SIGNAL mux_1922_nl : STD_LOGIC;
  SIGNAL or_1853_nl : STD_LOGIC;
  SIGNAL or_1852_nl : STD_LOGIC;
  SIGNAL nand_73_nl : STD_LOGIC;
  SIGNAL mux_1926_nl : STD_LOGIC;
  SIGNAL nor_874_nl : STD_LOGIC;
  SIGNAL nor_875_nl : STD_LOGIC;
  SIGNAL or_1857_nl : STD_LOGIC;
  SIGNAL mux_1925_nl : STD_LOGIC;
  SIGNAL or_1856_nl : STD_LOGIC;
  SIGNAL or_1855_nl : STD_LOGIC;
  SIGNAL mux_1929_nl : STD_LOGIC;
  SIGNAL nor_872_nl : STD_LOGIC;
  SIGNAL nor_873_nl : STD_LOGIC;
  SIGNAL or_1974_nl : STD_LOGIC;
  SIGNAL mux_2003_nl : STD_LOGIC;
  SIGNAL or_1973_nl : STD_LOGIC;
  SIGNAL or_1972_nl : STD_LOGIC;
  SIGNAL mux_2014_nl : STD_LOGIC;
  SIGNAL mux_2013_nl : STD_LOGIC;
  SIGNAL or_1990_nl : STD_LOGIC;
  SIGNAL or_1989_nl : STD_LOGIC;
  SIGNAL nand_426_nl : STD_LOGIC;
  SIGNAL or_1986_nl : STD_LOGIC;
  SIGNAL nand_414_nl : STD_LOGIC;
  SIGNAL or_1991_nl : STD_LOGIC;
  SIGNAL or_2073_nl : STD_LOGIC;
  SIGNAL mux_2070_nl : STD_LOGIC;
  SIGNAL or_2072_nl : STD_LOGIC;
  SIGNAL or_2071_nl : STD_LOGIC;
  SIGNAL mux_2075_nl : STD_LOGIC;
  SIGNAL mux_2074_nl : STD_LOGIC;
  SIGNAL or_2081_nl : STD_LOGIC;
  SIGNAL or_2080_nl : STD_LOGIC;
  SIGNAL nand_425_nl : STD_LOGIC;
  SIGNAL or_2077_nl : STD_LOGIC;
  SIGNAL nand_412_nl : STD_LOGIC;
  SIGNAL or_2083_nl : STD_LOGIC;
  SIGNAL or_2187_nl : STD_LOGIC;
  SIGNAL mux_2147_nl : STD_LOGIC;
  SIGNAL nand_291_nl : STD_LOGIC;
  SIGNAL or_2185_nl : STD_LOGIC;
  SIGNAL mux_2158_nl : STD_LOGIC;
  SIGNAL mux_2157_nl : STD_LOGIC;
  SIGNAL nand_288_nl : STD_LOGIC;
  SIGNAL nand_289_nl : STD_LOGIC;
  SIGNAL nand_424_nl : STD_LOGIC;
  SIGNAL or_2199_nl : STD_LOGIC;
  SIGNAL nand_410_nl : STD_LOGIC;
  SIGNAL or_2204_nl : STD_LOGIC;
  SIGNAL mux_2240_nl : STD_LOGIC;
  SIGNAL mux_2289_nl : STD_LOGIC;
  SIGNAL mux_2310_nl : STD_LOGIC;
  SIGNAL or_2393_nl : STD_LOGIC;
  SIGNAL mux_2427_nl : STD_LOGIC;
  SIGNAL or_2409_nl : STD_LOGIC;
  SIGNAL mux_2474_nl : STD_LOGIC;
  SIGNAL mux_2473_nl : STD_LOGIC;
  SIGNAL or_2425_nl : STD_LOGIC;
  SIGNAL mux_2472_nl : STD_LOGIC;
  SIGNAL or_2424_nl : STD_LOGIC;
  SIGNAL mux_2471_nl : STD_LOGIC;
  SIGNAL mux_2470_nl : STD_LOGIC;
  SIGNAL or_3285_nl : STD_LOGIC;
  SIGNAL mux_2469_nl : STD_LOGIC;
  SIGNAL or_2419_nl : STD_LOGIC;
  SIGNAL mux_2468_nl : STD_LOGIC;
  SIGNAL or_2417_nl : STD_LOGIC;
  SIGNAL mux_2467_nl : STD_LOGIC;
  SIGNAL nand_111_nl : STD_LOGIC;
  SIGNAL mux_2465_nl : STD_LOGIC;
  SIGNAL or_2412_nl : STD_LOGIC;
  SIGNAL mux_2464_nl : STD_LOGIC;
  SIGNAL nand_110_nl : STD_LOGIC;
  SIGNAL mux_2462_nl : STD_LOGIC;
  SIGNAL nor_756_nl : STD_LOGIC;
  SIGNAL nor_757_nl : STD_LOGIC;
  SIGNAL mux_2488_nl : STD_LOGIC;
  SIGNAL mux_2487_nl : STD_LOGIC;
  SIGNAL mux_2486_nl : STD_LOGIC;
  SIGNAL nor_743_nl : STD_LOGIC;
  SIGNAL nor_744_nl : STD_LOGIC;
  SIGNAL nor_745_nl : STD_LOGIC;
  SIGNAL mux_3706_nl : STD_LOGIC;
  SIGNAL or_3233_nl : STD_LOGIC;
  SIGNAL or_3232_nl : STD_LOGIC;
  SIGNAL mux_2484_nl : STD_LOGIC;
  SIGNAL nor_746_nl : STD_LOGIC;
  SIGNAL mux_2483_nl : STD_LOGIC;
  SIGNAL or_2441_nl : STD_LOGIC;
  SIGNAL or_2439_nl : STD_LOGIC;
  SIGNAL and_558_nl : STD_LOGIC;
  SIGNAL mux_89_nl : STD_LOGIC;
  SIGNAL nor_1285_nl : STD_LOGIC;
  SIGNAL nor_1286_nl : STD_LOGIC;
  SIGNAL mux_2481_nl : STD_LOGIC;
  SIGNAL mux_2480_nl : STD_LOGIC;
  SIGNAL mux_2479_nl : STD_LOGIC;
  SIGNAL mux_2478_nl : STD_LOGIC;
  SIGNAL nor_750_nl : STD_LOGIC;
  SIGNAL nor_1278_nl : STD_LOGIC;
  SIGNAL and_796_nl : STD_LOGIC;
  SIGNAL mux_94_nl : STD_LOGIC;
  SIGNAL mux_93_nl : STD_LOGIC;
  SIGNAL nor_1280_nl : STD_LOGIC;
  SIGNAL nor_1281_nl : STD_LOGIC;
  SIGNAL mux_2492_nl : STD_LOGIC;
  SIGNAL mux_2491_nl : STD_LOGIC;
  SIGNAL mux_2490_nl : STD_LOGIC;
  SIGNAL or_463_nl : STD_LOGIC;
  SIGNAL mux_2496_nl : STD_LOGIC;
  SIGNAL nor_741_nl : STD_LOGIC;
  SIGNAL nor_742_nl : STD_LOGIC;
  SIGNAL or_2468_nl : STD_LOGIC;
  SIGNAL or_2489_nl : STD_LOGIC;
  SIGNAL nand_117_nl : STD_LOGIC;
  SIGNAL nor_719_nl : STD_LOGIC;
  SIGNAL or_2556_nl : STD_LOGIC;
  SIGNAL or_2555_nl : STD_LOGIC;
  SIGNAL mux_2756_nl : STD_LOGIC;
  SIGNAL mux_2755_nl : STD_LOGIC;
  SIGNAL mux_2754_nl : STD_LOGIC;
  SIGNAL nor_702_nl : STD_LOGIC;
  SIGNAL mux_2753_nl : STD_LOGIC;
  SIGNAL nor_704_nl : STD_LOGIC;
  SIGNAL nor_705_nl : STD_LOGIC;
  SIGNAL mux_2752_nl : STD_LOGIC;
  SIGNAL nor_706_nl : STD_LOGIC;
  SIGNAL mux_2751_nl : STD_LOGIC;
  SIGNAL nor_707_nl : STD_LOGIC;
  SIGNAL mux_2750_nl : STD_LOGIC;
  SIGNAL nor_708_nl : STD_LOGIC;
  SIGNAL nor_1296_nl : STD_LOGIC;
  SIGNAL mux_2749_nl : STD_LOGIC;
  SIGNAL mux_2748_nl : STD_LOGIC;
  SIGNAL nor_710_nl : STD_LOGIC;
  SIGNAL mux_2747_nl : STD_LOGIC;
  SIGNAL nor_711_nl : STD_LOGIC;
  SIGNAL nor_712_nl : STD_LOGIC;
  SIGNAL nor_713_nl : STD_LOGIC;
  SIGNAL mux_2745_nl : STD_LOGIC;
  SIGNAL or_2553_nl : STD_LOGIC;
  SIGNAL mux_74_nl : STD_LOGIC;
  SIGNAL or_53_nl : STD_LOGIC;
  SIGNAL or_51_nl : STD_LOGIC;
  SIGNAL nand_120_nl : STD_LOGIC;
  SIGNAL or_2578_nl : STD_LOGIC;
  SIGNAL or_2621_nl : STD_LOGIC;
  SIGNAL mux_2799_nl : STD_LOGIC;
  SIGNAL mux_2871_nl : STD_LOGIC;
  SIGNAL or_207_nl : STD_LOGIC;
  SIGNAL mux_2880_nl : STD_LOGIC;
  SIGNAL and_503_nl : STD_LOGIC;
  SIGNAL mux_2879_nl : STD_LOGIC;
  SIGNAL mux_2878_nl : STD_LOGIC;
  SIGNAL nor_672_nl : STD_LOGIC;
  SIGNAL nor_673_nl : STD_LOGIC;
  SIGNAL nor_674_nl : STD_LOGIC;
  SIGNAL mux_2877_nl : STD_LOGIC;
  SIGNAL or_2662_nl : STD_LOGIC;
  SIGNAL mux_2876_nl : STD_LOGIC;
  SIGNAL or_2659_nl : STD_LOGIC;
  SIGNAL mux_2875_nl : STD_LOGIC;
  SIGNAL mux_2874_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL mux_2873_nl : STD_LOGIC;
  SIGNAL and_505_nl : STD_LOGIC;
  SIGNAL mux_2872_nl : STD_LOGIC;
  SIGNAL nor_676_nl : STD_LOGIC;
  SIGNAL mux_2870_nl : STD_LOGIC;
  SIGNAL or_2647_nl : STD_LOGIC;
  SIGNAL mux_2902_nl : STD_LOGIC;
  SIGNAL mux_2901_nl : STD_LOGIC;
  SIGNAL and_498_nl : STD_LOGIC;
  SIGNAL mux_2900_nl : STD_LOGIC;
  SIGNAL nor_654_nl : STD_LOGIC;
  SIGNAL mux_2899_nl : STD_LOGIC;
  SIGNAL nor_655_nl : STD_LOGIC;
  SIGNAL nor_656_nl : STD_LOGIC;
  SIGNAL mux_2898_nl : STD_LOGIC;
  SIGNAL nor_657_nl : STD_LOGIC;
  SIGNAL and_499_nl : STD_LOGIC;
  SIGNAL mux_2897_nl : STD_LOGIC;
  SIGNAL nor_658_nl : STD_LOGIC;
  SIGNAL mux_2896_nl : STD_LOGIC;
  SIGNAL or_2699_nl : STD_LOGIC;
  SIGNAL mux_2895_nl : STD_LOGIC;
  SIGNAL nor_659_nl : STD_LOGIC;
  SIGNAL nor_660_nl : STD_LOGIC;
  SIGNAL mux_2894_nl : STD_LOGIC;
  SIGNAL mux_2893_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL mux_2892_nl : STD_LOGIC;
  SIGNAL or_2693_nl : STD_LOGIC;
  SIGNAL and_500_nl : STD_LOGIC;
  SIGNAL mux_2891_nl : STD_LOGIC;
  SIGNAL nor_662_nl : STD_LOGIC;
  SIGNAL nor_663_nl : STD_LOGIC;
  SIGNAL mux_2890_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL nor_665_nl : STD_LOGIC;
  SIGNAL mux_523_nl : STD_LOGIC;
  SIGNAL or_248_nl : STD_LOGIC;
  SIGNAL mux_2910_nl : STD_LOGIC;
  SIGNAL mux_2920_nl : STD_LOGIC;
  SIGNAL mux_520_nl : STD_LOGIC;
  SIGNAL mux_3168_nl : STD_LOGIC;
  SIGNAL nor_627_nl : STD_LOGIC;
  SIGNAL nor_628_nl : STD_LOGIC;
  SIGNAL or_3260_nl : STD_LOGIC;
  SIGNAL mux_3213_nl : STD_LOGIC;
  SIGNAL or_2886_nl : STD_LOGIC;
  SIGNAL nand_220_nl : STD_LOGIC;
  SIGNAL mux_3212_nl : STD_LOGIC;
  SIGNAL or_2882_nl : STD_LOGIC;
  SIGNAL mux_3235_nl : STD_LOGIC;
  SIGNAL or_2905_nl : STD_LOGIC;
  SIGNAL or_2904_nl : STD_LOGIC;
  SIGNAL mux_3279_nl : STD_LOGIC;
  SIGNAL and_436_nl : STD_LOGIC;
  SIGNAL mux_3368_nl : STD_LOGIC;
  SIGNAL mux_3354_nl : STD_LOGIC;
  SIGNAL mux_3353_nl : STD_LOGIC;
  SIGNAL mux_3352_nl : STD_LOGIC;
  SIGNAL mux_3351_nl : STD_LOGIC;
  SIGNAL mux_3350_nl : STD_LOGIC;
  SIGNAL mux_3382_nl : STD_LOGIC;
  SIGNAL mux_3381_nl : STD_LOGIC;
  SIGNAL mux_3380_nl : STD_LOGIC;
  SIGNAL and_417_nl : STD_LOGIC;
  SIGNAL mux_3378_nl : STD_LOGIC;
  SIGNAL mux_3377_nl : STD_LOGIC;
  SIGNAL nor_591_nl : STD_LOGIC;
  SIGNAL nor_1295_nl : STD_LOGIC;
  SIGNAL mux_3376_nl : STD_LOGIC;
  SIGNAL mux_3375_nl : STD_LOGIC;
  SIGNAL and_418_nl : STD_LOGIC;
  SIGNAL mux_3374_nl : STD_LOGIC;
  SIGNAL nor_594_nl : STD_LOGIC;
  SIGNAL nor_595_nl : STD_LOGIC;
  SIGNAL nor_596_nl : STD_LOGIC;
  SIGNAL mux_3372_nl : STD_LOGIC;
  SIGNAL mux_3371_nl : STD_LOGIC;
  SIGNAL nor_1287_nl : STD_LOGIC;
  SIGNAL and_419_nl : STD_LOGIC;
  SIGNAL or_3007_nl : STD_LOGIC;
  SIGNAL or_3006_nl : STD_LOGIC;
  SIGNAL mux_3409_nl : STD_LOGIC;
  SIGNAL nor_573_nl : STD_LOGIC;
  SIGNAL mux_3408_nl : STD_LOGIC;
  SIGNAL mux_3407_nl : STD_LOGIC;
  SIGNAL or_3037_nl : STD_LOGIC;
  SIGNAL mux_3406_nl : STD_LOGIC;
  SIGNAL mux_3421_nl : STD_LOGIC;
  SIGNAL nor_568_nl : STD_LOGIC;
  SIGNAL mux_3613_nl : STD_LOGIC;
  SIGNAL mux_2664_nl : STD_LOGIC;
  SIGNAL mux_2663_nl : STD_LOGIC;
  SIGNAL mux_2662_nl : STD_LOGIC;
  SIGNAL nor_724_nl : STD_LOGIC;
  SIGNAL mux_2661_nl : STD_LOGIC;
  SIGNAL and_521_nl : STD_LOGIC;
  SIGNAL or_2522_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_acc_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL and_139_nl : STD_LOGIC;
  SIGNAL mux_1044_nl : STD_LOGIC;
  SIGNAL mux_1043_nl : STD_LOGIC;
  SIGNAL nor_1194_nl : STD_LOGIC;
  SIGNAL mux_1042_nl : STD_LOGIC;
  SIGNAL or_533_nl : STD_LOGIC;
  SIGNAL or_532_nl : STD_LOGIC;
  SIGNAL mux_1041_nl : STD_LOGIC;
  SIGNAL or_531_nl : STD_LOGIC;
  SIGNAL mux_1040_nl : STD_LOGIC;
  SIGNAL nor_1195_nl : STD_LOGIC;
  SIGNAL mux_1039_nl : STD_LOGIC;
  SIGNAL or_527_nl : STD_LOGIC;
  SIGNAL mux_1038_nl : STD_LOGIC;
  SIGNAL mux_1037_nl : STD_LOGIC;
  SIGNAL or_524_nl : STD_LOGIC;
  SIGNAL or_523_nl : STD_LOGIC;
  SIGNAL and_660_nl : STD_LOGIC;
  SIGNAL mux_1036_nl : STD_LOGIC;
  SIGNAL mux_1035_nl : STD_LOGIC;
  SIGNAL nor_1196_nl : STD_LOGIC;
  SIGNAL nor_1197_nl : STD_LOGIC;
  SIGNAL nor_1198_nl : STD_LOGIC;
  SIGNAL mux_1034_nl : STD_LOGIC;
  SIGNAL nor_1199_nl : STD_LOGIC;
  SIGNAL mux_1033_nl : STD_LOGIC;
  SIGNAL mux_1032_nl : STD_LOGIC;
  SIGNAL or_516_nl : STD_LOGIC;
  SIGNAL or_514_nl : STD_LOGIC;
  SIGNAL mux_1031_nl : STD_LOGIC;
  SIGNAL and_661_nl : STD_LOGIC;
  SIGNAL mux_1030_nl : STD_LOGIC;
  SIGNAL or_512_nl : STD_LOGIC;
  SIGNAL nor_1200_nl : STD_LOGIC;
  SIGNAL and_145_nl : STD_LOGIC;
  SIGNAL and_153_nl : STD_LOGIC;
  SIGNAL mux_1046_nl : STD_LOGIC;
  SIGNAL nor_1191_nl : STD_LOGIC;
  SIGNAL nor_1192_nl : STD_LOGIC;
  SIGNAL and_162_nl : STD_LOGIC;
  SIGNAL mux_1047_nl : STD_LOGIC;
  SIGNAL nor_1189_nl : STD_LOGIC;
  SIGNAL nor_1190_nl : STD_LOGIC;
  SIGNAL and_170_nl : STD_LOGIC;
  SIGNAL mux_1048_nl : STD_LOGIC;
  SIGNAL nor_1187_nl : STD_LOGIC;
  SIGNAL nor_1188_nl : STD_LOGIC;
  SIGNAL and_179_nl : STD_LOGIC;
  SIGNAL and_188_nl : STD_LOGIC;
  SIGNAL mux_1050_nl : STD_LOGIC;
  SIGNAL nor_1185_nl : STD_LOGIC;
  SIGNAL nor_1186_nl : STD_LOGIC;
  SIGNAL and_197_nl : STD_LOGIC;
  SIGNAL mux_1051_nl : STD_LOGIC;
  SIGNAL nor_1183_nl : STD_LOGIC;
  SIGNAL nor_1184_nl : STD_LOGIC;
  SIGNAL and_205_nl : STD_LOGIC;
  SIGNAL mux_1052_nl : STD_LOGIC;
  SIGNAL nor_1181_nl : STD_LOGIC;
  SIGNAL nor_1182_nl : STD_LOGIC;
  SIGNAL and_211_nl : STD_LOGIC;
  SIGNAL mux_1053_nl : STD_LOGIC;
  SIGNAL nor_1179_nl : STD_LOGIC;
  SIGNAL nor_1180_nl : STD_LOGIC;
  SIGNAL and_220_nl : STD_LOGIC;
  SIGNAL mux_1054_nl : STD_LOGIC;
  SIGNAL nor_1177_nl : STD_LOGIC;
  SIGNAL nor_1178_nl : STD_LOGIC;
  SIGNAL and_231_nl : STD_LOGIC;
  SIGNAL and_238_nl : STD_LOGIC;
  SIGNAL mux_1055_nl : STD_LOGIC;
  SIGNAL nor_1175_nl : STD_LOGIC;
  SIGNAL nor_1176_nl : STD_LOGIC;
  SIGNAL and_246_nl : STD_LOGIC;
  SIGNAL mux_1056_nl : STD_LOGIC;
  SIGNAL and_817_nl : STD_LOGIC;
  SIGNAL nor_1174_nl : STD_LOGIC;
  SIGNAL and_253_nl : STD_LOGIC;
  SIGNAL mux_1057_nl : STD_LOGIC;
  SIGNAL and_657_nl : STD_LOGIC;
  SIGNAL nor_1172_nl : STD_LOGIC;
  SIGNAL and_261_nl : STD_LOGIC;
  SIGNAL mux_1098_nl : STD_LOGIC;
  SIGNAL mux_1097_nl : STD_LOGIC;
  SIGNAL mux_1096_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL mux_1094_nl : STD_LOGIC;
  SIGNAL mux_1093_nl : STD_LOGIC;
  SIGNAL or_624_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL mux_1090_nl : STD_LOGIC;
  SIGNAL or_615_nl : STD_LOGIC;
  SIGNAL mux_1089_nl : STD_LOGIC;
  SIGNAL mux_1085_nl : STD_LOGIC;
  SIGNAL mux_1084_nl : STD_LOGIC;
  SIGNAL mux_1083_nl : STD_LOGIC;
  SIGNAL mux_1082_nl : STD_LOGIC;
  SIGNAL or_605_nl : STD_LOGIC;
  SIGNAL mux_1081_nl : STD_LOGIC;
  SIGNAL mux_1079_nl : STD_LOGIC;
  SIGNAL mux_1078_nl : STD_LOGIC;
  SIGNAL mux_1077_nl : STD_LOGIC;
  SIGNAL mux_1076_nl : STD_LOGIC;
  SIGNAL or_602_nl : STD_LOGIC;
  SIGNAL mux_1075_nl : STD_LOGIC;
  SIGNAL mux_1074_nl : STD_LOGIC;
  SIGNAL or_597_nl : STD_LOGIC;
  SIGNAL mux_1072_nl : STD_LOGIC;
  SIGNAL mux_1071_nl : STD_LOGIC;
  SIGNAL mux_1070_nl : STD_LOGIC;
  SIGNAL or_594_nl : STD_LOGIC;
  SIGNAL mux_1069_nl : STD_LOGIC;
  SIGNAL or_592_nl : STD_LOGIC;
  SIGNAL or_588_nl : STD_LOGIC;
  SIGNAL mux_1064_nl : STD_LOGIC;
  SIGNAL mux_1063_nl : STD_LOGIC;
  SIGNAL or_581_nl : STD_LOGIC;
  SIGNAL or_580_nl : STD_LOGIC;
  SIGNAL mux_1060_nl : STD_LOGIC;
  SIGNAL mux_1059_nl : STD_LOGIC;
  SIGNAL mux_1058_nl : STD_LOGIC;
  SIGNAL or_573_nl : STD_LOGIC;
  SIGNAL or_570_nl : STD_LOGIC;
  SIGNAL or_569_nl : STD_LOGIC;
  SIGNAL mux_1128_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL and_654_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL nor_1147_nl : STD_LOGIC;
  SIGNAL mux_1125_nl : STD_LOGIC;
  SIGNAL nor_1149_nl : STD_LOGIC;
  SIGNAL mux_1124_nl : STD_LOGIC;
  SIGNAL nor_1150_nl : STD_LOGIC;
  SIGNAL mux_1123_nl : STD_LOGIC;
  SIGNAL or_670_nl : STD_LOGIC;
  SIGNAL or_669_nl : STD_LOGIC;
  SIGNAL mux_1122_nl : STD_LOGIC;
  SIGNAL nor_1151_nl : STD_LOGIC;
  SIGNAL nor_1152_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL mux_1120_nl : STD_LOGIC;
  SIGNAL nor_1153_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL nor_1154_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL or_661_nl : STD_LOGIC;
  SIGNAL or_659_nl : STD_LOGIC;
  SIGNAL nor_1155_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL nor_1156_nl : STD_LOGIC;
  SIGNAL and_655_nl : STD_LOGIC;
  SIGNAL mux_1116_nl : STD_LOGIC;
  SIGNAL nor_1157_nl : STD_LOGIC;
  SIGNAL mux_1115_nl : STD_LOGIC;
  SIGNAL nor_1158_nl : STD_LOGIC;
  SIGNAL mux_1114_nl : STD_LOGIC;
  SIGNAL mux_1113_nl : STD_LOGIC;
  SIGNAL nor_1160_nl : STD_LOGIC;
  SIGNAL mux_1112_nl : STD_LOGIC;
  SIGNAL mux_1111_nl : STD_LOGIC;
  SIGNAL or_650_nl : STD_LOGIC;
  SIGNAL or_649_nl : STD_LOGIC;
  SIGNAL mux_1110_nl : STD_LOGIC;
  SIGNAL or_648_nl : STD_LOGIC;
  SIGNAL or_646_nl : STD_LOGIC;
  SIGNAL mux_1109_nl : STD_LOGIC;
  SIGNAL mux_1108_nl : STD_LOGIC;
  SIGNAL nor_1161_nl : STD_LOGIC;
  SIGNAL nor_1162_nl : STD_LOGIC;
  SIGNAL mux_1107_nl : STD_LOGIC;
  SIGNAL or_641_nl : STD_LOGIC;
  SIGNAL mux_1106_nl : STD_LOGIC;
  SIGNAL nor_1163_nl : STD_LOGIC;
  SIGNAL nor_1164_nl : STD_LOGIC;
  SIGNAL mux_1105_nl : STD_LOGIC;
  SIGNAL nor_1165_nl : STD_LOGIC;
  SIGNAL mux_1104_nl : STD_LOGIC;
  SIGNAL mux_1103_nl : STD_LOGIC;
  SIGNAL or_635_nl : STD_LOGIC;
  SIGNAL mux_1102_nl : STD_LOGIC;
  SIGNAL or_633_nl : STD_LOGIC;
  SIGNAL or_630_nl : STD_LOGIC;
  SIGNAL mux_1101_nl : STD_LOGIC;
  SIGNAL and_656_nl : STD_LOGIC;
  SIGNAL mux_1100_nl : STD_LOGIC;
  SIGNAL nor_1166_nl : STD_LOGIC;
  SIGNAL mux_1099_nl : STD_LOGIC;
  SIGNAL nor_1167_nl : STD_LOGIC;
  SIGNAL nor_1168_nl : STD_LOGIC;
  SIGNAL nor_1169_nl : STD_LOGIC;
  SIGNAL mux_1170_nl : STD_LOGIC;
  SIGNAL mux_1169_nl : STD_LOGIC;
  SIGNAL mux_1168_nl : STD_LOGIC;
  SIGNAL mux_1167_nl : STD_LOGIC;
  SIGNAL or_730_nl : STD_LOGIC;
  SIGNAL mux_1166_nl : STD_LOGIC;
  SIGNAL or_728_nl : STD_LOGIC;
  SIGNAL or_727_nl : STD_LOGIC;
  SIGNAL mux_1165_nl : STD_LOGIC;
  SIGNAL mux_1164_nl : STD_LOGIC;
  SIGNAL or_726_nl : STD_LOGIC;
  SIGNAL or_725_nl : STD_LOGIC;
  SIGNAL mux_1163_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL or_724_nl : STD_LOGIC;
  SIGNAL or_723_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL mux_1159_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL mux_1157_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL or_722_nl : STD_LOGIC;
  SIGNAL mux_1154_nl : STD_LOGIC;
  SIGNAL mux_1153_nl : STD_LOGIC;
  SIGNAL or_713_nl : STD_LOGIC;
  SIGNAL mux_1151_nl : STD_LOGIC;
  SIGNAL mux_1144_nl : STD_LOGIC;
  SIGNAL mux_1143_nl : STD_LOGIC;
  SIGNAL mux_1142_nl : STD_LOGIC;
  SIGNAL mux_1141_nl : STD_LOGIC;
  SIGNAL or_694_nl : STD_LOGIC;
  SIGNAL mux_1140_nl : STD_LOGIC;
  SIGNAL mux_1136_nl : STD_LOGIC;
  SIGNAL mux_1135_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL or_685_nl : STD_LOGIC;
  SIGNAL mux_1132_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL or_678_nl : STD_LOGIC;
  SIGNAL nor_224_nl : STD_LOGIC;
  SIGNAL mux_1200_nl : STD_LOGIC;
  SIGNAL mux_1199_nl : STD_LOGIC;
  SIGNAL and_651_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL nor_1122_nl : STD_LOGIC;
  SIGNAL mux_1197_nl : STD_LOGIC;
  SIGNAL nor_1124_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL nor_1125_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL or_776_nl : STD_LOGIC;
  SIGNAL or_775_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL nor_1126_nl : STD_LOGIC;
  SIGNAL nor_1127_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL nor_1128_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL nor_1129_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL or_767_nl : STD_LOGIC;
  SIGNAL or_765_nl : STD_LOGIC;
  SIGNAL nor_1130_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL nor_1131_nl : STD_LOGIC;
  SIGNAL and_652_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL nor_1132_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL nor_1133_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL mux_1185_nl : STD_LOGIC;
  SIGNAL nor_1135_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL mux_1183_nl : STD_LOGIC;
  SIGNAL or_756_nl : STD_LOGIC;
  SIGNAL or_755_nl : STD_LOGIC;
  SIGNAL mux_1182_nl : STD_LOGIC;
  SIGNAL or_754_nl : STD_LOGIC;
  SIGNAL or_752_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL mux_1180_nl : STD_LOGIC;
  SIGNAL nor_1136_nl : STD_LOGIC;
  SIGNAL nor_1137_nl : STD_LOGIC;
  SIGNAL mux_1179_nl : STD_LOGIC;
  SIGNAL or_747_nl : STD_LOGIC;
  SIGNAL mux_1178_nl : STD_LOGIC;
  SIGNAL nor_1138_nl : STD_LOGIC;
  SIGNAL nor_1139_nl : STD_LOGIC;
  SIGNAL mux_1177_nl : STD_LOGIC;
  SIGNAL nor_1140_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL mux_1175_nl : STD_LOGIC;
  SIGNAL or_741_nl : STD_LOGIC;
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL or_739_nl : STD_LOGIC;
  SIGNAL or_736_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL and_653_nl : STD_LOGIC;
  SIGNAL mux_1172_nl : STD_LOGIC;
  SIGNAL nor_1141_nl : STD_LOGIC;
  SIGNAL mux_1171_nl : STD_LOGIC;
  SIGNAL nor_1142_nl : STD_LOGIC;
  SIGNAL nor_1143_nl : STD_LOGIC;
  SIGNAL nor_1144_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL mux_1239_nl : STD_LOGIC;
  SIGNAL mux_1238_nl : STD_LOGIC;
  SIGNAL mux_1237_nl : STD_LOGIC;
  SIGNAL or_837_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL or_828_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL mux_1229_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL mux_1226_nl : STD_LOGIC;
  SIGNAL or_818_nl : STD_LOGIC;
  SIGNAL mux_1225_nl : STD_LOGIC;
  SIGNAL mux_1223_nl : STD_LOGIC;
  SIGNAL mux_1222_nl : STD_LOGIC;
  SIGNAL mux_1221_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL mux_1219_nl : STD_LOGIC;
  SIGNAL mux_1218_nl : STD_LOGIC;
  SIGNAL or_810_nl : STD_LOGIC;
  SIGNAL mux_1216_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL mux_1214_nl : STD_LOGIC;
  SIGNAL or_807_nl : STD_LOGIC;
  SIGNAL mux_1213_nl : STD_LOGIC;
  SIGNAL or_805_nl : STD_LOGIC;
  SIGNAL or_801_nl : STD_LOGIC;
  SIGNAL mux_1208_nl : STD_LOGIC;
  SIGNAL mux_1207_nl : STD_LOGIC;
  SIGNAL or_794_nl : STD_LOGIC;
  SIGNAL or_793_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL mux_1203_nl : STD_LOGIC;
  SIGNAL mux_1202_nl : STD_LOGIC;
  SIGNAL or_786_nl : STD_LOGIC;
  SIGNAL or_783_nl : STD_LOGIC;
  SIGNAL or_782_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL and_648_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL nor_1097_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL nor_1099_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL nor_1100_nl : STD_LOGIC;
  SIGNAL mux_1267_nl : STD_LOGIC;
  SIGNAL or_883_nl : STD_LOGIC;
  SIGNAL or_882_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL nor_1101_nl : STD_LOGIC;
  SIGNAL nor_1102_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL nor_1103_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL nor_1104_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL or_874_nl : STD_LOGIC;
  SIGNAL or_872_nl : STD_LOGIC;
  SIGNAL nor_1105_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL nor_1106_nl : STD_LOGIC;
  SIGNAL and_649_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL nor_1107_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL nor_1108_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL nor_1110_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL or_863_nl : STD_LOGIC;
  SIGNAL or_862_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL or_861_nl : STD_LOGIC;
  SIGNAL or_859_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL nor_1111_nl : STD_LOGIC;
  SIGNAL nor_1112_nl : STD_LOGIC;
  SIGNAL mux_1251_nl : STD_LOGIC;
  SIGNAL or_854_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL nor_1113_nl : STD_LOGIC;
  SIGNAL nor_1114_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL nor_1115_nl : STD_LOGIC;
  SIGNAL mux_1248_nl : STD_LOGIC;
  SIGNAL mux_1247_nl : STD_LOGIC;
  SIGNAL or_848_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL or_846_nl : STD_LOGIC;
  SIGNAL or_843_nl : STD_LOGIC;
  SIGNAL mux_1245_nl : STD_LOGIC;
  SIGNAL and_650_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL nor_1116_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL nor_1117_nl : STD_LOGIC;
  SIGNAL nor_1118_nl : STD_LOGIC;
  SIGNAL nor_1119_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL or_943_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL or_941_nl : STD_LOGIC;
  SIGNAL or_940_nl : STD_LOGIC;
  SIGNAL mux_1309_nl : STD_LOGIC;
  SIGNAL mux_1308_nl : STD_LOGIC;
  SIGNAL or_939_nl : STD_LOGIC;
  SIGNAL or_938_nl : STD_LOGIC;
  SIGNAL mux_1307_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL mux_1305_nl : STD_LOGIC;
  SIGNAL or_937_nl : STD_LOGIC;
  SIGNAL or_936_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL mux_1303_nl : STD_LOGIC;
  SIGNAL mux_1302_nl : STD_LOGIC;
  SIGNAL mux_1301_nl : STD_LOGIC;
  SIGNAL mux_1300_nl : STD_LOGIC;
  SIGNAL or_935_nl : STD_LOGIC;
  SIGNAL mux_1298_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL or_926_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL mux_1287_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL mux_1285_nl : STD_LOGIC;
  SIGNAL or_907_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL mux_1278_nl : STD_LOGIC;
  SIGNAL mux_1277_nl : STD_LOGIC;
  SIGNAL or_898_nl : STD_LOGIC;
  SIGNAL mux_1276_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL or_891_nl : STD_LOGIC;
  SIGNAL nor_231_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL mux_1343_nl : STD_LOGIC;
  SIGNAL and_645_nl : STD_LOGIC;
  SIGNAL mux_1342_nl : STD_LOGIC;
  SIGNAL nor_1072_nl : STD_LOGIC;
  SIGNAL mux_1341_nl : STD_LOGIC;
  SIGNAL nor_1074_nl : STD_LOGIC;
  SIGNAL mux_1340_nl : STD_LOGIC;
  SIGNAL nor_1075_nl : STD_LOGIC;
  SIGNAL mux_1339_nl : STD_LOGIC;
  SIGNAL or_989_nl : STD_LOGIC;
  SIGNAL or_988_nl : STD_LOGIC;
  SIGNAL mux_1338_nl : STD_LOGIC;
  SIGNAL nor_1076_nl : STD_LOGIC;
  SIGNAL nor_1077_nl : STD_LOGIC;
  SIGNAL mux_1337_nl : STD_LOGIC;
  SIGNAL mux_1336_nl : STD_LOGIC;
  SIGNAL nor_1078_nl : STD_LOGIC;
  SIGNAL mux_1335_nl : STD_LOGIC;
  SIGNAL nor_1079_nl : STD_LOGIC;
  SIGNAL mux_1334_nl : STD_LOGIC;
  SIGNAL or_980_nl : STD_LOGIC;
  SIGNAL or_978_nl : STD_LOGIC;
  SIGNAL nor_1080_nl : STD_LOGIC;
  SIGNAL mux_1333_nl : STD_LOGIC;
  SIGNAL nor_1081_nl : STD_LOGIC;
  SIGNAL and_646_nl : STD_LOGIC;
  SIGNAL mux_1332_nl : STD_LOGIC;
  SIGNAL nor_1082_nl : STD_LOGIC;
  SIGNAL mux_1331_nl : STD_LOGIC;
  SIGNAL nor_1083_nl : STD_LOGIC;
  SIGNAL mux_1330_nl : STD_LOGIC;
  SIGNAL mux_1329_nl : STD_LOGIC;
  SIGNAL nor_1085_nl : STD_LOGIC;
  SIGNAL mux_1328_nl : STD_LOGIC;
  SIGNAL mux_1327_nl : STD_LOGIC;
  SIGNAL or_969_nl : STD_LOGIC;
  SIGNAL or_968_nl : STD_LOGIC;
  SIGNAL mux_1326_nl : STD_LOGIC;
  SIGNAL or_967_nl : STD_LOGIC;
  SIGNAL or_965_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL nor_1086_nl : STD_LOGIC;
  SIGNAL nor_1087_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL or_960_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL nor_1088_nl : STD_LOGIC;
  SIGNAL nor_1089_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL nor_1090_nl : STD_LOGIC;
  SIGNAL mux_1320_nl : STD_LOGIC;
  SIGNAL mux_1319_nl : STD_LOGIC;
  SIGNAL or_954_nl : STD_LOGIC;
  SIGNAL mux_1318_nl : STD_LOGIC;
  SIGNAL or_952_nl : STD_LOGIC;
  SIGNAL or_949_nl : STD_LOGIC;
  SIGNAL mux_1317_nl : STD_LOGIC;
  SIGNAL and_647_nl : STD_LOGIC;
  SIGNAL mux_1316_nl : STD_LOGIC;
  SIGNAL nor_1091_nl : STD_LOGIC;
  SIGNAL mux_1315_nl : STD_LOGIC;
  SIGNAL nor_1092_nl : STD_LOGIC;
  SIGNAL nor_1093_nl : STD_LOGIC;
  SIGNAL nor_1094_nl : STD_LOGIC;
  SIGNAL mux_1386_nl : STD_LOGIC;
  SIGNAL mux_1385_nl : STD_LOGIC;
  SIGNAL mux_1384_nl : STD_LOGIC;
  SIGNAL mux_1383_nl : STD_LOGIC;
  SIGNAL mux_1382_nl : STD_LOGIC;
  SIGNAL mux_1381_nl : STD_LOGIC;
  SIGNAL or_1050_nl : STD_LOGIC;
  SIGNAL mux_1379_nl : STD_LOGIC;
  SIGNAL mux_1378_nl : STD_LOGIC;
  SIGNAL or_1041_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL mux_1373_nl : STD_LOGIC;
  SIGNAL mux_1372_nl : STD_LOGIC;
  SIGNAL mux_1371_nl : STD_LOGIC;
  SIGNAL mux_1370_nl : STD_LOGIC;
  SIGNAL or_1031_nl : STD_LOGIC;
  SIGNAL mux_1369_nl : STD_LOGIC;
  SIGNAL mux_1367_nl : STD_LOGIC;
  SIGNAL mux_1366_nl : STD_LOGIC;
  SIGNAL mux_1365_nl : STD_LOGIC;
  SIGNAL mux_1364_nl : STD_LOGIC;
  SIGNAL or_1028_nl : STD_LOGIC;
  SIGNAL mux_1363_nl : STD_LOGIC;
  SIGNAL mux_1362_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL mux_1360_nl : STD_LOGIC;
  SIGNAL mux_1359_nl : STD_LOGIC;
  SIGNAL mux_1358_nl : STD_LOGIC;
  SIGNAL or_1020_nl : STD_LOGIC;
  SIGNAL mux_1357_nl : STD_LOGIC;
  SIGNAL or_1018_nl : STD_LOGIC;
  SIGNAL or_1014_nl : STD_LOGIC;
  SIGNAL mux_1352_nl : STD_LOGIC;
  SIGNAL mux_1351_nl : STD_LOGIC;
  SIGNAL or_1007_nl : STD_LOGIC;
  SIGNAL or_1006_nl : STD_LOGIC;
  SIGNAL mux_1348_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL or_999_nl : STD_LOGIC;
  SIGNAL or_996_nl : STD_LOGIC;
  SIGNAL or_995_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL and_642_nl : STD_LOGIC;
  SIGNAL mux_1414_nl : STD_LOGIC;
  SIGNAL nor_1047_nl : STD_LOGIC;
  SIGNAL mux_1413_nl : STD_LOGIC;
  SIGNAL nor_1049_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL nor_1050_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL or_1096_nl : STD_LOGIC;
  SIGNAL or_1095_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL nor_1051_nl : STD_LOGIC;
  SIGNAL nor_1052_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL nor_1053_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL nor_1054_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL or_1087_nl : STD_LOGIC;
  SIGNAL or_1085_nl : STD_LOGIC;
  SIGNAL nor_1055_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL nor_1056_nl : STD_LOGIC;
  SIGNAL and_643_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL nor_1057_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL nor_1058_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL nor_1060_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL or_1076_nl : STD_LOGIC;
  SIGNAL or_1075_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL or_1074_nl : STD_LOGIC;
  SIGNAL or_1072_nl : STD_LOGIC;
  SIGNAL mux_1397_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL nor_1061_nl : STD_LOGIC;
  SIGNAL nor_1062_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL or_1067_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL nor_1063_nl : STD_LOGIC;
  SIGNAL nor_1064_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL nor_1065_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL or_1061_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL or_1059_nl : STD_LOGIC;
  SIGNAL or_1056_nl : STD_LOGIC;
  SIGNAL mux_1389_nl : STD_LOGIC;
  SIGNAL and_644_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL nor_1066_nl : STD_LOGIC;
  SIGNAL mux_1387_nl : STD_LOGIC;
  SIGNAL nor_1067_nl : STD_LOGIC;
  SIGNAL nor_1068_nl : STD_LOGIC;
  SIGNAL nor_1069_nl : STD_LOGIC;
  SIGNAL mux_1458_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL or_1156_nl : STD_LOGIC;
  SIGNAL mux_1454_nl : STD_LOGIC;
  SIGNAL or_1154_nl : STD_LOGIC;
  SIGNAL or_1153_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL or_1152_nl : STD_LOGIC;
  SIGNAL or_1151_nl : STD_LOGIC;
  SIGNAL mux_1451_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL or_1150_nl : STD_LOGIC;
  SIGNAL or_1149_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL or_1148_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL mux_1441_nl : STD_LOGIC;
  SIGNAL or_1139_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL or_1120_nl : STD_LOGIC;
  SIGNAL mux_1428_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL mux_1421_nl : STD_LOGIC;
  SIGNAL or_1111_nl : STD_LOGIC;
  SIGNAL mux_1420_nl : STD_LOGIC;
  SIGNAL mux_1419_nl : STD_LOGIC;
  SIGNAL or_1104_nl : STD_LOGIC;
  SIGNAL nor_238_nl : STD_LOGIC;
  SIGNAL mux_1488_nl : STD_LOGIC;
  SIGNAL mux_1487_nl : STD_LOGIC;
  SIGNAL and_639_nl : STD_LOGIC;
  SIGNAL mux_1486_nl : STD_LOGIC;
  SIGNAL nor_1022_nl : STD_LOGIC;
  SIGNAL mux_1485_nl : STD_LOGIC;
  SIGNAL nor_1024_nl : STD_LOGIC;
  SIGNAL mux_1484_nl : STD_LOGIC;
  SIGNAL nor_1025_nl : STD_LOGIC;
  SIGNAL mux_1483_nl : STD_LOGIC;
  SIGNAL or_1202_nl : STD_LOGIC;
  SIGNAL or_1201_nl : STD_LOGIC;
  SIGNAL mux_1482_nl : STD_LOGIC;
  SIGNAL nor_1026_nl : STD_LOGIC;
  SIGNAL nor_1027_nl : STD_LOGIC;
  SIGNAL mux_1481_nl : STD_LOGIC;
  SIGNAL mux_1480_nl : STD_LOGIC;
  SIGNAL nor_1028_nl : STD_LOGIC;
  SIGNAL mux_1479_nl : STD_LOGIC;
  SIGNAL nor_1029_nl : STD_LOGIC;
  SIGNAL mux_1478_nl : STD_LOGIC;
  SIGNAL or_1193_nl : STD_LOGIC;
  SIGNAL or_1191_nl : STD_LOGIC;
  SIGNAL nor_1030_nl : STD_LOGIC;
  SIGNAL mux_1477_nl : STD_LOGIC;
  SIGNAL nor_1031_nl : STD_LOGIC;
  SIGNAL and_640_nl : STD_LOGIC;
  SIGNAL mux_1476_nl : STD_LOGIC;
  SIGNAL nor_1032_nl : STD_LOGIC;
  SIGNAL mux_1475_nl : STD_LOGIC;
  SIGNAL nor_1033_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL nor_1035_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL or_1182_nl : STD_LOGIC;
  SIGNAL or_1181_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL or_1180_nl : STD_LOGIC;
  SIGNAL or_1178_nl : STD_LOGIC;
  SIGNAL mux_1469_nl : STD_LOGIC;
  SIGNAL mux_1468_nl : STD_LOGIC;
  SIGNAL nor_1036_nl : STD_LOGIC;
  SIGNAL nor_1037_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL or_1173_nl : STD_LOGIC;
  SIGNAL mux_1466_nl : STD_LOGIC;
  SIGNAL nor_1038_nl : STD_LOGIC;
  SIGNAL nor_1039_nl : STD_LOGIC;
  SIGNAL mux_1465_nl : STD_LOGIC;
  SIGNAL nor_1040_nl : STD_LOGIC;
  SIGNAL mux_1464_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL or_1167_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL or_1165_nl : STD_LOGIC;
  SIGNAL or_1162_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL and_641_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL nor_1041_nl : STD_LOGIC;
  SIGNAL mux_1459_nl : STD_LOGIC;
  SIGNAL nor_1042_nl : STD_LOGIC;
  SIGNAL nor_1043_nl : STD_LOGIC;
  SIGNAL nor_1044_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL mux_1529_nl : STD_LOGIC;
  SIGNAL mux_1528_nl : STD_LOGIC;
  SIGNAL mux_1527_nl : STD_LOGIC;
  SIGNAL mux_1526_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL or_1263_nl : STD_LOGIC;
  SIGNAL mux_1523_nl : STD_LOGIC;
  SIGNAL mux_1522_nl : STD_LOGIC;
  SIGNAL or_1254_nl : STD_LOGIC;
  SIGNAL mux_1521_nl : STD_LOGIC;
  SIGNAL mux_1517_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL mux_1515_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL or_1244_nl : STD_LOGIC;
  SIGNAL mux_1513_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL or_1241_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL mux_1506_nl : STD_LOGIC;
  SIGNAL or_1236_nl : STD_LOGIC;
  SIGNAL mux_1504_nl : STD_LOGIC;
  SIGNAL mux_1503_nl : STD_LOGIC;
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL or_1233_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL or_1231_nl : STD_LOGIC;
  SIGNAL or_1227_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL mux_1495_nl : STD_LOGIC;
  SIGNAL or_1220_nl : STD_LOGIC;
  SIGNAL or_1219_nl : STD_LOGIC;
  SIGNAL mux_1492_nl : STD_LOGIC;
  SIGNAL mux_1491_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL or_1212_nl : STD_LOGIC;
  SIGNAL or_1209_nl : STD_LOGIC;
  SIGNAL or_1208_nl : STD_LOGIC;
  SIGNAL mux_1560_nl : STD_LOGIC;
  SIGNAL mux_1559_nl : STD_LOGIC;
  SIGNAL and_636_nl : STD_LOGIC;
  SIGNAL mux_1558_nl : STD_LOGIC;
  SIGNAL nor_997_nl : STD_LOGIC;
  SIGNAL mux_1557_nl : STD_LOGIC;
  SIGNAL nor_999_nl : STD_LOGIC;
  SIGNAL mux_1556_nl : STD_LOGIC;
  SIGNAL nor_1000_nl : STD_LOGIC;
  SIGNAL mux_1555_nl : STD_LOGIC;
  SIGNAL or_1309_nl : STD_LOGIC;
  SIGNAL or_1308_nl : STD_LOGIC;
  SIGNAL mux_1554_nl : STD_LOGIC;
  SIGNAL nor_1001_nl : STD_LOGIC;
  SIGNAL nor_1002_nl : STD_LOGIC;
  SIGNAL mux_1553_nl : STD_LOGIC;
  SIGNAL mux_1552_nl : STD_LOGIC;
  SIGNAL nor_1003_nl : STD_LOGIC;
  SIGNAL mux_1551_nl : STD_LOGIC;
  SIGNAL nor_1004_nl : STD_LOGIC;
  SIGNAL mux_1550_nl : STD_LOGIC;
  SIGNAL or_1300_nl : STD_LOGIC;
  SIGNAL or_1298_nl : STD_LOGIC;
  SIGNAL nor_1005_nl : STD_LOGIC;
  SIGNAL mux_1549_nl : STD_LOGIC;
  SIGNAL nor_1006_nl : STD_LOGIC;
  SIGNAL and_637_nl : STD_LOGIC;
  SIGNAL mux_1548_nl : STD_LOGIC;
  SIGNAL nor_1007_nl : STD_LOGIC;
  SIGNAL mux_1547_nl : STD_LOGIC;
  SIGNAL nor_1008_nl : STD_LOGIC;
  SIGNAL mux_1546_nl : STD_LOGIC;
  SIGNAL mux_1545_nl : STD_LOGIC;
  SIGNAL nor_1010_nl : STD_LOGIC;
  SIGNAL mux_1544_nl : STD_LOGIC;
  SIGNAL mux_1543_nl : STD_LOGIC;
  SIGNAL or_1289_nl : STD_LOGIC;
  SIGNAL or_1288_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL or_1287_nl : STD_LOGIC;
  SIGNAL or_1285_nl : STD_LOGIC;
  SIGNAL mux_1541_nl : STD_LOGIC;
  SIGNAL mux_1540_nl : STD_LOGIC;
  SIGNAL nor_1011_nl : STD_LOGIC;
  SIGNAL nor_1012_nl : STD_LOGIC;
  SIGNAL mux_1539_nl : STD_LOGIC;
  SIGNAL or_1280_nl : STD_LOGIC;
  SIGNAL mux_1538_nl : STD_LOGIC;
  SIGNAL nor_1013_nl : STD_LOGIC;
  SIGNAL nor_1014_nl : STD_LOGIC;
  SIGNAL mux_1537_nl : STD_LOGIC;
  SIGNAL nor_1015_nl : STD_LOGIC;
  SIGNAL mux_1536_nl : STD_LOGIC;
  SIGNAL mux_1535_nl : STD_LOGIC;
  SIGNAL or_1274_nl : STD_LOGIC;
  SIGNAL mux_1534_nl : STD_LOGIC;
  SIGNAL or_1272_nl : STD_LOGIC;
  SIGNAL or_1269_nl : STD_LOGIC;
  SIGNAL mux_1533_nl : STD_LOGIC;
  SIGNAL and_638_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL nor_1016_nl : STD_LOGIC;
  SIGNAL mux_1531_nl : STD_LOGIC;
  SIGNAL nor_1017_nl : STD_LOGIC;
  SIGNAL nor_1018_nl : STD_LOGIC;
  SIGNAL nor_1019_nl : STD_LOGIC;
  SIGNAL mux_1602_nl : STD_LOGIC;
  SIGNAL mux_1601_nl : STD_LOGIC;
  SIGNAL mux_1600_nl : STD_LOGIC;
  SIGNAL mux_1599_nl : STD_LOGIC;
  SIGNAL or_1369_nl : STD_LOGIC;
  SIGNAL mux_1598_nl : STD_LOGIC;
  SIGNAL or_1367_nl : STD_LOGIC;
  SIGNAL or_1366_nl : STD_LOGIC;
  SIGNAL mux_1597_nl : STD_LOGIC;
  SIGNAL mux_1596_nl : STD_LOGIC;
  SIGNAL nand_336_nl : STD_LOGIC;
  SIGNAL or_1364_nl : STD_LOGIC;
  SIGNAL mux_1595_nl : STD_LOGIC;
  SIGNAL mux_1594_nl : STD_LOGIC;
  SIGNAL mux_1593_nl : STD_LOGIC;
  SIGNAL or_1363_nl : STD_LOGIC;
  SIGNAL or_1362_nl : STD_LOGIC;
  SIGNAL mux_1592_nl : STD_LOGIC;
  SIGNAL mux_1591_nl : STD_LOGIC;
  SIGNAL mux_1590_nl : STD_LOGIC;
  SIGNAL mux_1589_nl : STD_LOGIC;
  SIGNAL mux_1588_nl : STD_LOGIC;
  SIGNAL or_1361_nl : STD_LOGIC;
  SIGNAL mux_1586_nl : STD_LOGIC;
  SIGNAL mux_1585_nl : STD_LOGIC;
  SIGNAL or_1352_nl : STD_LOGIC;
  SIGNAL mux_1583_nl : STD_LOGIC;
  SIGNAL mux_1576_nl : STD_LOGIC;
  SIGNAL mux_1575_nl : STD_LOGIC;
  SIGNAL mux_1574_nl : STD_LOGIC;
  SIGNAL mux_1573_nl : STD_LOGIC;
  SIGNAL nand_338_nl : STD_LOGIC;
  SIGNAL mux_1572_nl : STD_LOGIC;
  SIGNAL mux_1568_nl : STD_LOGIC;
  SIGNAL mux_1567_nl : STD_LOGIC;
  SIGNAL mux_1566_nl : STD_LOGIC;
  SIGNAL mux_1565_nl : STD_LOGIC;
  SIGNAL or_1324_nl : STD_LOGIC;
  SIGNAL mux_1564_nl : STD_LOGIC;
  SIGNAL mux_1563_nl : STD_LOGIC;
  SIGNAL or_1317_nl : STD_LOGIC;
  SIGNAL and_635_nl : STD_LOGIC;
  SIGNAL mux_1632_nl : STD_LOGIC;
  SIGNAL mux_1631_nl : STD_LOGIC;
  SIGNAL and_630_nl : STD_LOGIC;
  SIGNAL mux_1630_nl : STD_LOGIC;
  SIGNAL nor_974_nl : STD_LOGIC;
  SIGNAL mux_1629_nl : STD_LOGIC;
  SIGNAL nor_976_nl : STD_LOGIC;
  SIGNAL mux_1628_nl : STD_LOGIC;
  SIGNAL nor_977_nl : STD_LOGIC;
  SIGNAL mux_1627_nl : STD_LOGIC;
  SIGNAL nand_333_nl : STD_LOGIC;
  SIGNAL or_1414_nl : STD_LOGIC;
  SIGNAL mux_1626_nl : STD_LOGIC;
  SIGNAL nor_978_nl : STD_LOGIC;
  SIGNAL nor_979_nl : STD_LOGIC;
  SIGNAL mux_1625_nl : STD_LOGIC;
  SIGNAL mux_1624_nl : STD_LOGIC;
  SIGNAL and_631_nl : STD_LOGIC;
  SIGNAL mux_1623_nl : STD_LOGIC;
  SIGNAL nor_980_nl : STD_LOGIC;
  SIGNAL mux_1622_nl : STD_LOGIC;
  SIGNAL or_1406_nl : STD_LOGIC;
  SIGNAL or_1404_nl : STD_LOGIC;
  SIGNAL nor_981_nl : STD_LOGIC;
  SIGNAL mux_1621_nl : STD_LOGIC;
  SIGNAL nor_982_nl : STD_LOGIC;
  SIGNAL and_632_nl : STD_LOGIC;
  SIGNAL mux_1620_nl : STD_LOGIC;
  SIGNAL and_828_nl : STD_LOGIC;
  SIGNAL mux_1619_nl : STD_LOGIC;
  SIGNAL nor_984_nl : STD_LOGIC;
  SIGNAL mux_1618_nl : STD_LOGIC;
  SIGNAL mux_1617_nl : STD_LOGIC;
  SIGNAL nor_986_nl : STD_LOGIC;
  SIGNAL mux_1616_nl : STD_LOGIC;
  SIGNAL mux_1615_nl : STD_LOGIC;
  SIGNAL or_1395_nl : STD_LOGIC;
  SIGNAL or_1394_nl : STD_LOGIC;
  SIGNAL mux_1614_nl : STD_LOGIC;
  SIGNAL or_1393_nl : STD_LOGIC;
  SIGNAL or_1391_nl : STD_LOGIC;
  SIGNAL mux_1613_nl : STD_LOGIC;
  SIGNAL mux_1612_nl : STD_LOGIC;
  SIGNAL nor_987_nl : STD_LOGIC;
  SIGNAL nor_988_nl : STD_LOGIC;
  SIGNAL mux_1611_nl : STD_LOGIC;
  SIGNAL or_1386_nl : STD_LOGIC;
  SIGNAL mux_1610_nl : STD_LOGIC;
  SIGNAL nor_989_nl : STD_LOGIC;
  SIGNAL nor_990_nl : STD_LOGIC;
  SIGNAL mux_1609_nl : STD_LOGIC;
  SIGNAL nor_991_nl : STD_LOGIC;
  SIGNAL mux_1608_nl : STD_LOGIC;
  SIGNAL mux_1607_nl : STD_LOGIC;
  SIGNAL nand_417_nl : STD_LOGIC;
  SIGNAL mux_1606_nl : STD_LOGIC;
  SIGNAL or_1378_nl : STD_LOGIC;
  SIGNAL or_1375_nl : STD_LOGIC;
  SIGNAL mux_1605_nl : STD_LOGIC;
  SIGNAL and_633_nl : STD_LOGIC;
  SIGNAL mux_1604_nl : STD_LOGIC;
  SIGNAL nor_992_nl : STD_LOGIC;
  SIGNAL mux_1603_nl : STD_LOGIC;
  SIGNAL and_634_nl : STD_LOGIC;
  SIGNAL nor_993_nl : STD_LOGIC;
  SIGNAL nor_994_nl : STD_LOGIC;
  SIGNAL mux_1674_nl : STD_LOGIC;
  SIGNAL mux_1673_nl : STD_LOGIC;
  SIGNAL mux_1672_nl : STD_LOGIC;
  SIGNAL mux_1671_nl : STD_LOGIC;
  SIGNAL mux_1670_nl : STD_LOGIC;
  SIGNAL mux_1669_nl : STD_LOGIC;
  SIGNAL or_1476_nl : STD_LOGIC;
  SIGNAL mux_1667_nl : STD_LOGIC;
  SIGNAL mux_1666_nl : STD_LOGIC;
  SIGNAL or_1467_nl : STD_LOGIC;
  SIGNAL mux_1665_nl : STD_LOGIC;
  SIGNAL mux_1661_nl : STD_LOGIC;
  SIGNAL mux_1660_nl : STD_LOGIC;
  SIGNAL mux_1659_nl : STD_LOGIC;
  SIGNAL mux_1658_nl : STD_LOGIC;
  SIGNAL or_1457_nl : STD_LOGIC;
  SIGNAL mux_1657_nl : STD_LOGIC;
  SIGNAL mux_1655_nl : STD_LOGIC;
  SIGNAL mux_1654_nl : STD_LOGIC;
  SIGNAL mux_1653_nl : STD_LOGIC;
  SIGNAL mux_1652_nl : STD_LOGIC;
  SIGNAL or_1454_nl : STD_LOGIC;
  SIGNAL mux_1651_nl : STD_LOGIC;
  SIGNAL mux_1650_nl : STD_LOGIC;
  SIGNAL or_1449_nl : STD_LOGIC;
  SIGNAL mux_1648_nl : STD_LOGIC;
  SIGNAL mux_1647_nl : STD_LOGIC;
  SIGNAL mux_1646_nl : STD_LOGIC;
  SIGNAL or_1446_nl : STD_LOGIC;
  SIGNAL mux_1645_nl : STD_LOGIC;
  SIGNAL or_1444_nl : STD_LOGIC;
  SIGNAL or_1440_nl : STD_LOGIC;
  SIGNAL mux_1640_nl : STD_LOGIC;
  SIGNAL mux_1639_nl : STD_LOGIC;
  SIGNAL or_1433_nl : STD_LOGIC;
  SIGNAL or_1432_nl : STD_LOGIC;
  SIGNAL mux_1636_nl : STD_LOGIC;
  SIGNAL mux_1635_nl : STD_LOGIC;
  SIGNAL mux_1634_nl : STD_LOGIC;
  SIGNAL or_1425_nl : STD_LOGIC;
  SIGNAL or_1422_nl : STD_LOGIC;
  SIGNAL or_1421_nl : STD_LOGIC;
  SIGNAL mux_1704_nl : STD_LOGIC;
  SIGNAL mux_1703_nl : STD_LOGIC;
  SIGNAL and_627_nl : STD_LOGIC;
  SIGNAL mux_1702_nl : STD_LOGIC;
  SIGNAL nor_949_nl : STD_LOGIC;
  SIGNAL mux_1701_nl : STD_LOGIC;
  SIGNAL nor_951_nl : STD_LOGIC;
  SIGNAL mux_1700_nl : STD_LOGIC;
  SIGNAL nor_952_nl : STD_LOGIC;
  SIGNAL mux_1699_nl : STD_LOGIC;
  SIGNAL or_1522_nl : STD_LOGIC;
  SIGNAL or_1521_nl : STD_LOGIC;
  SIGNAL mux_1698_nl : STD_LOGIC;
  SIGNAL nor_953_nl : STD_LOGIC;
  SIGNAL nor_954_nl : STD_LOGIC;
  SIGNAL mux_1697_nl : STD_LOGIC;
  SIGNAL mux_1696_nl : STD_LOGIC;
  SIGNAL nor_955_nl : STD_LOGIC;
  SIGNAL mux_1695_nl : STD_LOGIC;
  SIGNAL nor_956_nl : STD_LOGIC;
  SIGNAL mux_1694_nl : STD_LOGIC;
  SIGNAL or_1513_nl : STD_LOGIC;
  SIGNAL or_1511_nl : STD_LOGIC;
  SIGNAL nor_957_nl : STD_LOGIC;
  SIGNAL mux_1693_nl : STD_LOGIC;
  SIGNAL nor_958_nl : STD_LOGIC;
  SIGNAL and_628_nl : STD_LOGIC;
  SIGNAL mux_1692_nl : STD_LOGIC;
  SIGNAL nor_959_nl : STD_LOGIC;
  SIGNAL mux_1691_nl : STD_LOGIC;
  SIGNAL nor_960_nl : STD_LOGIC;
  SIGNAL mux_1690_nl : STD_LOGIC;
  SIGNAL mux_1689_nl : STD_LOGIC;
  SIGNAL nor_962_nl : STD_LOGIC;
  SIGNAL mux_1688_nl : STD_LOGIC;
  SIGNAL mux_1687_nl : STD_LOGIC;
  SIGNAL or_1502_nl : STD_LOGIC;
  SIGNAL or_1501_nl : STD_LOGIC;
  SIGNAL mux_1686_nl : STD_LOGIC;
  SIGNAL or_1500_nl : STD_LOGIC;
  SIGNAL or_1498_nl : STD_LOGIC;
  SIGNAL mux_1685_nl : STD_LOGIC;
  SIGNAL mux_1684_nl : STD_LOGIC;
  SIGNAL nor_963_nl : STD_LOGIC;
  SIGNAL nor_964_nl : STD_LOGIC;
  SIGNAL mux_1683_nl : STD_LOGIC;
  SIGNAL or_1493_nl : STD_LOGIC;
  SIGNAL mux_1682_nl : STD_LOGIC;
  SIGNAL nor_965_nl : STD_LOGIC;
  SIGNAL nor_966_nl : STD_LOGIC;
  SIGNAL mux_1681_nl : STD_LOGIC;
  SIGNAL nor_967_nl : STD_LOGIC;
  SIGNAL mux_1680_nl : STD_LOGIC;
  SIGNAL mux_1679_nl : STD_LOGIC;
  SIGNAL or_1487_nl : STD_LOGIC;
  SIGNAL mux_1678_nl : STD_LOGIC;
  SIGNAL or_1485_nl : STD_LOGIC;
  SIGNAL or_1482_nl : STD_LOGIC;
  SIGNAL mux_1677_nl : STD_LOGIC;
  SIGNAL and_629_nl : STD_LOGIC;
  SIGNAL mux_1676_nl : STD_LOGIC;
  SIGNAL nor_968_nl : STD_LOGIC;
  SIGNAL mux_1675_nl : STD_LOGIC;
  SIGNAL nor_969_nl : STD_LOGIC;
  SIGNAL nor_970_nl : STD_LOGIC;
  SIGNAL nor_971_nl : STD_LOGIC;
  SIGNAL mux_1746_nl : STD_LOGIC;
  SIGNAL mux_1745_nl : STD_LOGIC;
  SIGNAL mux_1744_nl : STD_LOGIC;
  SIGNAL mux_1743_nl : STD_LOGIC;
  SIGNAL or_1582_nl : STD_LOGIC;
  SIGNAL mux_1742_nl : STD_LOGIC;
  SIGNAL or_1580_nl : STD_LOGIC;
  SIGNAL or_1579_nl : STD_LOGIC;
  SIGNAL mux_1741_nl : STD_LOGIC;
  SIGNAL mux_1740_nl : STD_LOGIC;
  SIGNAL or_1578_nl : STD_LOGIC;
  SIGNAL or_1577_nl : STD_LOGIC;
  SIGNAL mux_1739_nl : STD_LOGIC;
  SIGNAL mux_1738_nl : STD_LOGIC;
  SIGNAL mux_1737_nl : STD_LOGIC;
  SIGNAL or_1576_nl : STD_LOGIC;
  SIGNAL or_1575_nl : STD_LOGIC;
  SIGNAL mux_1736_nl : STD_LOGIC;
  SIGNAL mux_1735_nl : STD_LOGIC;
  SIGNAL mux_1734_nl : STD_LOGIC;
  SIGNAL mux_1733_nl : STD_LOGIC;
  SIGNAL mux_1732_nl : STD_LOGIC;
  SIGNAL or_1574_nl : STD_LOGIC;
  SIGNAL mux_1730_nl : STD_LOGIC;
  SIGNAL mux_1729_nl : STD_LOGIC;
  SIGNAL or_1565_nl : STD_LOGIC;
  SIGNAL mux_1727_nl : STD_LOGIC;
  SIGNAL mux_1720_nl : STD_LOGIC;
  SIGNAL mux_1719_nl : STD_LOGIC;
  SIGNAL mux_1718_nl : STD_LOGIC;
  SIGNAL mux_1717_nl : STD_LOGIC;
  SIGNAL or_1546_nl : STD_LOGIC;
  SIGNAL mux_1716_nl : STD_LOGIC;
  SIGNAL mux_1712_nl : STD_LOGIC;
  SIGNAL mux_1711_nl : STD_LOGIC;
  SIGNAL mux_1710_nl : STD_LOGIC;
  SIGNAL mux_1709_nl : STD_LOGIC;
  SIGNAL or_1537_nl : STD_LOGIC;
  SIGNAL mux_1708_nl : STD_LOGIC;
  SIGNAL mux_1707_nl : STD_LOGIC;
  SIGNAL or_1530_nl : STD_LOGIC;
  SIGNAL nor_252_nl : STD_LOGIC;
  SIGNAL mux_1776_nl : STD_LOGIC;
  SIGNAL mux_1775_nl : STD_LOGIC;
  SIGNAL and_624_nl : STD_LOGIC;
  SIGNAL mux_1774_nl : STD_LOGIC;
  SIGNAL nor_924_nl : STD_LOGIC;
  SIGNAL mux_1773_nl : STD_LOGIC;
  SIGNAL nor_926_nl : STD_LOGIC;
  SIGNAL mux_1772_nl : STD_LOGIC;
  SIGNAL nor_927_nl : STD_LOGIC;
  SIGNAL mux_1771_nl : STD_LOGIC;
  SIGNAL or_1628_nl : STD_LOGIC;
  SIGNAL or_1627_nl : STD_LOGIC;
  SIGNAL mux_1770_nl : STD_LOGIC;
  SIGNAL nor_928_nl : STD_LOGIC;
  SIGNAL nor_929_nl : STD_LOGIC;
  SIGNAL mux_1769_nl : STD_LOGIC;
  SIGNAL mux_1768_nl : STD_LOGIC;
  SIGNAL nor_930_nl : STD_LOGIC;
  SIGNAL mux_1767_nl : STD_LOGIC;
  SIGNAL nor_931_nl : STD_LOGIC;
  SIGNAL mux_1766_nl : STD_LOGIC;
  SIGNAL or_1619_nl : STD_LOGIC;
  SIGNAL or_1617_nl : STD_LOGIC;
  SIGNAL nor_932_nl : STD_LOGIC;
  SIGNAL mux_1765_nl : STD_LOGIC;
  SIGNAL nor_933_nl : STD_LOGIC;
  SIGNAL and_625_nl : STD_LOGIC;
  SIGNAL mux_1764_nl : STD_LOGIC;
  SIGNAL nor_934_nl : STD_LOGIC;
  SIGNAL mux_1763_nl : STD_LOGIC;
  SIGNAL nor_935_nl : STD_LOGIC;
  SIGNAL mux_1762_nl : STD_LOGIC;
  SIGNAL mux_1761_nl : STD_LOGIC;
  SIGNAL nor_937_nl : STD_LOGIC;
  SIGNAL mux_1760_nl : STD_LOGIC;
  SIGNAL mux_1759_nl : STD_LOGIC;
  SIGNAL or_1608_nl : STD_LOGIC;
  SIGNAL or_1607_nl : STD_LOGIC;
  SIGNAL mux_1758_nl : STD_LOGIC;
  SIGNAL or_1606_nl : STD_LOGIC;
  SIGNAL or_1604_nl : STD_LOGIC;
  SIGNAL mux_1757_nl : STD_LOGIC;
  SIGNAL mux_1756_nl : STD_LOGIC;
  SIGNAL nor_938_nl : STD_LOGIC;
  SIGNAL nor_939_nl : STD_LOGIC;
  SIGNAL mux_1755_nl : STD_LOGIC;
  SIGNAL or_1599_nl : STD_LOGIC;
  SIGNAL mux_1754_nl : STD_LOGIC;
  SIGNAL nor_940_nl : STD_LOGIC;
  SIGNAL nor_941_nl : STD_LOGIC;
  SIGNAL mux_1753_nl : STD_LOGIC;
  SIGNAL nor_942_nl : STD_LOGIC;
  SIGNAL mux_1752_nl : STD_LOGIC;
  SIGNAL mux_1751_nl : STD_LOGIC;
  SIGNAL or_1593_nl : STD_LOGIC;
  SIGNAL mux_1750_nl : STD_LOGIC;
  SIGNAL or_1591_nl : STD_LOGIC;
  SIGNAL or_1588_nl : STD_LOGIC;
  SIGNAL mux_1749_nl : STD_LOGIC;
  SIGNAL and_626_nl : STD_LOGIC;
  SIGNAL mux_1748_nl : STD_LOGIC;
  SIGNAL nor_943_nl : STD_LOGIC;
  SIGNAL mux_1747_nl : STD_LOGIC;
  SIGNAL nor_944_nl : STD_LOGIC;
  SIGNAL nor_945_nl : STD_LOGIC;
  SIGNAL nor_946_nl : STD_LOGIC;
  SIGNAL mux_1818_nl : STD_LOGIC;
  SIGNAL mux_1817_nl : STD_LOGIC;
  SIGNAL mux_1816_nl : STD_LOGIC;
  SIGNAL mux_1815_nl : STD_LOGIC;
  SIGNAL mux_1814_nl : STD_LOGIC;
  SIGNAL mux_1813_nl : STD_LOGIC;
  SIGNAL or_1689_nl : STD_LOGIC;
  SIGNAL mux_1811_nl : STD_LOGIC;
  SIGNAL mux_1810_nl : STD_LOGIC;
  SIGNAL or_1680_nl : STD_LOGIC;
  SIGNAL mux_1809_nl : STD_LOGIC;
  SIGNAL mux_1805_nl : STD_LOGIC;
  SIGNAL mux_1804_nl : STD_LOGIC;
  SIGNAL mux_1803_nl : STD_LOGIC;
  SIGNAL mux_1802_nl : STD_LOGIC;
  SIGNAL or_1670_nl : STD_LOGIC;
  SIGNAL mux_1801_nl : STD_LOGIC;
  SIGNAL mux_1799_nl : STD_LOGIC;
  SIGNAL mux_1798_nl : STD_LOGIC;
  SIGNAL mux_1797_nl : STD_LOGIC;
  SIGNAL mux_1796_nl : STD_LOGIC;
  SIGNAL or_1667_nl : STD_LOGIC;
  SIGNAL mux_1795_nl : STD_LOGIC;
  SIGNAL mux_1794_nl : STD_LOGIC;
  SIGNAL or_1662_nl : STD_LOGIC;
  SIGNAL mux_1792_nl : STD_LOGIC;
  SIGNAL mux_1791_nl : STD_LOGIC;
  SIGNAL mux_1790_nl : STD_LOGIC;
  SIGNAL or_1659_nl : STD_LOGIC;
  SIGNAL mux_1789_nl : STD_LOGIC;
  SIGNAL or_1657_nl : STD_LOGIC;
  SIGNAL or_1653_nl : STD_LOGIC;
  SIGNAL mux_1784_nl : STD_LOGIC;
  SIGNAL mux_1783_nl : STD_LOGIC;
  SIGNAL or_1646_nl : STD_LOGIC;
  SIGNAL or_1645_nl : STD_LOGIC;
  SIGNAL mux_1780_nl : STD_LOGIC;
  SIGNAL mux_1779_nl : STD_LOGIC;
  SIGNAL mux_1778_nl : STD_LOGIC;
  SIGNAL or_1638_nl : STD_LOGIC;
  SIGNAL or_1635_nl : STD_LOGIC;
  SIGNAL or_1634_nl : STD_LOGIC;
  SIGNAL mux_1848_nl : STD_LOGIC;
  SIGNAL mux_1847_nl : STD_LOGIC;
  SIGNAL and_621_nl : STD_LOGIC;
  SIGNAL mux_1846_nl : STD_LOGIC;
  SIGNAL nor_899_nl : STD_LOGIC;
  SIGNAL mux_1845_nl : STD_LOGIC;
  SIGNAL nor_901_nl : STD_LOGIC;
  SIGNAL mux_1844_nl : STD_LOGIC;
  SIGNAL nor_902_nl : STD_LOGIC;
  SIGNAL mux_1843_nl : STD_LOGIC;
  SIGNAL or_1735_nl : STD_LOGIC;
  SIGNAL or_1734_nl : STD_LOGIC;
  SIGNAL mux_1842_nl : STD_LOGIC;
  SIGNAL nor_903_nl : STD_LOGIC;
  SIGNAL nor_904_nl : STD_LOGIC;
  SIGNAL mux_1841_nl : STD_LOGIC;
  SIGNAL mux_1840_nl : STD_LOGIC;
  SIGNAL nor_905_nl : STD_LOGIC;
  SIGNAL mux_1839_nl : STD_LOGIC;
  SIGNAL nor_906_nl : STD_LOGIC;
  SIGNAL mux_1838_nl : STD_LOGIC;
  SIGNAL or_1726_nl : STD_LOGIC;
  SIGNAL or_1724_nl : STD_LOGIC;
  SIGNAL nor_907_nl : STD_LOGIC;
  SIGNAL mux_1837_nl : STD_LOGIC;
  SIGNAL nor_908_nl : STD_LOGIC;
  SIGNAL and_622_nl : STD_LOGIC;
  SIGNAL mux_1836_nl : STD_LOGIC;
  SIGNAL nor_909_nl : STD_LOGIC;
  SIGNAL mux_1835_nl : STD_LOGIC;
  SIGNAL nor_910_nl : STD_LOGIC;
  SIGNAL mux_1834_nl : STD_LOGIC;
  SIGNAL mux_1833_nl : STD_LOGIC;
  SIGNAL nor_912_nl : STD_LOGIC;
  SIGNAL mux_1832_nl : STD_LOGIC;
  SIGNAL mux_1831_nl : STD_LOGIC;
  SIGNAL or_1715_nl : STD_LOGIC;
  SIGNAL or_1714_nl : STD_LOGIC;
  SIGNAL mux_1830_nl : STD_LOGIC;
  SIGNAL or_1713_nl : STD_LOGIC;
  SIGNAL or_1711_nl : STD_LOGIC;
  SIGNAL mux_1829_nl : STD_LOGIC;
  SIGNAL mux_1828_nl : STD_LOGIC;
  SIGNAL nor_913_nl : STD_LOGIC;
  SIGNAL nor_914_nl : STD_LOGIC;
  SIGNAL mux_1827_nl : STD_LOGIC;
  SIGNAL or_1706_nl : STD_LOGIC;
  SIGNAL mux_1826_nl : STD_LOGIC;
  SIGNAL nor_915_nl : STD_LOGIC;
  SIGNAL nor_916_nl : STD_LOGIC;
  SIGNAL mux_1825_nl : STD_LOGIC;
  SIGNAL nor_917_nl : STD_LOGIC;
  SIGNAL mux_1824_nl : STD_LOGIC;
  SIGNAL mux_1823_nl : STD_LOGIC;
  SIGNAL or_1700_nl : STD_LOGIC;
  SIGNAL mux_1822_nl : STD_LOGIC;
  SIGNAL or_1698_nl : STD_LOGIC;
  SIGNAL or_1695_nl : STD_LOGIC;
  SIGNAL mux_1821_nl : STD_LOGIC;
  SIGNAL and_623_nl : STD_LOGIC;
  SIGNAL mux_1820_nl : STD_LOGIC;
  SIGNAL nor_918_nl : STD_LOGIC;
  SIGNAL mux_1819_nl : STD_LOGIC;
  SIGNAL nor_919_nl : STD_LOGIC;
  SIGNAL nor_920_nl : STD_LOGIC;
  SIGNAL nor_921_nl : STD_LOGIC;
  SIGNAL mux_1890_nl : STD_LOGIC;
  SIGNAL mux_1889_nl : STD_LOGIC;
  SIGNAL mux_1888_nl : STD_LOGIC;
  SIGNAL mux_1887_nl : STD_LOGIC;
  SIGNAL or_1795_nl : STD_LOGIC;
  SIGNAL mux_1886_nl : STD_LOGIC;
  SIGNAL or_1793_nl : STD_LOGIC;
  SIGNAL or_1792_nl : STD_LOGIC;
  SIGNAL mux_1885_nl : STD_LOGIC;
  SIGNAL mux_1884_nl : STD_LOGIC;
  SIGNAL nand_319_nl : STD_LOGIC;
  SIGNAL or_1790_nl : STD_LOGIC;
  SIGNAL mux_1883_nl : STD_LOGIC;
  SIGNAL mux_1882_nl : STD_LOGIC;
  SIGNAL mux_1881_nl : STD_LOGIC;
  SIGNAL or_1789_nl : STD_LOGIC;
  SIGNAL or_1788_nl : STD_LOGIC;
  SIGNAL mux_1880_nl : STD_LOGIC;
  SIGNAL mux_1879_nl : STD_LOGIC;
  SIGNAL mux_1878_nl : STD_LOGIC;
  SIGNAL mux_1877_nl : STD_LOGIC;
  SIGNAL mux_1876_nl : STD_LOGIC;
  SIGNAL or_1787_nl : STD_LOGIC;
  SIGNAL mux_1874_nl : STD_LOGIC;
  SIGNAL mux_1873_nl : STD_LOGIC;
  SIGNAL or_1778_nl : STD_LOGIC;
  SIGNAL mux_1871_nl : STD_LOGIC;
  SIGNAL mux_1864_nl : STD_LOGIC;
  SIGNAL mux_1863_nl : STD_LOGIC;
  SIGNAL mux_1862_nl : STD_LOGIC;
  SIGNAL mux_1861_nl : STD_LOGIC;
  SIGNAL nand_321_nl : STD_LOGIC;
  SIGNAL mux_1860_nl : STD_LOGIC;
  SIGNAL mux_1856_nl : STD_LOGIC;
  SIGNAL mux_1855_nl : STD_LOGIC;
  SIGNAL mux_1854_nl : STD_LOGIC;
  SIGNAL mux_1853_nl : STD_LOGIC;
  SIGNAL or_1750_nl : STD_LOGIC;
  SIGNAL mux_1852_nl : STD_LOGIC;
  SIGNAL mux_1851_nl : STD_LOGIC;
  SIGNAL or_1743_nl : STD_LOGIC;
  SIGNAL and_620_nl : STD_LOGIC;
  SIGNAL mux_1920_nl : STD_LOGIC;
  SIGNAL mux_1919_nl : STD_LOGIC;
  SIGNAL and_615_nl : STD_LOGIC;
  SIGNAL mux_1918_nl : STD_LOGIC;
  SIGNAL nor_876_nl : STD_LOGIC;
  SIGNAL mux_1917_nl : STD_LOGIC;
  SIGNAL nor_878_nl : STD_LOGIC;
  SIGNAL mux_1916_nl : STD_LOGIC;
  SIGNAL nor_879_nl : STD_LOGIC;
  SIGNAL mux_1915_nl : STD_LOGIC;
  SIGNAL nand_316_nl : STD_LOGIC;
  SIGNAL or_1840_nl : STD_LOGIC;
  SIGNAL mux_1914_nl : STD_LOGIC;
  SIGNAL nor_880_nl : STD_LOGIC;
  SIGNAL nor_881_nl : STD_LOGIC;
  SIGNAL mux_1913_nl : STD_LOGIC;
  SIGNAL mux_1912_nl : STD_LOGIC;
  SIGNAL and_616_nl : STD_LOGIC;
  SIGNAL mux_1911_nl : STD_LOGIC;
  SIGNAL nor_882_nl : STD_LOGIC;
  SIGNAL mux_1910_nl : STD_LOGIC;
  SIGNAL or_1832_nl : STD_LOGIC;
  SIGNAL or_1830_nl : STD_LOGIC;
  SIGNAL nor_883_nl : STD_LOGIC;
  SIGNAL mux_1909_nl : STD_LOGIC;
  SIGNAL nor_884_nl : STD_LOGIC;
  SIGNAL and_617_nl : STD_LOGIC;
  SIGNAL mux_1908_nl : STD_LOGIC;
  SIGNAL and_827_nl : STD_LOGIC;
  SIGNAL mux_1907_nl : STD_LOGIC;
  SIGNAL nor_886_nl : STD_LOGIC;
  SIGNAL mux_1906_nl : STD_LOGIC;
  SIGNAL mux_1905_nl : STD_LOGIC;
  SIGNAL nor_888_nl : STD_LOGIC;
  SIGNAL mux_1904_nl : STD_LOGIC;
  SIGNAL mux_1903_nl : STD_LOGIC;
  SIGNAL or_1821_nl : STD_LOGIC;
  SIGNAL or_1820_nl : STD_LOGIC;
  SIGNAL mux_1902_nl : STD_LOGIC;
  SIGNAL or_1819_nl : STD_LOGIC;
  SIGNAL or_1817_nl : STD_LOGIC;
  SIGNAL mux_1901_nl : STD_LOGIC;
  SIGNAL mux_1900_nl : STD_LOGIC;
  SIGNAL nor_889_nl : STD_LOGIC;
  SIGNAL nor_890_nl : STD_LOGIC;
  SIGNAL mux_1899_nl : STD_LOGIC;
  SIGNAL or_1812_nl : STD_LOGIC;
  SIGNAL mux_1898_nl : STD_LOGIC;
  SIGNAL nor_891_nl : STD_LOGIC;
  SIGNAL nor_892_nl : STD_LOGIC;
  SIGNAL mux_1897_nl : STD_LOGIC;
  SIGNAL nor_893_nl : STD_LOGIC;
  SIGNAL mux_1896_nl : STD_LOGIC;
  SIGNAL mux_1895_nl : STD_LOGIC;
  SIGNAL nand_415_nl : STD_LOGIC;
  SIGNAL mux_1894_nl : STD_LOGIC;
  SIGNAL or_1804_nl : STD_LOGIC;
  SIGNAL or_1801_nl : STD_LOGIC;
  SIGNAL mux_1893_nl : STD_LOGIC;
  SIGNAL and_618_nl : STD_LOGIC;
  SIGNAL mux_1892_nl : STD_LOGIC;
  SIGNAL nor_894_nl : STD_LOGIC;
  SIGNAL mux_1891_nl : STD_LOGIC;
  SIGNAL and_619_nl : STD_LOGIC;
  SIGNAL nor_895_nl : STD_LOGIC;
  SIGNAL nor_896_nl : STD_LOGIC;
  SIGNAL mux_1963_nl : STD_LOGIC;
  SIGNAL mux_1962_nl : STD_LOGIC;
  SIGNAL mux_1961_nl : STD_LOGIC;
  SIGNAL mux_1960_nl : STD_LOGIC;
  SIGNAL mux_1959_nl : STD_LOGIC;
  SIGNAL mux_1958_nl : STD_LOGIC;
  SIGNAL or_1905_nl : STD_LOGIC;
  SIGNAL or_1903_nl : STD_LOGIC;
  SIGNAL or_1902_nl : STD_LOGIC;
  SIGNAL mux_1957_nl : STD_LOGIC;
  SIGNAL nand_311_nl : STD_LOGIC;
  SIGNAL or_1900_nl : STD_LOGIC;
  SIGNAL mux_1956_nl : STD_LOGIC;
  SIGNAL mux_1955_nl : STD_LOGIC;
  SIGNAL mux_1954_nl : STD_LOGIC;
  SIGNAL or_1898_nl : STD_LOGIC;
  SIGNAL or_1896_nl : STD_LOGIC;
  SIGNAL mux_1953_nl : STD_LOGIC;
  SIGNAL or_1894_nl : STD_LOGIC;
  SIGNAL mux_1952_nl : STD_LOGIC;
  SIGNAL nand_437_nl : STD_LOGIC;
  SIGNAL mux_1951_nl : STD_LOGIC;
  SIGNAL or_1891_nl : STD_LOGIC;
  SIGNAL mux_1950_nl : STD_LOGIC;
  SIGNAL mux_1949_nl : STD_LOGIC;
  SIGNAL or_1890_nl : STD_LOGIC;
  SIGNAL mux_1948_nl : STD_LOGIC;
  SIGNAL or_1889_nl : STD_LOGIC;
  SIGNAL or_1888_nl : STD_LOGIC;
  SIGNAL mux_1947_nl : STD_LOGIC;
  SIGNAL mux_1946_nl : STD_LOGIC;
  SIGNAL mux_1945_nl : STD_LOGIC;
  SIGNAL mux_1944_nl : STD_LOGIC;
  SIGNAL or_1887_nl : STD_LOGIC;
  SIGNAL or_1886_nl : STD_LOGIC;
  SIGNAL mux_1943_nl : STD_LOGIC;
  SIGNAL or_1884_nl : STD_LOGIC;
  SIGNAL or_1883_nl : STD_LOGIC;
  SIGNAL mux_1942_nl : STD_LOGIC;
  SIGNAL mux_1941_nl : STD_LOGIC;
  SIGNAL mux_1940_nl : STD_LOGIC;
  SIGNAL or_1882_nl : STD_LOGIC;
  SIGNAL or_1881_nl : STD_LOGIC;
  SIGNAL mux_1939_nl : STD_LOGIC;
  SIGNAL mux_1938_nl : STD_LOGIC;
  SIGNAL mux_1937_nl : STD_LOGIC;
  SIGNAL or_1879_nl : STD_LOGIC;
  SIGNAL or_1876_nl : STD_LOGIC;
  SIGNAL or_1875_nl : STD_LOGIC;
  SIGNAL mux_1936_nl : STD_LOGIC;
  SIGNAL mux_1935_nl : STD_LOGIC;
  SIGNAL mux_1934_nl : STD_LOGIC;
  SIGNAL or_1873_nl : STD_LOGIC;
  SIGNAL mux_1933_nl : STD_LOGIC;
  SIGNAL mux_1932_nl : STD_LOGIC;
  SIGNAL or_1871_nl : STD_LOGIC;
  SIGNAL mux_1931_nl : STD_LOGIC;
  SIGNAL or_1867_nl : STD_LOGIC;
  SIGNAL mux_1930_nl : STD_LOGIC;
  SIGNAL or_1866_nl : STD_LOGIC;
  SIGNAL mux_1928_nl : STD_LOGIC;
  SIGNAL or_1862_nl : STD_LOGIC;
  SIGNAL mux_1924_nl : STD_LOGIC;
  SIGNAL mux_1923_nl : STD_LOGIC;
  SIGNAL or_1850_nl : STD_LOGIC;
  SIGNAL or_1848_nl : STD_LOGIC;
  SIGNAL or_1847_nl : STD_LOGIC;
  SIGNAL mux_1993_nl : STD_LOGIC;
  SIGNAL mux_1992_nl : STD_LOGIC;
  SIGNAL and_612_nl : STD_LOGIC;
  SIGNAL mux_1991_nl : STD_LOGIC;
  SIGNAL nor_849_nl : STD_LOGIC;
  SIGNAL mux_1990_nl : STD_LOGIC;
  SIGNAL nor_851_nl : STD_LOGIC;
  SIGNAL mux_1989_nl : STD_LOGIC;
  SIGNAL nor_852_nl : STD_LOGIC;
  SIGNAL mux_1988_nl : STD_LOGIC;
  SIGNAL or_1951_nl : STD_LOGIC;
  SIGNAL or_1950_nl : STD_LOGIC;
  SIGNAL mux_1987_nl : STD_LOGIC;
  SIGNAL nor_853_nl : STD_LOGIC;
  SIGNAL nor_854_nl : STD_LOGIC;
  SIGNAL mux_1986_nl : STD_LOGIC;
  SIGNAL mux_1985_nl : STD_LOGIC;
  SIGNAL nor_855_nl : STD_LOGIC;
  SIGNAL mux_1984_nl : STD_LOGIC;
  SIGNAL nor_856_nl : STD_LOGIC;
  SIGNAL mux_1983_nl : STD_LOGIC;
  SIGNAL or_1942_nl : STD_LOGIC;
  SIGNAL or_1940_nl : STD_LOGIC;
  SIGNAL nor_857_nl : STD_LOGIC;
  SIGNAL mux_1982_nl : STD_LOGIC;
  SIGNAL nor_858_nl : STD_LOGIC;
  SIGNAL and_613_nl : STD_LOGIC;
  SIGNAL mux_1981_nl : STD_LOGIC;
  SIGNAL nor_859_nl : STD_LOGIC;
  SIGNAL mux_1980_nl : STD_LOGIC;
  SIGNAL nor_860_nl : STD_LOGIC;
  SIGNAL mux_1979_nl : STD_LOGIC;
  SIGNAL mux_1978_nl : STD_LOGIC;
  SIGNAL nor_862_nl : STD_LOGIC;
  SIGNAL mux_1977_nl : STD_LOGIC;
  SIGNAL mux_1976_nl : STD_LOGIC;
  SIGNAL or_1931_nl : STD_LOGIC;
  SIGNAL or_1930_nl : STD_LOGIC;
  SIGNAL mux_1975_nl : STD_LOGIC;
  SIGNAL or_1929_nl : STD_LOGIC;
  SIGNAL or_1927_nl : STD_LOGIC;
  SIGNAL mux_1974_nl : STD_LOGIC;
  SIGNAL mux_1973_nl : STD_LOGIC;
  SIGNAL nor_863_nl : STD_LOGIC;
  SIGNAL nor_864_nl : STD_LOGIC;
  SIGNAL mux_1972_nl : STD_LOGIC;
  SIGNAL or_1922_nl : STD_LOGIC;
  SIGNAL mux_1971_nl : STD_LOGIC;
  SIGNAL nor_865_nl : STD_LOGIC;
  SIGNAL nor_866_nl : STD_LOGIC;
  SIGNAL mux_1970_nl : STD_LOGIC;
  SIGNAL nor_867_nl : STD_LOGIC;
  SIGNAL mux_1969_nl : STD_LOGIC;
  SIGNAL mux_1968_nl : STD_LOGIC;
  SIGNAL or_1916_nl : STD_LOGIC;
  SIGNAL mux_1967_nl : STD_LOGIC;
  SIGNAL or_1914_nl : STD_LOGIC;
  SIGNAL or_1911_nl : STD_LOGIC;
  SIGNAL mux_1966_nl : STD_LOGIC;
  SIGNAL and_614_nl : STD_LOGIC;
  SIGNAL mux_1965_nl : STD_LOGIC;
  SIGNAL nor_868_nl : STD_LOGIC;
  SIGNAL mux_1964_nl : STD_LOGIC;
  SIGNAL nor_869_nl : STD_LOGIC;
  SIGNAL nor_870_nl : STD_LOGIC;
  SIGNAL nor_871_nl : STD_LOGIC;
  SIGNAL mux_2035_nl : STD_LOGIC;
  SIGNAL mux_2034_nl : STD_LOGIC;
  SIGNAL mux_2033_nl : STD_LOGIC;
  SIGNAL mux_2032_nl : STD_LOGIC;
  SIGNAL or_2011_nl : STD_LOGIC;
  SIGNAL mux_2031_nl : STD_LOGIC;
  SIGNAL or_2009_nl : STD_LOGIC;
  SIGNAL or_2008_nl : STD_LOGIC;
  SIGNAL mux_2030_nl : STD_LOGIC;
  SIGNAL mux_2029_nl : STD_LOGIC;
  SIGNAL nand_305_nl : STD_LOGIC;
  SIGNAL or_2006_nl : STD_LOGIC;
  SIGNAL mux_2028_nl : STD_LOGIC;
  SIGNAL mux_2027_nl : STD_LOGIC;
  SIGNAL mux_2026_nl : STD_LOGIC;
  SIGNAL or_2005_nl : STD_LOGIC;
  SIGNAL or_2004_nl : STD_LOGIC;
  SIGNAL mux_2025_nl : STD_LOGIC;
  SIGNAL mux_2024_nl : STD_LOGIC;
  SIGNAL mux_2023_nl : STD_LOGIC;
  SIGNAL mux_2022_nl : STD_LOGIC;
  SIGNAL mux_2021_nl : STD_LOGIC;
  SIGNAL or_2003_nl : STD_LOGIC;
  SIGNAL mux_2019_nl : STD_LOGIC;
  SIGNAL mux_2018_nl : STD_LOGIC;
  SIGNAL or_1994_nl : STD_LOGIC;
  SIGNAL mux_2016_nl : STD_LOGIC;
  SIGNAL mux_2009_nl : STD_LOGIC;
  SIGNAL mux_2008_nl : STD_LOGIC;
  SIGNAL mux_2007_nl : STD_LOGIC;
  SIGNAL mux_2006_nl : STD_LOGIC;
  SIGNAL nand_307_nl : STD_LOGIC;
  SIGNAL mux_2005_nl : STD_LOGIC;
  SIGNAL mux_2001_nl : STD_LOGIC;
  SIGNAL mux_2000_nl : STD_LOGIC;
  SIGNAL mux_1999_nl : STD_LOGIC;
  SIGNAL mux_1998_nl : STD_LOGIC;
  SIGNAL or_1966_nl : STD_LOGIC;
  SIGNAL mux_1997_nl : STD_LOGIC;
  SIGNAL mux_1996_nl : STD_LOGIC;
  SIGNAL or_1959_nl : STD_LOGIC;
  SIGNAL and_611_nl : STD_LOGIC;
  SIGNAL mux_2065_nl : STD_LOGIC;
  SIGNAL mux_2064_nl : STD_LOGIC;
  SIGNAL and_606_nl : STD_LOGIC;
  SIGNAL mux_2063_nl : STD_LOGIC;
  SIGNAL nor_826_nl : STD_LOGIC;
  SIGNAL mux_2062_nl : STD_LOGIC;
  SIGNAL nor_828_nl : STD_LOGIC;
  SIGNAL mux_2061_nl : STD_LOGIC;
  SIGNAL nor_829_nl : STD_LOGIC;
  SIGNAL mux_2060_nl : STD_LOGIC;
  SIGNAL nand_302_nl : STD_LOGIC;
  SIGNAL or_2056_nl : STD_LOGIC;
  SIGNAL mux_2059_nl : STD_LOGIC;
  SIGNAL nor_830_nl : STD_LOGIC;
  SIGNAL nor_831_nl : STD_LOGIC;
  SIGNAL mux_2058_nl : STD_LOGIC;
  SIGNAL mux_2057_nl : STD_LOGIC;
  SIGNAL and_607_nl : STD_LOGIC;
  SIGNAL mux_2056_nl : STD_LOGIC;
  SIGNAL nor_832_nl : STD_LOGIC;
  SIGNAL mux_2055_nl : STD_LOGIC;
  SIGNAL or_2048_nl : STD_LOGIC;
  SIGNAL or_2046_nl : STD_LOGIC;
  SIGNAL nor_833_nl : STD_LOGIC;
  SIGNAL mux_2054_nl : STD_LOGIC;
  SIGNAL nor_834_nl : STD_LOGIC;
  SIGNAL and_608_nl : STD_LOGIC;
  SIGNAL mux_2053_nl : STD_LOGIC;
  SIGNAL and_826_nl : STD_LOGIC;
  SIGNAL mux_2052_nl : STD_LOGIC;
  SIGNAL nor_836_nl : STD_LOGIC;
  SIGNAL mux_2051_nl : STD_LOGIC;
  SIGNAL mux_2050_nl : STD_LOGIC;
  SIGNAL nor_838_nl : STD_LOGIC;
  SIGNAL mux_2049_nl : STD_LOGIC;
  SIGNAL mux_2048_nl : STD_LOGIC;
  SIGNAL or_2037_nl : STD_LOGIC;
  SIGNAL or_2036_nl : STD_LOGIC;
  SIGNAL mux_2047_nl : STD_LOGIC;
  SIGNAL or_2035_nl : STD_LOGIC;
  SIGNAL or_2033_nl : STD_LOGIC;
  SIGNAL mux_2046_nl : STD_LOGIC;
  SIGNAL mux_2045_nl : STD_LOGIC;
  SIGNAL nor_839_nl : STD_LOGIC;
  SIGNAL nor_840_nl : STD_LOGIC;
  SIGNAL mux_2044_nl : STD_LOGIC;
  SIGNAL or_2028_nl : STD_LOGIC;
  SIGNAL mux_2043_nl : STD_LOGIC;
  SIGNAL nor_841_nl : STD_LOGIC;
  SIGNAL nor_842_nl : STD_LOGIC;
  SIGNAL mux_2042_nl : STD_LOGIC;
  SIGNAL nor_843_nl : STD_LOGIC;
  SIGNAL mux_2041_nl : STD_LOGIC;
  SIGNAL mux_2040_nl : STD_LOGIC;
  SIGNAL nand_413_nl : STD_LOGIC;
  SIGNAL mux_2039_nl : STD_LOGIC;
  SIGNAL or_2020_nl : STD_LOGIC;
  SIGNAL or_2017_nl : STD_LOGIC;
  SIGNAL mux_2038_nl : STD_LOGIC;
  SIGNAL and_609_nl : STD_LOGIC;
  SIGNAL mux_2037_nl : STD_LOGIC;
  SIGNAL nor_844_nl : STD_LOGIC;
  SIGNAL mux_2036_nl : STD_LOGIC;
  SIGNAL and_610_nl : STD_LOGIC;
  SIGNAL nor_845_nl : STD_LOGIC;
  SIGNAL nor_846_nl : STD_LOGIC;
  SIGNAL mux_2107_nl : STD_LOGIC;
  SIGNAL mux_2106_nl : STD_LOGIC;
  SIGNAL mux_2105_nl : STD_LOGIC;
  SIGNAL mux_2104_nl : STD_LOGIC;
  SIGNAL mux_2103_nl : STD_LOGIC;
  SIGNAL mux_2102_nl : STD_LOGIC;
  SIGNAL or_2118_nl : STD_LOGIC;
  SIGNAL mux_2100_nl : STD_LOGIC;
  SIGNAL mux_2099_nl : STD_LOGIC;
  SIGNAL or_2109_nl : STD_LOGIC;
  SIGNAL mux_2098_nl : STD_LOGIC;
  SIGNAL mux_2094_nl : STD_LOGIC;
  SIGNAL mux_2093_nl : STD_LOGIC;
  SIGNAL mux_2092_nl : STD_LOGIC;
  SIGNAL mux_2091_nl : STD_LOGIC;
  SIGNAL nand_297_nl : STD_LOGIC;
  SIGNAL mux_2090_nl : STD_LOGIC;
  SIGNAL mux_2088_nl : STD_LOGIC;
  SIGNAL mux_2087_nl : STD_LOGIC;
  SIGNAL mux_2086_nl : STD_LOGIC;
  SIGNAL mux_2085_nl : STD_LOGIC;
  SIGNAL or_2096_nl : STD_LOGIC;
  SIGNAL mux_2084_nl : STD_LOGIC;
  SIGNAL mux_2083_nl : STD_LOGIC;
  SIGNAL or_2091_nl : STD_LOGIC;
  SIGNAL mux_2081_nl : STD_LOGIC;
  SIGNAL mux_2080_nl : STD_LOGIC;
  SIGNAL mux_2079_nl : STD_LOGIC;
  SIGNAL or_2088_nl : STD_LOGIC;
  SIGNAL mux_2078_nl : STD_LOGIC;
  SIGNAL or_2086_nl : STD_LOGIC;
  SIGNAL or_2082_nl : STD_LOGIC;
  SIGNAL mux_2073_nl : STD_LOGIC;
  SIGNAL mux_2072_nl : STD_LOGIC;
  SIGNAL nand_298_nl : STD_LOGIC;
  SIGNAL or_2074_nl : STD_LOGIC;
  SIGNAL mux_2069_nl : STD_LOGIC;
  SIGNAL mux_2068_nl : STD_LOGIC;
  SIGNAL mux_2067_nl : STD_LOGIC;
  SIGNAL or_2067_nl : STD_LOGIC;
  SIGNAL or_2064_nl : STD_LOGIC;
  SIGNAL nand_299_nl : STD_LOGIC;
  SIGNAL mux_2137_nl : STD_LOGIC;
  SIGNAL mux_2136_nl : STD_LOGIC;
  SIGNAL and_601_nl : STD_LOGIC;
  SIGNAL mux_2135_nl : STD_LOGIC;
  SIGNAL nor_803_nl : STD_LOGIC;
  SIGNAL mux_2134_nl : STD_LOGIC;
  SIGNAL nor_805_nl : STD_LOGIC;
  SIGNAL mux_2133_nl : STD_LOGIC;
  SIGNAL nor_806_nl : STD_LOGIC;
  SIGNAL mux_2132_nl : STD_LOGIC;
  SIGNAL nand_293_nl : STD_LOGIC;
  SIGNAL or_2163_nl : STD_LOGIC;
  SIGNAL mux_2131_nl : STD_LOGIC;
  SIGNAL nor_807_nl : STD_LOGIC;
  SIGNAL nor_808_nl : STD_LOGIC;
  SIGNAL mux_2130_nl : STD_LOGIC;
  SIGNAL mux_2129_nl : STD_LOGIC;
  SIGNAL and_602_nl : STD_LOGIC;
  SIGNAL mux_2128_nl : STD_LOGIC;
  SIGNAL nor_809_nl : STD_LOGIC;
  SIGNAL mux_2127_nl : STD_LOGIC;
  SIGNAL or_2155_nl : STD_LOGIC;
  SIGNAL or_2153_nl : STD_LOGIC;
  SIGNAL nor_810_nl : STD_LOGIC;
  SIGNAL mux_2126_nl : STD_LOGIC;
  SIGNAL nor_811_nl : STD_LOGIC;
  SIGNAL and_603_nl : STD_LOGIC;
  SIGNAL mux_2125_nl : STD_LOGIC;
  SIGNAL and_825_nl : STD_LOGIC;
  SIGNAL mux_2124_nl : STD_LOGIC;
  SIGNAL nor_813_nl : STD_LOGIC;
  SIGNAL mux_2123_nl : STD_LOGIC;
  SIGNAL mux_2122_nl : STD_LOGIC;
  SIGNAL nor_815_nl : STD_LOGIC;
  SIGNAL mux_2121_nl : STD_LOGIC;
  SIGNAL mux_2120_nl : STD_LOGIC;
  SIGNAL or_2144_nl : STD_LOGIC;
  SIGNAL or_2143_nl : STD_LOGIC;
  SIGNAL mux_2119_nl : STD_LOGIC;
  SIGNAL or_2142_nl : STD_LOGIC;
  SIGNAL or_2140_nl : STD_LOGIC;
  SIGNAL mux_2118_nl : STD_LOGIC;
  SIGNAL mux_2117_nl : STD_LOGIC;
  SIGNAL nor_816_nl : STD_LOGIC;
  SIGNAL nor_817_nl : STD_LOGIC;
  SIGNAL mux_2116_nl : STD_LOGIC;
  SIGNAL or_2135_nl : STD_LOGIC;
  SIGNAL mux_2115_nl : STD_LOGIC;
  SIGNAL nor_818_nl : STD_LOGIC;
  SIGNAL nor_819_nl : STD_LOGIC;
  SIGNAL mux_2114_nl : STD_LOGIC;
  SIGNAL nor_820_nl : STD_LOGIC;
  SIGNAL mux_2113_nl : STD_LOGIC;
  SIGNAL mux_2112_nl : STD_LOGIC;
  SIGNAL nand_411_nl : STD_LOGIC;
  SIGNAL mux_2111_nl : STD_LOGIC;
  SIGNAL or_2127_nl : STD_LOGIC;
  SIGNAL or_2124_nl : STD_LOGIC;
  SIGNAL mux_2110_nl : STD_LOGIC;
  SIGNAL and_604_nl : STD_LOGIC;
  SIGNAL mux_2109_nl : STD_LOGIC;
  SIGNAL nor_821_nl : STD_LOGIC;
  SIGNAL mux_2108_nl : STD_LOGIC;
  SIGNAL and_605_nl : STD_LOGIC;
  SIGNAL nor_822_nl : STD_LOGIC;
  SIGNAL nor_823_nl : STD_LOGIC;
  SIGNAL mux_2179_nl : STD_LOGIC;
  SIGNAL mux_2178_nl : STD_LOGIC;
  SIGNAL mux_2177_nl : STD_LOGIC;
  SIGNAL mux_2176_nl : STD_LOGIC;
  SIGNAL or_2224_nl : STD_LOGIC;
  SIGNAL mux_2175_nl : STD_LOGIC;
  SIGNAL or_2222_nl : STD_LOGIC;
  SIGNAL or_2221_nl : STD_LOGIC;
  SIGNAL mux_2174_nl : STD_LOGIC;
  SIGNAL mux_2173_nl : STD_LOGIC;
  SIGNAL nand_284_nl : STD_LOGIC;
  SIGNAL or_2219_nl : STD_LOGIC;
  SIGNAL mux_2172_nl : STD_LOGIC;
  SIGNAL mux_2171_nl : STD_LOGIC;
  SIGNAL mux_2170_nl : STD_LOGIC;
  SIGNAL or_2218_nl : STD_LOGIC;
  SIGNAL or_2217_nl : STD_LOGIC;
  SIGNAL mux_2169_nl : STD_LOGIC;
  SIGNAL mux_2168_nl : STD_LOGIC;
  SIGNAL mux_2167_nl : STD_LOGIC;
  SIGNAL mux_2166_nl : STD_LOGIC;
  SIGNAL mux_2165_nl : STD_LOGIC;
  SIGNAL nand_438_nl : STD_LOGIC;
  SIGNAL mux_2163_nl : STD_LOGIC;
  SIGNAL mux_2162_nl : STD_LOGIC;
  SIGNAL or_2207_nl : STD_LOGIC;
  SIGNAL mux_2160_nl : STD_LOGIC;
  SIGNAL mux_2153_nl : STD_LOGIC;
  SIGNAL mux_2152_nl : STD_LOGIC;
  SIGNAL mux_2151_nl : STD_LOGIC;
  SIGNAL mux_2150_nl : STD_LOGIC;
  SIGNAL nand_286_nl : STD_LOGIC;
  SIGNAL mux_2149_nl : STD_LOGIC;
  SIGNAL mux_2145_nl : STD_LOGIC;
  SIGNAL mux_2144_nl : STD_LOGIC;
  SIGNAL mux_2143_nl : STD_LOGIC;
  SIGNAL mux_2142_nl : STD_LOGIC;
  SIGNAL or_2179_nl : STD_LOGIC;
  SIGNAL mux_2141_nl : STD_LOGIC;
  SIGNAL mux_2140_nl : STD_LOGIC;
  SIGNAL or_2172_nl : STD_LOGIC;
  SIGNAL and_600_nl : STD_LOGIC;
  SIGNAL mux_2209_nl : STD_LOGIC;
  SIGNAL mux_2208_nl : STD_LOGIC;
  SIGNAL and_590_nl : STD_LOGIC;
  SIGNAL mux_2207_nl : STD_LOGIC;
  SIGNAL and_823_nl : STD_LOGIC;
  SIGNAL mux_2206_nl : STD_LOGIC;
  SIGNAL nor_786_nl : STD_LOGIC;
  SIGNAL mux_2205_nl : STD_LOGIC;
  SIGNAL nor_787_nl : STD_LOGIC;
  SIGNAL mux_2204_nl : STD_LOGIC;
  SIGNAL nand_269_nl : STD_LOGIC;
  SIGNAL or_2269_nl : STD_LOGIC;
  SIGNAL mux_2203_nl : STD_LOGIC;
  SIGNAL nor_788_nl : STD_LOGIC;
  SIGNAL nor_789_nl : STD_LOGIC;
  SIGNAL mux_2202_nl : STD_LOGIC;
  SIGNAL mux_2201_nl : STD_LOGIC;
  SIGNAL and_592_nl : STD_LOGIC;
  SIGNAL mux_2200_nl : STD_LOGIC;
  SIGNAL nor_790_nl : STD_LOGIC;
  SIGNAL mux_2199_nl : STD_LOGIC;
  SIGNAL nand_436_nl : STD_LOGIC;
  SIGNAL nand_434_nl : STD_LOGIC;
  SIGNAL nor_791_nl : STD_LOGIC;
  SIGNAL mux_2198_nl : STD_LOGIC;
  SIGNAL nor_792_nl : STD_LOGIC;
  SIGNAL and_593_nl : STD_LOGIC;
  SIGNAL mux_2197_nl : STD_LOGIC;
  SIGNAL and_824_nl : STD_LOGIC;
  SIGNAL mux_2196_nl : STD_LOGIC;
  SIGNAL and_594_nl : STD_LOGIC;
  SIGNAL mux_2195_nl : STD_LOGIC;
  SIGNAL mux_2194_nl : STD_LOGIC;
  SIGNAL nor_794_nl : STD_LOGIC;
  SIGNAL mux_2193_nl : STD_LOGIC;
  SIGNAL mux_2192_nl : STD_LOGIC;
  SIGNAL nand_274_nl : STD_LOGIC;
  SIGNAL nand_275_nl : STD_LOGIC;
  SIGNAL mux_2191_nl : STD_LOGIC;
  SIGNAL or_2248_nl : STD_LOGIC;
  SIGNAL nand_277_nl : STD_LOGIC;
  SIGNAL mux_2190_nl : STD_LOGIC;
  SIGNAL mux_2189_nl : STD_LOGIC;
  SIGNAL nor_795_nl : STD_LOGIC;
  SIGNAL nor_796_nl : STD_LOGIC;
  SIGNAL mux_2188_nl : STD_LOGIC;
  SIGNAL or_2241_nl : STD_LOGIC;
  SIGNAL mux_2187_nl : STD_LOGIC;
  SIGNAL nor_797_nl : STD_LOGIC;
  SIGNAL and_596_nl : STD_LOGIC;
  SIGNAL mux_2186_nl : STD_LOGIC;
  SIGNAL nor_798_nl : STD_LOGIC;
  SIGNAL mux_2185_nl : STD_LOGIC;
  SIGNAL mux_2184_nl : STD_LOGIC;
  SIGNAL nand_409_nl : STD_LOGIC;
  SIGNAL mux_2183_nl : STD_LOGIC;
  SIGNAL or_2233_nl : STD_LOGIC;
  SIGNAL or_2230_nl : STD_LOGIC;
  SIGNAL mux_2182_nl : STD_LOGIC;
  SIGNAL and_597_nl : STD_LOGIC;
  SIGNAL mux_2181_nl : STD_LOGIC;
  SIGNAL and_598_nl : STD_LOGIC;
  SIGNAL mux_2180_nl : STD_LOGIC;
  SIGNAL and_599_nl : STD_LOGIC;
  SIGNAL nor_799_nl : STD_LOGIC;
  SIGNAL nor_800_nl : STD_LOGIC;
  SIGNAL nand_450_nl : STD_LOGIC;
  SIGNAL or_3357_nl : STD_LOGIC;
  SIGNAL mux_3723_nl : STD_LOGIC;
  SIGNAL mux_3722_nl : STD_LOGIC;
  SIGNAL mux_3721_nl : STD_LOGIC;
  SIGNAL nand_439_nl : STD_LOGIC;
  SIGNAL or_3373_nl : STD_LOGIC;
  SIGNAL mux_3720_nl : STD_LOGIC;
  SIGNAL or_3371_nl : STD_LOGIC;
  SIGNAL or_3369_nl : STD_LOGIC;
  SIGNAL or_3368_nl : STD_LOGIC;
  SIGNAL mux_3719_nl : STD_LOGIC;
  SIGNAL mux_3718_nl : STD_LOGIC;
  SIGNAL or_3367_nl : STD_LOGIC;
  SIGNAL or_3366_nl : STD_LOGIC;
  SIGNAL or_3365_nl : STD_LOGIC;
  SIGNAL mux_3717_nl : STD_LOGIC;
  SIGNAL nand_445_nl : STD_LOGIC;
  SIGNAL mux_3716_nl : STD_LOGIC;
  SIGNAL mux_3715_nl : STD_LOGIC;
  SIGNAL nor_1381_nl : STD_LOGIC;
  SIGNAL nor_1382_nl : STD_LOGIC;
  SIGNAL nor_1383_nl : STD_LOGIC;
  SIGNAL mux_3714_nl : STD_LOGIC;
  SIGNAL or_3358_nl : STD_LOGIC;
  SIGNAL mux_3713_nl : STD_LOGIC;
  SIGNAL mux_3712_nl : STD_LOGIC;
  SIGNAL or_3356_nl : STD_LOGIC;
  SIGNAL or_3355_nl : STD_LOGIC;
  SIGNAL nand_455_nl : STD_LOGIC;
  SIGNAL or_3396_nl : STD_LOGIC;
  SIGNAL or_3406_nl : STD_LOGIC;
  SIGNAL or_3409_nl : STD_LOGIC;
  SIGNAL mux_3771_nl : STD_LOGIC;
  SIGNAL or_3413_nl : STD_LOGIC;
  SIGNAL mux_3787_nl : STD_LOGIC;
  SIGNAL mux_3786_nl : STD_LOGIC;
  SIGNAL mux_3785_nl : STD_LOGIC;
  SIGNAL mux_3784_nl : STD_LOGIC;
  SIGNAL mux_3783_nl : STD_LOGIC;
  SIGNAL or_3420_nl : STD_LOGIC;
  SIGNAL mux_3782_nl : STD_LOGIC;
  SIGNAL or_3418_nl : STD_LOGIC;
  SIGNAL mux_3781_nl : STD_LOGIC;
  SIGNAL mux_3780_nl : STD_LOGIC;
  SIGNAL mux_3779_nl : STD_LOGIC;
  SIGNAL mux_3778_nl : STD_LOGIC;
  SIGNAL mux_3777_nl : STD_LOGIC;
  SIGNAL or_3417_nl : STD_LOGIC;
  SIGNAL mux_3776_nl : STD_LOGIC;
  SIGNAL or_3415_nl : STD_LOGIC;
  SIGNAL mux_3775_nl : STD_LOGIC;
  SIGNAL mux_3774_nl : STD_LOGIC;
  SIGNAL mux_3773_nl : STD_LOGIC;
  SIGNAL mux_3770_nl : STD_LOGIC;
  SIGNAL mux_3769_nl : STD_LOGIC;
  SIGNAL mux_3768_nl : STD_LOGIC;
  SIGNAL or_3411_nl : STD_LOGIC;
  SIGNAL mux_3767_nl : STD_LOGIC;
  SIGNAL mux_3766_nl : STD_LOGIC;
  SIGNAL mux_3765_nl : STD_LOGIC;
  SIGNAL mux_3764_nl : STD_LOGIC;
  SIGNAL mux_3762_nl : STD_LOGIC;
  SIGNAL mux_3761_nl : STD_LOGIC;
  SIGNAL mux_3760_nl : STD_LOGIC;
  SIGNAL or_3407_nl : STD_LOGIC;
  SIGNAL mux_3759_nl : STD_LOGIC;
  SIGNAL mux_3758_nl : STD_LOGIC;
  SIGNAL mux_3757_nl : STD_LOGIC;
  SIGNAL mux_3756_nl : STD_LOGIC;
  SIGNAL mux_3755_nl : STD_LOGIC;
  SIGNAL mux_3753_nl : STD_LOGIC;
  SIGNAL mux_3751_nl : STD_LOGIC;
  SIGNAL or_3403_nl : STD_LOGIC;
  SIGNAL mux_3750_nl : STD_LOGIC;
  SIGNAL mux_3749_nl : STD_LOGIC;
  SIGNAL mux_3748_nl : STD_LOGIC;
  SIGNAL or_3401_nl : STD_LOGIC;
  SIGNAL mux_3747_nl : STD_LOGIC;
  SIGNAL mux_3746_nl : STD_LOGIC;
  SIGNAL mux_3745_nl : STD_LOGIC;
  SIGNAL mux_3742_nl : STD_LOGIC;
  SIGNAL mux_3741_nl : STD_LOGIC;
  SIGNAL mux_3740_nl : STD_LOGIC;
  SIGNAL or_3395_nl : STD_LOGIC;
  SIGNAL mux_3739_nl : STD_LOGIC;
  SIGNAL or_3392_nl : STD_LOGIC;
  SIGNAL mux_3737_nl : STD_LOGIC;
  SIGNAL mux_3735_nl : STD_LOGIC;
  SIGNAL mux_3733_nl : STD_LOGIC;
  SIGNAL mux_3732_nl : STD_LOGIC;
  SIGNAL mux_3731_nl : STD_LOGIC;
  SIGNAL mux_3730_nl : STD_LOGIC;
  SIGNAL or_3384_nl : STD_LOGIC;
  SIGNAL mux_3728_nl : STD_LOGIC;
  SIGNAL mux_3727_nl : STD_LOGIC;
  SIGNAL or_3376_nl : STD_LOGIC;
  SIGNAL mux_3801_nl : STD_LOGIC;
  SIGNAL and_1248_nl : STD_LOGIC;
  SIGNAL mux_3800_nl : STD_LOGIC;
  SIGNAL nor_1369_nl : STD_LOGIC;
  SIGNAL and_1249_nl : STD_LOGIC;
  SIGNAL mux_3799_nl : STD_LOGIC;
  SIGNAL nor_1370_nl : STD_LOGIC;
  SIGNAL nor_1371_nl : STD_LOGIC;
  SIGNAL nor_1372_nl : STD_LOGIC;
  SIGNAL mux_3798_nl : STD_LOGIC;
  SIGNAL or_3441_nl : STD_LOGIC;
  SIGNAL mux_3797_nl : STD_LOGIC;
  SIGNAL or_3439_nl : STD_LOGIC;
  SIGNAL or_3438_nl : STD_LOGIC;
  SIGNAL mux_3796_nl : STD_LOGIC;
  SIGNAL mux_3795_nl : STD_LOGIC;
  SIGNAL mux_3794_nl : STD_LOGIC;
  SIGNAL mux_3793_nl : STD_LOGIC;
  SIGNAL nor_1373_nl : STD_LOGIC;
  SIGNAL nor_1374_nl : STD_LOGIC;
  SIGNAL nor_1375_nl : STD_LOGIC;
  SIGNAL nor_1376_nl : STD_LOGIC;
  SIGNAL mux_3792_nl : STD_LOGIC;
  SIGNAL or_3431_nl : STD_LOGIC;
  SIGNAL or_3430_nl : STD_LOGIC;
  SIGNAL mux_3791_nl : STD_LOGIC;
  SIGNAL and_1250_nl : STD_LOGIC;
  SIGNAL mux_3790_nl : STD_LOGIC;
  SIGNAL nor_1378_nl : STD_LOGIC;
  SIGNAL nor_1379_nl : STD_LOGIC;
  SIGNAL mux_3789_nl : STD_LOGIC;
  SIGNAL or_3424_nl : STD_LOGIC;
  SIGNAL or_3422_nl : STD_LOGIC;
  SIGNAL nor_1460_nl : STD_LOGIC;
  SIGNAL and_1267_nl : STD_LOGIC;
  SIGNAL mux_3898_nl : STD_LOGIC;
  SIGNAL or_3516_nl : STD_LOGIC;
  SIGNAL mux_3902_nl : STD_LOGIC;
  SIGNAL nand_470_nl : STD_LOGIC;
  SIGNAL or_3531_nl : STD_LOGIC;
  SIGNAL or_3530_nl : STD_LOGIC;
  SIGNAL mux_3906_nl : STD_LOGIC;
  SIGNAL acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_18_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_or_77_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_19_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_84_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_mux_20_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_20_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_85_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_585_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_1278_nl : STD_LOGIC;
  SIGNAL and_1279_nl : STD_LOGIC;
  SIGNAL and_1280_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_78_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_86_nl : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL and_1281_nl : STD_LOGIC;
  SIGNAL and_1282_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_586_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_1283_nl : STD_LOGIC;
  SIGNAL and_1284_nl : STD_LOGIC;
  SIGNAL and_1285_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_587_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_588_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_64_false_1_mux1h_2_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_64_false_1_or_1_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL operator_64_false_1_mux1h_3_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_104_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_105_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_589_nl : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_or_79_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_285_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_590_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL not_8636_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_591_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_or_80_nl : STD_LOGIC;
  SIGNAL acc_8_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_87_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_592_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_593_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_594_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_595_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_596_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_597_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_81_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_82_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_990_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_23_nl : STD_LOGIC;
  SIGNAL acc_9_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_24_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_598_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_or_83_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_22_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_or_84_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_25_nl : STD_LOGIC;
  SIGNAL modExp_while_if_mux_1_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_3954_nl : STD_LOGIC;
  SIGNAL mux_3955_nl : STD_LOGIC;
  SIGNAL mux_3956_nl : STD_LOGIC;
  SIGNAL mux_3957_nl : STD_LOGIC;
  SIGNAL mux_3958_nl : STD_LOGIC;
  SIGNAL nor_1463_nl : STD_LOGIC;
  SIGNAL nor_1464_nl : STD_LOGIC;
  SIGNAL nor_1465_nl : STD_LOGIC;
  SIGNAL mux_3959_nl : STD_LOGIC;
  SIGNAL nor_1466_nl : STD_LOGIC;
  SIGNAL mux_3960_nl : STD_LOGIC;
  SIGNAL nor_1467_nl : STD_LOGIC;
  SIGNAL nor_1468_nl : STD_LOGIC;
  SIGNAL mux_3961_nl : STD_LOGIC;
  SIGNAL mux_3962_nl : STD_LOGIC;
  SIGNAL nor_1469_nl : STD_LOGIC;
  SIGNAL nor_1470_nl : STD_LOGIC;
  SIGNAL mux_3963_nl : STD_LOGIC;
  SIGNAL nor_1471_nl : STD_LOGIC;
  SIGNAL nor_1472_nl : STD_LOGIC;
  SIGNAL mux_3964_nl : STD_LOGIC;
  SIGNAL or_3612_nl : STD_LOGIC;
  SIGNAL or_3613_nl : STD_LOGIC;
  SIGNAL mux_3965_nl : STD_LOGIC;
  SIGNAL mux_3966_nl : STD_LOGIC;
  SIGNAL and_1286_nl : STD_LOGIC;
  SIGNAL mux_3967_nl : STD_LOGIC;
  SIGNAL nor_1473_nl : STD_LOGIC;
  SIGNAL nor_1474_nl : STD_LOGIC;
  SIGNAL nor_1475_nl : STD_LOGIC;
  SIGNAL mux_3968_nl : STD_LOGIC;
  SIGNAL nor_1476_nl : STD_LOGIC;
  SIGNAL mux_3969_nl : STD_LOGIC;
  SIGNAL and_1287_nl : STD_LOGIC;
  SIGNAL nor_1477_nl : STD_LOGIC;
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL r_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL modulo_result_rem_cmp_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_result_rem_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL operator_66_true_div_cmp_a_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_b : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL STAGE_LOOP_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_rg_z : STD_LOGIC_VECTOR (9 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
      STAGE_LOOP_C_8_tr0 : IN STD_LOGIC;
      modExp_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_1_tr0 : IN STD_LOGIC;
      COMP_LOOP_1_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_62_tr0 : IN STD_LOGIC;
      COMP_LOOP_2_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_124_tr0 : IN STD_LOGIC;
      COMP_LOOP_3_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_186_tr0 : IN STD_LOGIC;
      COMP_LOOP_4_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_248_tr0 : IN STD_LOGIC;
      COMP_LOOP_5_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_310_tr0 : IN STD_LOGIC;
      COMP_LOOP_6_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_372_tr0 : IN STD_LOGIC;
      COMP_LOOP_7_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_434_tr0 : IN STD_LOGIC;
      COMP_LOOP_8_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_496_tr0 : IN STD_LOGIC;
      COMP_LOOP_9_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_558_tr0 : IN STD_LOGIC;
      COMP_LOOP_10_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_620_tr0 : IN STD_LOGIC;
      COMP_LOOP_11_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_682_tr0 : IN STD_LOGIC;
      COMP_LOOP_12_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_744_tr0 : IN STD_LOGIC;
      COMP_LOOP_13_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_806_tr0 : IN STD_LOGIC;
      COMP_LOOP_14_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_868_tr0 : IN STD_LOGIC;
      COMP_LOOP_15_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_930_tr0 : IN STD_LOGIC;
      COMP_LOOP_16_modExp_1_while_C_38_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_992_tr0 : IN STD_LOGIC;
      VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_9_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (10 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_496_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_558_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_620_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_682_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_744_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_806_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_868_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_930_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0 :
      STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_6_2(input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_12_3_2(input_2 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(11 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(11 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_7_2(input_6 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_4_2(input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_17_2(input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(16 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_21_2(input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(20 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_3_2(input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_4_2(input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_6_2(input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_65_3_2(input_2 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(64 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(64 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_4_2(input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_7_7_2(input_6 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_8_19_2(input_18 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(18 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(7 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(7 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_12_2_2(input_0 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(11 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_2_2_2(input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_63_2_2(input_0 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(62 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(62 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_65_2_2(input_0 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(64 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_9_2_2(input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  r_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      dat => r_rsci_dat,
      idat => r_rsci_idat_1
    );
  r_rsci_dat <= r_rsc_dat;
  r_rsci_idat <= r_rsci_idat_1;

  vec_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_15_lz
    );
  vec_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_14_lz
    );
  vec_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_13_lz
    );
  vec_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_12_lz
    );
  vec_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_11_lz
    );
  vec_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_10_lz
    );
  vec_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_9_lz
    );
  vec_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_8_lz
    );
  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_7_lz
    );
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_6_lz
    );
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_5_lz
    );
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_4_lz
    );
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_3_lz
    );
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_2_lz
    );
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_1_lz
    );
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  modulo_result_rem_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 1
      )
    PORT MAP(
      a => modulo_result_rem_cmp_a_1,
      b => modulo_result_rem_cmp_b_1,
      z => modulo_result_rem_cmp_z_1
    );
  modulo_result_rem_cmp_a_1 <= modulo_result_rem_cmp_a;
  modulo_result_rem_cmp_b_1 <= modulo_result_rem_cmp_b;
  modulo_result_rem_cmp_z <= modulo_result_rem_cmp_z_1;

  operator_66_true_div_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 65,
      width_b => 11,
      signd => 1
      )
    PORT MAP(
      a => operator_66_true_div_cmp_a_1,
      b => operator_66_true_div_cmp_b,
      z => operator_66_true_div_cmp_z_1
    );
  operator_66_true_div_cmp_a_1 <= operator_66_true_div_cmp_a;
  operator_66_true_div_cmp_b <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(operator_66_true_div_cmp_b_9_0));
  operator_66_true_div_cmp_z <= operator_66_true_div_cmp_z_1;

  STAGE_LOOP_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 10
      )
    PORT MAP(
      a => STAGE_LOOP_lshift_rg_a,
      s => STAGE_LOOP_lshift_rg_s,
      z => STAGE_LOOP_lshift_rg_z
    );
  STAGE_LOOP_lshift_rg_a(0) <= '1';
  STAGE_LOOP_lshift_rg_s <= STAGE_LOOP_i_3_0_sva;
  STAGE_LOOP_lshift_psp_sva_mx0w0 <= STAGE_LOOP_lshift_rg_z;

  inPlaceNTT_DIT_core_core_fsm_inst : inPlaceNTT_DIT_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => inPlaceNTT_DIT_core_core_fsm_inst_fsm_output,
      STAGE_LOOP_C_8_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0,
      modExp_while_C_38_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_1_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_1_while_C_38_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_62_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0,
      COMP_LOOP_2_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_124_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0,
      COMP_LOOP_3_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_186_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0,
      COMP_LOOP_4_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_248_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0,
      COMP_LOOP_5_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_310_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0,
      COMP_LOOP_6_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_372_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0,
      COMP_LOOP_7_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_434_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0,
      COMP_LOOP_8_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_496_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_496_tr0,
      COMP_LOOP_9_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_558_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_558_tr0,
      COMP_LOOP_10_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_620_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_620_tr0,
      COMP_LOOP_11_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_682_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_682_tr0,
      COMP_LOOP_12_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_744_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_744_tr0,
      COMP_LOOP_13_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_806_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_806_tr0,
      COMP_LOOP_14_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_868_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_868_tr0,
      COMP_LOOP_15_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_930_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_930_tr0,
      COMP_LOOP_16_modExp_1_while_C_38_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_992_tr0 => COMP_LOOP_COMP_LOOP_and_10_itm,
      VEC_LOOP_C_0_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_9_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0
    );
  fsm_output <= inPlaceNTT_DIT_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 <= NOT (z_out_7(64));
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 <= NOT COMP_LOOP_nor_11_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_62_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_124_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_186_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_248_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_310_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_372_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_434_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_496_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_558_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_620_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_682_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_744_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_806_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_868_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_930_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 <= z_out_6(12);
  inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 <= NOT STAGE_LOOP_acc_itm_2_1;

  nand_360_nl <= NOT((fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9)) AND
      (fsm_output(8)) AND (NOT (fsm_output(10))));
  or_619_nl <= (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR not_tmp_51;
  mux_1092_nl <= MUX_s_1_2_2(nand_360_nl, or_619_nl, fsm_output(0));
  or_621_cse <= (fsm_output(5)) OR mux_1092_nl;
  or_596_cse <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR not_tmp_51;
  nor_223_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  and_574_cse <= (fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(1));
  or_2348_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  and_573_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_563_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  or_2385_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  and_565_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  nand_257_cse <= NOT((fsm_output(8)) AND (fsm_output(6)));
  nand_375_cse <= NOT((fsm_output(7)) AND (fsm_output(9)) AND (fsm_output(10)));
  or_495_cse <= CONV_SL_1_1(fsm_output(6 DOWNTO 2)/=STD_LOGIC_VECTOR'("00000"));
  nand_376_cse <= NOT(CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("11")));
  nor_412_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")));
  and_528_cse <= (fsm_output(6)) AND (fsm_output(3));
  nor_422_cse <= NOT((fsm_output(3)) OR (NOT (fsm_output(6))));
  and_472_cse <= (fsm_output(9)) AND (fsm_output(4));
  or_2778_nl <= (fsm_output(7)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(4)))
      OR (fsm_output(10));
  mux_3143_cse <= MUX_s_1_2_2(or_tmp_2516, or_2778_nl, fsm_output(9));
  nor_637_nl <= NOT((NOT (fsm_output(9))) OR (NOT (fsm_output(7))) OR (fsm_output(2))
      OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_638_nl <= NOT((fsm_output(9)) OR (fsm_output(7)) OR (NOT (fsm_output(2))) OR
      (fsm_output(4)) OR (NOT (fsm_output(10))));
  mux_3145_nl <= MUX_s_1_2_2(nor_637_nl, nor_638_nl, fsm_output(5));
  and_466_nl <= (fsm_output(1)) AND mux_3145_nl;
  nor_639_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR
      (NOT (fsm_output(7))) OR (fsm_output(2)) OR nand_398_cse);
  mux_3146_nl <= MUX_s_1_2_2(and_466_nl, nor_639_nl, fsm_output(6));
  and_467_nl <= (fsm_output(6)) AND (fsm_output(1)) AND (fsm_output(5)) AND (NOT
      (fsm_output(9))) AND (fsm_output(7)) AND (fsm_output(2)) AND (fsm_output(4))
      AND (NOT (fsm_output(10)));
  mux_3147_nl <= MUX_s_1_2_2(mux_3146_nl, and_467_nl, fsm_output(3));
  nor_640_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (NOT (fsm_output(7))) OR (fsm_output(2)) OR nand_398_cse);
  nor_641_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR mux_3143_cse);
  mux_3144_nl <= MUX_s_1_2_2(nor_640_nl, nor_641_nl, fsm_output(6));
  and_468_nl <= (fsm_output(3)) AND mux_3144_nl;
  mux_3148_nl <= MUX_s_1_2_2(mux_3147_nl, and_468_nl, fsm_output(8));
  nor_642_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (fsm_output(7)) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  and_469_nl <= (fsm_output(1)) AND (fsm_output(5)) AND (fsm_output(9)) AND (fsm_output(7))
      AND (fsm_output(2)) AND (fsm_output(4)) AND (NOT (fsm_output(10)));
  mux_3140_nl <= MUX_s_1_2_2(nor_642_nl, and_469_nl, fsm_output(6));
  or_2773_nl <= (fsm_output(9)) OR (NOT (fsm_output(7))) OR (fsm_output(2)) OR (NOT
      (fsm_output(4))) OR (fsm_output(10));
  or_2772_nl <= (NOT (fsm_output(9))) OR (fsm_output(7)) OR (NOT (fsm_output(2)))
      OR (fsm_output(4)) OR (fsm_output(10));
  mux_3138_nl <= MUX_s_1_2_2(or_2773_nl, or_2772_nl, fsm_output(5));
  or_2770_nl <= (NOT (fsm_output(7))) OR (fsm_output(2)) OR (fsm_output(4)) OR (NOT
      (fsm_output(10)));
  mux_3137_nl <= MUX_s_1_2_2(or_2770_nl, or_tmp_2707, fsm_output(9));
  or_2771_nl <= (fsm_output(5)) OR mux_3137_nl;
  mux_3139_nl <= MUX_s_1_2_2(mux_3138_nl, or_2771_nl, fsm_output(1));
  nor_643_nl <= NOT((fsm_output(6)) OR mux_3139_nl);
  mux_3141_nl <= MUX_s_1_2_2(mux_3140_nl, nor_643_nl, fsm_output(3));
  mux_3135_nl <= MUX_s_1_2_2(or_tmp_2707, or_tmp_2516, fsm_output(9));
  nor_644_nl <= NOT((fsm_output(5)) OR mux_3135_nl);
  nor_645_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(7)) OR
      (fsm_output(2)) OR (fsm_output(4)) OR (fsm_output(10)));
  mux_3136_nl <= MUX_s_1_2_2(nor_644_nl, nor_645_nl, fsm_output(1));
  and_470_nl <= nor_422_cse AND mux_3136_nl;
  mux_3142_nl <= MUX_s_1_2_2(mux_3141_nl, and_470_nl, fsm_output(8));
  mux_3149_nl <= MUX_s_1_2_2(mux_3148_nl, mux_3142_nl, fsm_output(0));
  and_353_nl <= mux_3149_nl AND COMP_LOOP_nor_11_itm;
  modExp_while_if_and_nl <= modExp_while_and_3 AND not_tmp_646;
  modExp_while_if_and_1_nl <= modExp_while_and_5 AND not_tmp_646;
  modExp_while_if_mux1h_nl <= MUX1HOT_v_64_6_2(z_out_10, STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
      COMP_LOOP_1_modExp_1_while_if_mul_mut_1, modulo_result_rem_cmp_z, (z_out_6(63
      DOWNTO 0)), z_out_5, STD_LOGIC_VECTOR'( and_dcpl_260 & not_tmp_596 & and_353_nl
      & modExp_while_if_and_nl & modExp_while_if_and_1_nl & (NOT mux_2475_itm)));
  and_284_nl <= and_dcpl_118 AND and_dcpl_98;
  mux_2560_nl <= MUX_s_1_2_2(not_tmp_529, mux_tmp_2502, fsm_output(1));
  mux_2559_nl <= MUX_s_1_2_2(mux_tmp_2519, nor_tmp_342, and_573_cse);
  mux_2561_nl <= MUX_s_1_2_2(mux_2560_nl, mux_2559_nl, fsm_output(9));
  and_532_nl <= (fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(10));
  and_533_nl <= (and_565_cse OR (fsm_output(3))) AND (fsm_output(10));
  mux_2558_nl <= MUX_s_1_2_2(and_532_nl, and_533_nl, fsm_output(9));
  mux_2562_nl <= MUX_s_1_2_2(mux_2561_nl, mux_2558_nl, fsm_output(6));
  mux_2556_nl <= MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, or_3308_cse);
  or_2494_nl <= (fsm_output(9)) OR (NOT mux_2556_nl);
  mux_2553_nl <= MUX_s_1_2_2(mux_tmp_2519, nor_tmp_342, fsm_output(1));
  and_535_nl <= (and_563_cse OR (fsm_output(3))) AND (fsm_output(10));
  mux_2554_nl <= MUX_s_1_2_2(mux_2553_nl, and_535_nl, fsm_output(0));
  or_2491_nl <= nor_784_cse OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR
      (fsm_output(10));
  mux_2555_nl <= MUX_s_1_2_2((NOT mux_2554_nl), or_2491_nl, fsm_output(9));
  mux_2557_nl <= MUX_s_1_2_2(or_2494_nl, mux_2555_nl, fsm_output(6));
  mux_2563_nl <= MUX_s_1_2_2(mux_2562_nl, mux_2557_nl, fsm_output(7));
  mux_2551_nl <= MUX_s_1_2_2(and_816_cse, mux_tmp_2549, fsm_output(6));
  nor_731_nl <= NOT(and_563_cse OR (fsm_output(3)) OR (fsm_output(10)));
  mux_2548_nl <= MUX_s_1_2_2(nor_731_nl, (fsm_output(10)), fsm_output(9));
  mux_2550_nl <= MUX_s_1_2_2(mux_tmp_2549, mux_2548_nl, fsm_output(6));
  mux_2552_nl <= MUX_s_1_2_2(mux_2551_nl, mux_2550_nl, fsm_output(7));
  mux_2564_nl <= MUX_s_1_2_2(mux_2563_nl, mux_2552_nl, fsm_output(8));
  mux_2544_nl <= MUX_s_1_2_2(nor_tmp_342, or_tmp_2429, fsm_output(9));
  mux_2542_nl <= MUX_s_1_2_2(nor_tmp_338, or_tmp_2416, fsm_output(0));
  mux_2543_nl <= MUX_s_1_2_2((NOT mux_2542_nl), mux_tmp_2502, fsm_output(9));
  mux_2545_nl <= MUX_s_1_2_2((NOT mux_2544_nl), mux_2543_nl, fsm_output(6));
  mux_2540_nl <= MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, and_563_cse);
  or_2484_nl <= (fsm_output(9)) OR (NOT mux_2540_nl);
  mux_2541_nl <= MUX_s_1_2_2(and_816_cse, or_2484_nl, fsm_output(6));
  mux_2546_nl <= MUX_s_1_2_2(mux_2545_nl, mux_2541_nl, fsm_output(7));
  mux_2536_nl <= MUX_s_1_2_2(mux_tmp_2502, mux_tmp_2523, fsm_output(1));
  mux_2537_nl <= MUX_s_1_2_2(mux_2536_nl, mux_tmp_2525, fsm_output(0));
  or_2483_nl <= (fsm_output(9)) OR (NOT mux_2537_nl);
  nor_732_nl <= NOT((fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(3))
      OR (fsm_output(10)));
  mux_2535_nl <= MUX_s_1_2_2(nor_732_nl, (fsm_output(10)), fsm_output(9));
  mux_2538_nl <= MUX_s_1_2_2(or_2483_nl, mux_2535_nl, fsm_output(6));
  or_2480_nl <= (or_3308_cse AND (fsm_output(3))) OR (fsm_output(10));
  mux_2534_nl <= MUX_s_1_2_2(nor_tmp_338, or_2480_nl, fsm_output(9));
  mux_2539_nl <= MUX_s_1_2_2(mux_2538_nl, mux_2534_nl, fsm_output(7));
  mux_2547_nl <= MUX_s_1_2_2(mux_2546_nl, mux_2539_nl, fsm_output(8));
  mux_2565_nl <= MUX_s_1_2_2(mux_2564_nl, mux_2547_nl, fsm_output(5));
  mux_2528_nl <= MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, and_540_cse);
  mux_2529_nl <= MUX_s_1_2_2(not_tmp_529, mux_2528_nl, fsm_output(9));
  mux_2524_nl <= MUX_s_1_2_2(mux_tmp_2523, mux_tmp_2519, fsm_output(1));
  mux_2526_nl <= MUX_s_1_2_2(mux_tmp_2525, mux_2524_nl, fsm_output(0));
  mux_2527_nl <= MUX_s_1_2_2(not_tmp_529, mux_2526_nl, fsm_output(9));
  mux_2530_nl <= MUX_s_1_2_2(mux_2529_nl, mux_2527_nl, fsm_output(6));
  nor_733_nl <= NOT(and_565_cse OR (fsm_output(3)) OR (fsm_output(10)));
  mux_2521_nl <= MUX_s_1_2_2(nor_733_nl, (fsm_output(10)), fsm_output(9));
  mux_2520_nl <= MUX_s_1_2_2(mux_tmp_2519, or_tmp_2419, fsm_output(9));
  mux_2522_nl <= MUX_s_1_2_2(mux_2521_nl, mux_2520_nl, fsm_output(6));
  mux_2531_nl <= MUX_s_1_2_2((NOT mux_2530_nl), mux_2522_nl, fsm_output(7));
  mux_2516_nl <= MUX_s_1_2_2(nor_tmp_6, or_tmp_2419, fsm_output(9));
  or_2475_nl <= (NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))))
      OR (NOT (fsm_output(3))) OR (fsm_output(10));
  mux_2515_nl <= MUX_s_1_2_2((NOT nor_tmp_330), or_2475_nl, fsm_output(9));
  mux_2517_nl <= MUX_s_1_2_2(mux_2516_nl, mux_2515_nl, fsm_output(6));
  or_2472_nl <= (NOT(and_565_cse OR (fsm_output(3)))) OR (fsm_output(10));
  mux_2513_nl <= MUX_s_1_2_2((NOT or_tmp_2416), or_2472_nl, fsm_output(9));
  mux_2514_nl <= MUX_s_1_2_2(mux_2513_nl, and_816_cse, fsm_output(6));
  mux_2518_nl <= MUX_s_1_2_2(mux_2517_nl, mux_2514_nl, fsm_output(7));
  mux_2532_nl <= MUX_s_1_2_2(mux_2531_nl, mux_2518_nl, fsm_output(8));
  mux_2510_nl <= MUX_s_1_2_2(nor_1203_cse, mux_tmp_2508, fsm_output(6));
  or_2466_nl <= (NOT(and_540_cse OR (fsm_output(3)))) OR (fsm_output(10));
  mux_2507_nl <= MUX_s_1_2_2(not_tmp_529, or_2466_nl, fsm_output(9));
  mux_2509_nl <= MUX_s_1_2_2(mux_tmp_2508, mux_2507_nl, fsm_output(6));
  mux_2511_nl <= MUX_s_1_2_2(mux_2510_nl, mux_2509_nl, fsm_output(7));
  mux_2503_nl <= MUX_s_1_2_2(not_tmp_529, mux_tmp_2502, or_2348_cse);
  or_2460_nl <= nor_738_cse OR (fsm_output(10));
  mux_2504_nl <= MUX_s_1_2_2(mux_2503_nl, or_2460_nl, fsm_output(9));
  and_544_nl <= or_2348_cse AND (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(10));
  mux_2500_nl <= MUX_s_1_2_2(and_544_nl, (fsm_output(10)), fsm_output(9));
  mux_2505_nl <= MUX_s_1_2_2(mux_2504_nl, mux_2500_nl, fsm_output(6));
  nand_247_nl <= NOT((fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(2)) AND
      (fsm_output(3)) AND (NOT (fsm_output(10))));
  mux_2498_nl <= MUX_s_1_2_2((NOT nor_tmp_6), nand_247_nl, fsm_output(9));
  nand_248_nl <= NOT((and_540_cse OR (fsm_output(3))) AND (fsm_output(10)));
  or_2454_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(10));
  mux_2497_nl <= MUX_s_1_2_2(nand_248_nl, or_2454_nl, fsm_output(9));
  mux_2499_nl <= MUX_s_1_2_2(mux_2498_nl, mux_2497_nl, fsm_output(6));
  mux_2506_nl <= MUX_s_1_2_2(mux_2505_nl, mux_2499_nl, fsm_output(7));
  mux_2512_nl <= MUX_s_1_2_2(mux_2511_nl, mux_2506_nl, fsm_output(8));
  mux_2533_nl <= MUX_s_1_2_2(mux_2532_nl, mux_2512_nl, fsm_output(5));
  mux_2566_nl <= MUX_s_1_2_2(mux_2565_nl, mux_2533_nl, fsm_output(4));
  operator_64_false_mux1h_2_rgt <= MUX1HOT_v_65_3_2(z_out_6, (STD_LOGIC_VECTOR'(
      "00") & operator_64_false_slc_modExp_exp_63_1_3), ('0' & modExp_while_if_mux1h_nl),
      STD_LOGIC_VECTOR'( and_284_nl & and_dcpl_273 & (NOT mux_2566_nl)));
  and_1262_cse <= (fsm_output(3)) AND (fsm_output(9));
  nor_1450_cse <= NOT((NOT (fsm_output(1))) OR COMP_LOOP_nor_11_itm);
  or_3328_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00"));
  or_2520_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  and_754_cse <= or_3328_cse AND (fsm_output(10));
  and_300_m1c <= and_dcpl_191 AND and_dcpl_279;
  and_816_cse <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)=STD_LOGIC_VECTOR'("11"));
  and_815_cse <= (fsm_output(7)) AND (fsm_output(9)) AND (fsm_output(10));
  modExp_result_and_rgt <= (NOT modExp_while_and_5) AND and_300_m1c;
  modExp_result_and_1_rgt <= modExp_while_and_5 AND and_300_m1c;
  or_15_cse <= (NOT((fsm_output(6)) OR (NOT (fsm_output(3))))) OR (fsm_output(10));
  nand_402_cse <= NOT((fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(1)) AND
      (NOT (fsm_output(10))));
  mux_28_cse <= MUX_s_1_2_2((NOT (fsm_output(10))), or_tmp_21, fsm_output(6));
  or_36_cse <= (fsm_output(6)) OR (NOT nor_tmp_6);
  mux_3_cse <= MUX_s_1_2_2(or_tmp_4, or_tmp_3, fsm_output(7));
  mux_7_cse <= MUX_s_1_2_2(or_tmp_9, (fsm_output(10)), fsm_output(6));
  mux_9_cse <= MUX_s_1_2_2((fsm_output(10)), nand_402_cse, fsm_output(6));
  nand_240_cse <= NOT((fsm_output(7)) AND (fsm_output(4)) AND (fsm_output(10)));
  or_2591_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR (fsm_output(9))
      OR (fsm_output(2)) OR nand_240_cse;
  or_2588_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(7))
      OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  mux_2767_nl <= MUX_s_1_2_2(mux_3143_cse, or_2588_nl, fsm_output(1));
  or_2589_nl <= (fsm_output(5)) OR mux_2767_nl;
  mux_2768_nl <= MUX_s_1_2_2(or_2591_nl, or_2589_nl, fsm_output(6));
  nor_694_nl <= NOT((fsm_output(3)) OR mux_2768_nl);
  nor_695_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(1))) OR mux_3143_cse);
  nor_696_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(1)) OR mux_tmp_2758);
  mux_2766_nl <= MUX_s_1_2_2(nor_695_nl, nor_696_nl, fsm_output(6));
  and_513_nl <= (fsm_output(3)) AND mux_2766_nl;
  mux_2769_nl <= MUX_s_1_2_2(nor_694_nl, and_513_nl, fsm_output(8));
  nor_697_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(1)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  or_2581_nl <= (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(4))
      OR (NOT (fsm_output(10)));
  or_2579_nl <= (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(4)))
      OR (fsm_output(10));
  mux_2762_nl <= MUX_s_1_2_2(or_2581_nl, or_2579_nl, fsm_output(1));
  nor_698_nl <= NOT((fsm_output(5)) OR mux_2762_nl);
  mux_2763_nl <= MUX_s_1_2_2(nor_697_nl, nor_698_nl, fsm_output(6));
  and_514_nl <= (fsm_output(3)) AND mux_2763_nl;
  and_515_nl <= (fsm_output(1)) AND (NOT mux_tmp_2758);
  nor_699_nl <= NOT((fsm_output(1)) OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR
      (fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(10)));
  mux_2759_nl <= MUX_s_1_2_2(and_515_nl, nor_699_nl, fsm_output(5));
  nor_700_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(1)) OR (fsm_output(9)) OR
      (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  mux_2760_nl <= MUX_s_1_2_2(mux_2759_nl, nor_700_nl, fsm_output(6));
  nor_701_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(1)))
      OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(4))
      OR (fsm_output(10)));
  mux_2761_nl <= MUX_s_1_2_2(mux_2760_nl, nor_701_nl, fsm_output(3));
  mux_2764_nl <= MUX_s_1_2_2(and_514_nl, mux_2761_nl, fsm_output(8));
  mux_2770_m1c <= MUX_s_1_2_2(mux_2769_nl, mux_2764_nl, fsm_output(0));
  and_517_cse <= (fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(3));
  nand_398_cse <= NOT((fsm_output(4)) AND (fsm_output(10)));
  nand_237_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")));
  modulo_result_mux_1_cse <= MUX_v_64_2_2(modulo_result_rem_cmp_z, (z_out_6(63 DOWNTO
      0)), modulo_result_rem_cmp_z(63));
  nor_1302_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(4)) OR (fsm_output(10)));
  and_801_nl <= (fsm_output(7)) AND (fsm_output(9)) AND (fsm_output(8)) AND (fsm_output(4))
      AND (NOT (fsm_output(10)));
  mux_71_cse <= MUX_s_1_2_2(nor_1302_nl, and_801_nl, fsm_output(2));
  nor_715_nl <= NOT((fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(3)));
  mux_2742_nl <= MUX_s_1_2_2(and_517_cse, nor_715_nl, fsm_output(5));
  and_345_m1c <= mux_2742_nl AND and_dcpl_26 AND (NOT (fsm_output(7))) AND (NOT (fsm_output(2)))
      AND (NOT (fsm_output(8))) AND and_dcpl_30;
  or_2679_cse <= (fsm_output(8)) OR (NOT (fsm_output(9))) OR (fsm_output(5)) OR (fsm_output(10));
  nor_381_cse <= NOT((fsm_output(4)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(6))));
  nor_670_cse <= NOT((NOT (fsm_output(8))) OR (fsm_output(9)) OR (fsm_output(5))
      OR (fsm_output(10)));
  or_212_cse <= (fsm_output(8)) OR (fsm_output(4));
  and_491_cse <= (fsm_output(4)) AND (fsm_output(10));
  or_2729_cse <= (fsm_output(8)) OR and_491_cse;
  or_199_nl <= (fsm_output(8)) OR (NOT or_tmp_182);
  mux_384_cse <= MUX_s_1_2_2(or_199_nl, nand_tmp_12, fsm_output(6));
  mux_382_cse <= MUX_s_1_2_2(mux_tmp_381, mux_tmp_379, fsm_output(1));
  COMP_LOOP_or_32_cse <= and_dcpl_126 OR and_dcpl_141 OR and_dcpl_147 OR and_dcpl_158
      OR and_dcpl_164 OR and_dcpl_175 OR and_dcpl_182 OR and_dcpl_192 OR and_dcpl_198
      OR and_dcpl_206 OR and_dcpl_217 OR and_dcpl_225 OR and_dcpl_232 OR and_dcpl_242
      OR and_dcpl_247 OR and_dcpl_255;
  or_2824_cse <= (fsm_output(3)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(4))) OR (fsm_output(10));
  nand_226_cse <= NOT((fsm_output(3)) AND (fsm_output(1)) AND (fsm_output(9)) AND
      (fsm_output(4)) AND (fsm_output(10)));
  or_2826_cse <= (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(4))
      OR (NOT (fsm_output(10)));
  or_2839_cse <= (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(1)))
      OR (fsm_output(9)) OR (fsm_output(4)) OR (fsm_output(10));
  and_464_cse <= (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(1)) AND (fsm_output(9))
      AND (fsm_output(4)) AND (NOT (fsm_output(10)));
  or_2819_cse <= (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(9))
      OR nand_398_cse;
  or_2894_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"));
  and_458_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"));
  and_459_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"));
  and_359_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11")) AND
      or_2894_cse;
  and_456_cse <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"));
  or_2898_cse <= (fsm_output(3)) OR (fsm_output(6));
  and_450_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  or_2902_cse <= and_573_cse OR (fsm_output(3));
  nor_1316_cse <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000")));
  nor_610_cse <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00")));
  and_440_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
  or_2935_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  mux_726_cse <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), fsm_output(9));
  or_3308_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  or_2951_cse <= CONV_SL_1_1(fsm_output(8 DOWNTO 6)/=STD_LOGIC_VECTOR'("000"));
  nor_1203_cse <= NOT((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(10)));
  nor_601_cse <= NOT(CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00")));
  or_3002_cse <= (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(8)) OR (NOT (fsm_output(4)))
      OR (fsm_output(10));
  or_3018_cse <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(8)) OR nand_398_cse;
  or_3016_cse <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR not_tmp_34;
  or_3014_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(7)) OR (NOT
      (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  mux_3393_nl <= MUX_s_1_2_2(or_3016_cse, or_3014_nl, fsm_output(5));
  mux_3394_cse <= MUX_s_1_2_2(or_3018_cse, mux_3393_nl, fsm_output(0));
  or_3004_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(8)) OR (fsm_output(4))
      OR (NOT (fsm_output(10)));
  mux_3384_nl <= MUX_s_1_2_2(or_3004_nl, or_3002_cse, fsm_output(1));
  or_3001_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  mux_3385_cse <= MUX_s_1_2_2(mux_3384_nl, or_3001_nl, fsm_output(5));
  nor_581_nl <= NOT((fsm_output(0)) OR mux_tmp_3386);
  nor_582_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR (fsm_output(2))
      OR (fsm_output(7)) OR not_tmp_34);
  nor_583_nl <= NOT((fsm_output(7)) OR (fsm_output(8)) OR (fsm_output(4)) OR (NOT
      (fsm_output(10))));
  and_415_nl <= (fsm_output(7)) AND (fsm_output(8)) AND (fsm_output(4)) AND (fsm_output(10));
  mux_3389_nl <= MUX_s_1_2_2(nor_583_nl, and_415_nl, fsm_output(2));
  and_414_nl <= (fsm_output(1)) AND mux_3389_nl;
  nor_584_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10)));
  mux_3390_nl <= MUX_s_1_2_2(and_414_nl, nor_584_nl, fsm_output(5));
  mux_3391_nl <= MUX_s_1_2_2(nor_582_nl, mux_3390_nl, fsm_output(0));
  mux_3392_cse <= MUX_s_1_2_2(nor_581_nl, mux_3391_nl, fsm_output(6));
  and_416_nl <= (fsm_output(0)) AND (NOT mux_tmp_3386);
  nor_585_nl <= NOT((fsm_output(0)) OR mux_3385_cse);
  mux_3387_nl <= MUX_s_1_2_2(and_416_nl, nor_585_nl, fsm_output(6));
  nor_586_nl <= NOT((fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(8))) OR (NOT
      (fsm_output(4))) OR (fsm_output(10)));
  mux_3388_cse <= MUX_s_1_2_2(mux_3387_nl, nor_586_nl, fsm_output(3));
  or_3241_nl <= (fsm_output(7)) OR (fsm_output(8)) OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  nand_205_nl <= NOT((fsm_output(7)) AND (fsm_output(8)) AND (fsm_output(4)) AND
      (fsm_output(10)));
  mux_3498_cse <= MUX_s_1_2_2(or_3241_nl, nand_205_nl, fsm_output(2));
  mux_3556_nl <= MUX_s_1_2_2(nand_tmp_157, nand_tmp_12, fsm_output(1));
  mux_3557_cse <= MUX_s_1_2_2(or_tmp_191, mux_3556_nl, fsm_output(6));
  mux_3056_nl <= MUX_s_1_2_2(and_491_cse, (fsm_output(4)), fsm_output(9));
  or_3120_nl <= (fsm_output(8)) OR mux_3056_nl;
  mux_3572_nl <= MUX_s_1_2_2(or_2729_cse, or_3120_nl, fsm_output(1));
  mux_3573_nl <= MUX_s_1_2_2(nand_tmp_157, mux_3572_nl, fsm_output(6));
  mux_433_nl <= MUX_s_1_2_2((NOT mux_tmp_380), or_tmp_182, fsm_output(8));
  or_3119_nl <= (fsm_output(8)) OR (NOT mux_tmp_380);
  mux_3569_nl <= MUX_s_1_2_2(mux_433_nl, or_3119_nl, and_573_cse);
  mux_3567_nl <= MUX_s_1_2_2(nand_tmp_14, nand_tmp_157, fsm_output(1));
  mux_3570_nl <= MUX_s_1_2_2(mux_3569_nl, mux_3567_nl, fsm_output(6));
  mux_3574_nl <= MUX_s_1_2_2(mux_3573_nl, mux_3570_nl, fsm_output(5));
  mux_437_nl <= MUX_s_1_2_2(mux_tmp_399, mux_tmp_375, or_2348_cse);
  mux_438_nl <= MUX_s_1_2_2(mux_437_nl, nand_tmp_14, fsm_output(6));
  mux_431_nl <= MUX_s_1_2_2(or_tmp_189, mux_tmp_399, fsm_output(6));
  mux_3566_nl <= MUX_s_1_2_2(mux_438_nl, mux_431_nl, fsm_output(5));
  mux_3575_cse <= MUX_s_1_2_2(mux_3574_nl, mux_3566_nl, fsm_output(7));
  mux_3554_nl <= MUX_s_1_2_2(mux_tmp_373, nand_tmp_157, fsm_output(6));
  mux_419_nl <= MUX_s_1_2_2(or_tmp_188, mux_tmp_381, or_2348_cse);
  mux_420_nl <= MUX_s_1_2_2(mux_419_nl, mux_tmp_375, fsm_output(6));
  mux_3555_cse <= MUX_s_1_2_2(mux_3554_nl, mux_420_nl, fsm_output(5));
  nand_201_cse <= NOT((fsm_output(9)) AND (fsm_output(4)) AND (fsm_output(10)));
  mux_3547_nl <= MUX_s_1_2_2(nand_tmp_157, nand_tmp_12, or_2348_cse);
  mux_3548_nl <= MUX_s_1_2_2(mux_3547_nl, mux_tmp_381, fsm_output(6));
  or_3115_nl <= (fsm_output(8)) OR (NOT mux_tmp_378);
  mux_403_nl <= MUX_s_1_2_2(or_3115_nl, or_tmp_191, or_2348_cse);
  mux_3546_nl <= MUX_s_1_2_2(mux_403_nl, nand_tmp_157, fsm_output(6));
  mux_3549_nl <= MUX_s_1_2_2(mux_3548_nl, mux_3546_nl, fsm_output(5));
  mux_3542_nl <= MUX_s_1_2_2(nand_tmp_14, nand_tmp_157, and_573_cse);
  mux_3543_nl <= MUX_s_1_2_2(mux_tmp_375, mux_3542_nl, fsm_output(6));
  mux_401_nl <= MUX_s_1_2_2(or_tmp_189, or_tmp_188, and_573_cse);
  mux_400_nl <= MUX_s_1_2_2(mux_tmp_399, mux_tmp_375, fsm_output(1));
  mux_402_nl <= MUX_s_1_2_2(mux_401_nl, mux_400_nl, fsm_output(6));
  mux_3544_nl <= MUX_s_1_2_2(mux_3543_nl, mux_402_nl, fsm_output(5));
  mux_3550_nl <= MUX_s_1_2_2(mux_3549_nl, mux_3544_nl, fsm_output(7));
  nand_173_nl <= NOT((fsm_output(8)) AND (NOT mux_tmp_380));
  mux_3532_nl <= MUX_s_1_2_2(nand_201_cse, mux_tmp_380, fsm_output(8));
  mux_3533_nl <= MUX_s_1_2_2(nand_173_nl, mux_3532_nl, fsm_output(1));
  mux_3534_nl <= MUX_s_1_2_2(mux_3533_nl, mux_tmp_3323, fsm_output(6));
  mux_3535_nl <= MUX_s_1_2_2(mux_3534_nl, mux_384_cse, fsm_output(5));
  mux_3527_nl <= MUX_s_1_2_2(nand_tmp_157, nand_tmp_12, and_573_cse);
  mux_3528_nl <= MUX_s_1_2_2(or_tmp_180, mux_3527_nl, fsm_output(6));
  mux_376_nl <= MUX_s_1_2_2(mux_tmp_375, or_tmp_181, fsm_output(1));
  mux_377_nl <= MUX_s_1_2_2(mux_376_nl, mux_tmp_373, fsm_output(0));
  mux_383_nl <= MUX_s_1_2_2(mux_382_cse, mux_377_nl, fsm_output(6));
  mux_3529_nl <= MUX_s_1_2_2(mux_3528_nl, mux_383_nl, fsm_output(5));
  mux_3536_nl <= MUX_s_1_2_2(mux_3535_nl, mux_3529_nl, fsm_output(7));
  mux_3551_cse <= MUX_s_1_2_2(mux_3550_nl, mux_3536_nl, fsm_output(3));
  nor_544_cse <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(2)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  nor_539_cse <= NOT((fsm_output(7)) OR (NOT (fsm_output(2))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  nor_515_cse <= NOT((fsm_output(5)) OR (NOT (fsm_output(3))));
  nor_540_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(2)) OR (fsm_output(9)) OR
      not_tmp_34);
  mux_3603_cse <= MUX_s_1_2_2(nor_539_cse, nor_540_nl, fsm_output(3));
  nor_545_cse <= NOT((fsm_output(5)) OR (fsm_output(3)) OR (fsm_output(7)) OR (fsm_output(2))
      OR (fsm_output(9)) OR not_tmp_34);
  STAGE_LOOP_i_3_0_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_i_3_0_sva)
      + UNSIGNED'( "0001"), 4));
  COMP_LOOP_acc_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
      DOWNTO 4)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0),
      5), 8), 8));
  or_529_cse <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3)))
      OR (fsm_output(4)) OR (fsm_output(10));
  or_525_cse <= (NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3)))
      OR (fsm_output(4)) OR (fsm_output(10));
  COMP_LOOP_1_modExp_1_while_if_mul_mut_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'(
      SIGNED(operator_64_false_acc_mut_63_0) * SIGNED(COMP_LOOP_10_mul_mut)), 64));
  operator_64_false_slc_modExp_exp_63_1_3 <= MUX_v_63_2_2((operator_66_true_div_cmp_z(63
      DOWNTO 1)), (tmp_10_lpi_4_dfm(63 DOWNTO 1)), and_dcpl_281);
  nor_1276_cse <= NOT((fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (fsm_output(10)));
  nor_1279_cse <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(9))
      OR (fsm_output(10)));
  COMP_LOOP_acc_1_cse_6_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0101")), 9), 12), 12));
  COMP_LOOP_acc_1_cse_2_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0001")), 9), 12), 12));
  or_163_cse <= (fsm_output(4)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  COMP_LOOP_k_9_4_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0),
      5), 6) + UNSIGNED'( "000001"), 6));
  modExp_while_and_3 <= (NOT (modulo_result_rem_cmp_z(63))) AND COMP_LOOP_nor_11_itm;
  modExp_while_and_5 <= (modulo_result_rem_cmp_z(63)) AND COMP_LOOP_nor_11_itm;
  or_tmp_3 <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(10));
  or_tmp_4 <= (NOT (fsm_output(6))) OR (fsm_output(10));
  or_tmp_8 <= nor_422_cse OR (fsm_output(10));
  or_tmp_9 <= (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(10));
  or_tmp_14 <= (fsm_output(6)) OR (fsm_output(10));
  nor_tmp_6 <= (fsm_output(3)) AND (fsm_output(10));
  or_tmp_21 <= (fsm_output(3)) OR (fsm_output(10));
  nor_tmp_9 <= ((fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3))) AND (fsm_output(10));
  not_tmp_34 <= NOT((fsm_output(8)) AND (fsm_output(4)) AND (fsm_output(10)));
  not_tmp_45 <= NOT((fsm_output(5)) AND (fsm_output(10)));
  or_tmp_110 <= (fsm_output(8)) OR (fsm_output(10));
  not_tmp_51 <= NOT((fsm_output(8)) AND (fsm_output(10)));
  or_tmp_118 <= (NOT (fsm_output(8))) OR (fsm_output(10));
  or_tmp_141 <= (fsm_output(4)) OR (fsm_output(8)) OR (fsm_output(10));
  or_154_cse <= (NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_tmp_207 <= MUX_s_1_2_2(or_154_cse, or_tmp_141, fsm_output(5));
  mux_tmp_226 <= MUX_s_1_2_2(or_tmp_141, or_tmp_118, fsm_output(5));
  or_tmp_150 <= (NOT (fsm_output(4))) OR (fsm_output(8));
  or_tmp_178 <= (NOT (fsm_output(4))) OR (fsm_output(10));
  or_tmp_179 <= (fsm_output(4)) OR (fsm_output(10));
  mux_371_nl <= MUX_s_1_2_2((NOT or_tmp_179), or_tmp_178, fsm_output(9));
  or_tmp_180 <= (fsm_output(8)) OR mux_371_nl;
  mux_372_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), or_tmp_178, fsm_output(9));
  or_tmp_181 <= (fsm_output(8)) OR mux_372_nl;
  mux_tmp_373 <= MUX_s_1_2_2(or_tmp_181, or_tmp_180, fsm_output(1));
  or_tmp_182 <= (fsm_output(9)) OR (fsm_output(4)) OR (fsm_output(10));
  mux_tmp_374 <= MUX_s_1_2_2((NOT and_491_cse), or_tmp_178, fsm_output(9));
  mux_tmp_375 <= MUX_s_1_2_2(mux_tmp_374, or_tmp_182, fsm_output(8));
  or_tmp_183 <= (fsm_output(9)) OR (NOT and_491_cse);
  mux_tmp_378 <= MUX_s_1_2_2((fsm_output(4)), or_tmp_179, fsm_output(9));
  mux_tmp_379 <= MUX_s_1_2_2(mux_tmp_378, or_tmp_183, fsm_output(8));
  mux_tmp_380 <= MUX_s_1_2_2(and_491_cse, or_tmp_179, fsm_output(9));
  mux_tmp_381 <= MUX_s_1_2_2(mux_tmp_380, or_tmp_183, fsm_output(8));
  or_2747_cse <= (fsm_output(9)) OR (fsm_output(4));
  nor_tmp_46 <= or_2747_cse AND (fsm_output(10));
  nand_tmp_12 <= NOT((fsm_output(8)) AND (NOT nor_tmp_46));
  nand_tmp_13 <= NOT((fsm_output(8)) AND (NOT and_816_cse));
  or_tmp_187 <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_399 <= MUX_s_1_2_2(or_tmp_183, or_tmp_179, fsm_output(8));
  or_tmp_188 <= (fsm_output(8)) OR mux_tmp_380;
  or_tmp_189 <= (fsm_output(8)) OR nor_tmp_46;
  or_tmp_191 <= (fsm_output(8)) OR (NOT or_tmp_179);
  mux_406_nl <= MUX_s_1_2_2(or_tmp_179, (NOT (fsm_output(10))), fsm_output(9));
  nand_tmp_14 <= NOT((fsm_output(8)) AND mux_406_nl);
  or_tmp_195 <= (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_tmp_412 <= MUX_s_1_2_2(or_tmp_195, nor_tmp_46, fsm_output(8));
  mux_tmp_413 <= MUX_s_1_2_2(or_tmp_195, and_816_cse, fsm_output(8));
  and_dcpl <= NOT((fsm_output(4)) OR (fsm_output(9)));
  and_dcpl_1 <= (fsm_output(5)) AND (fsm_output(2));
  and_dcpl_2 <= and_dcpl_1 AND (NOT (fsm_output(8)));
  or_tmp_237 <= (NOT (fsm_output(3))) OR (fsm_output(10));
  nor_tmp_116 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("11"));
  mux_tmp_741 <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), or_3328_cse);
  or_tmp_434 <= (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_tmp_893 <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), fsm_output(6));
  mux_tmp_917 <= MUX_s_1_2_2(or_tmp_434, or_tmp_4, fsm_output(8));
  and_dcpl_21 <= (NOT (fsm_output(5))) AND (fsm_output(2));
  and_dcpl_22 <= and_dcpl_21 AND (fsm_output(8));
  and_dcpl_26 <= NOT((fsm_output(10)) OR (fsm_output(1)));
  and_dcpl_30 <= (fsm_output(4)) AND (NOT (fsm_output(9)));
  and_dcpl_31 <= (fsm_output(5)) AND (NOT (fsm_output(2)));
  and_dcpl_32 <= and_dcpl_31 AND (fsm_output(8));
  and_dcpl_40 <= and_dcpl_21 AND (NOT (fsm_output(8)));
  and_dcpl_46 <= and_dcpl_31 AND (NOT (fsm_output(8)));
  and_dcpl_50 <= (NOT (fsm_output(4))) AND (fsm_output(9));
  or_3295_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(7)) OR (fsm_output(9))
      OR (fsm_output(10));
  mux_1027_nl <= MUX_s_1_2_2(or_3295_nl, nand_375_cse, or_495_cse);
  not_tmp_219 <= MUX_s_1_2_2(mux_1027_nl, nand_376_cse, fsm_output(8));
  and_dcpl_96 <= NOT((fsm_output(5)) OR (fsm_output(2)));
  and_dcpl_97 <= and_dcpl_96 AND (NOT (fsm_output(8)));
  and_dcpl_98 <= and_dcpl_97 AND and_dcpl;
  and_dcpl_99 <= NOT((fsm_output(0)) OR (fsm_output(6)));
  and_dcpl_100 <= and_dcpl_99 AND (NOT (fsm_output(7)));
  and_dcpl_101 <= NOT((fsm_output(10)) OR (fsm_output(3)));
  and_dcpl_102 <= and_dcpl_101 AND (NOT (fsm_output(1)));
  and_dcpl_103 <= and_dcpl_102 AND and_dcpl_100;
  and_dcpl_106 <= and_dcpl_97 AND and_dcpl_50;
  and_dcpl_107 <= (fsm_output(0)) AND (NOT (fsm_output(6)));
  and_dcpl_108 <= and_dcpl_107 AND (fsm_output(7));
  and_dcpl_109 <= (fsm_output(10)) AND (NOT (fsm_output(3)));
  and_dcpl_110 <= and_dcpl_109 AND (fsm_output(1));
  and_dcpl_111 <= and_dcpl_110 AND and_dcpl_108;
  and_dcpl_116 <= and_dcpl_46 AND and_dcpl_30;
  and_dcpl_117 <= and_dcpl_107 AND (NOT (fsm_output(7)));
  and_dcpl_118 <= and_dcpl_102 AND and_dcpl_117;
  and_dcpl_119 <= and_dcpl_118 AND and_dcpl_116;
  and_dcpl_121 <= (NOT (fsm_output(0))) AND (fsm_output(6));
  and_dcpl_122 <= and_dcpl_121 AND (NOT (fsm_output(7)));
  and_dcpl_123 <= (NOT (fsm_output(10))) AND (fsm_output(3));
  and_dcpl_124 <= and_dcpl_123 AND (fsm_output(1));
  and_dcpl_125 <= and_dcpl_124 AND and_dcpl_122;
  and_dcpl_126 <= and_dcpl_125 AND and_dcpl_97 AND and_dcpl_30;
  and_dcpl_127 <= and_dcpl_99 AND (fsm_output(7));
  and_dcpl_128 <= and_dcpl_101 AND (fsm_output(1));
  and_dcpl_129 <= and_dcpl_128 AND and_dcpl_127;
  or_tmp_453 <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(4))) OR (fsm_output(10));
  and_659_nl <= (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(0));
  nor_1193_nl <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(0)));
  not_tmp_240 <= MUX_s_1_2_2(and_659_nl, nor_1193_nl, fsm_output(4));
  and_dcpl_139 <= and_dcpl_2 AND and_dcpl_30;
  and_dcpl_140 <= and_dcpl_124 AND and_dcpl_108;
  and_dcpl_141 <= and_dcpl_140 AND and_dcpl_139;
  and_dcpl_145 <= and_dcpl_1 AND (fsm_output(8));
  and_dcpl_146 <= and_dcpl_145 AND and_dcpl;
  and_dcpl_147 <= and_dcpl_103 AND and_dcpl_146;
  and_dcpl_148 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_154 <= and_dcpl_96 AND (fsm_output(8));
  and_dcpl_156 <= and_dcpl_123 AND (NOT (fsm_output(1)));
  and_dcpl_158 <= and_dcpl_156 AND and_dcpl_108 AND and_dcpl_154 AND and_dcpl;
  and_dcpl_162 <= and_dcpl_121 AND (fsm_output(7));
  and_dcpl_164 <= and_dcpl_124 AND and_dcpl_162 AND and_dcpl_146;
  and_dcpl_165 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("10"));
  nor_tmp_217 <= (fsm_output(6)) AND (fsm_output(0));
  mux_tmp_1049 <= MUX_s_1_2_2(and_dcpl_99, nor_tmp_217, fsm_output(4));
  and_dcpl_172 <= and_dcpl_97 AND and_472_cse;
  and_dcpl_173 <= nor_tmp_217 AND (NOT (fsm_output(7)));
  and_dcpl_175 <= and_dcpl_128 AND and_dcpl_173 AND and_dcpl_172;
  and_dcpl_182 <= and_dcpl_156 AND and_dcpl_127 AND and_dcpl_46 AND and_472_cse;
  and_dcpl_191 <= and_dcpl_156 AND and_dcpl_117;
  and_dcpl_192 <= and_dcpl_191 AND and_dcpl_22 AND and_472_cse;
  and_dcpl_198 <= and_dcpl_129 AND and_dcpl_154 AND and_dcpl_50;
  and_dcpl_204 <= nor_tmp_217 AND (fsm_output(7));
  and_dcpl_206 <= and_dcpl_128 AND and_dcpl_204 AND and_dcpl_145 AND and_dcpl_50;
  and_dcpl_215 <= nor_tmp_6 AND (NOT (fsm_output(1)));
  and_dcpl_217 <= and_dcpl_215 AND and_dcpl_122 AND and_dcpl_40 AND and_dcpl;
  and_dcpl_223 <= and_dcpl_109 AND (NOT (fsm_output(1)));
  and_dcpl_225 <= and_dcpl_223 AND and_dcpl_108 AND and_dcpl_116;
  and_dcpl_232 <= and_dcpl_110 AND and_dcpl_100 AND and_dcpl_22 AND and_dcpl_30;
  and_dcpl_239 <= and_dcpl_32 AND and_dcpl_30;
  and_dcpl_240 <= nor_tmp_6 AND (fsm_output(1));
  and_dcpl_242 <= and_dcpl_240 AND and_dcpl_173 AND and_dcpl_239;
  and_dcpl_243 <= (fsm_output(10)) AND (NOT (fsm_output(6)));
  and_dcpl_245 <= and_dcpl_32 AND and_dcpl;
  and_dcpl_247 <= and_dcpl_223 AND and_dcpl_162 AND and_dcpl_245;
  and_dcpl_255 <= and_dcpl_223 AND and_dcpl_173 AND and_dcpl_40 AND and_dcpl_50;
  or_tmp_515 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_518 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_579_nl <= (VEC_LOOP_j_sva_11_0(3)) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_578_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_577_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1061_nl <= MUX_s_1_2_2(or_578_nl, or_577_nl, fsm_output(0));
  mux_tmp_1062 <= MUX_s_1_2_2(or_579_nl, mux_1061_nl, fsm_output(5));
  or_587_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_586_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1065_nl <= MUX_s_1_2_2(or_587_nl, or_586_nl, fsm_output(0));
  or_585_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1066_nl <= MUX_s_1_2_2(mux_1065_nl, or_585_nl, fsm_output(5));
  or_583_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1067 <= MUX_s_1_2_2(mux_1066_nl, or_583_nl, fsm_output(4));
  or_591_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_589_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1068 <= MUX_s_1_2_2(or_591_nl, or_589_nl, fsm_output(5));
  or_622_cse <= (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_617_cse <= (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9)))
      OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_614_nl <= (fsm_output(0)) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_613_nl <= (fsm_output(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1087_nl <= MUX_s_1_2_2(or_614_nl, or_613_nl, fsm_output(5));
  or_611_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  or_610_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_1086_nl <= MUX_s_1_2_2(or_611_nl, or_610_nl, fsm_output(5));
  mux_1088_cse <= MUX_s_1_2_2(mux_1087_nl, mux_1086_nl, fsm_output(4));
  or_609_cse <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_607_cse <= (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  nor_1170_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10)));
  nor_1171_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9)))
      OR (fsm_output(8)) OR (fsm_output(10)));
  mux_1080_nl <= MUX_s_1_2_2(nor_1170_nl, nor_1171_nl, fsm_output(0));
  nand_25_cse <= NOT((fsm_output(5)) AND mux_1080_nl);
  or_601_cse <= (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_600_nl <= (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9)))
      OR (fsm_output(8)) OR (fsm_output(10));
  or_599_nl <= (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_1073_cse <= MUX_s_1_2_2(or_600_nl, or_599_nl, fsm_output(0));
  not_tmp_260 <= NOT((fsm_output(1)) AND (fsm_output(10)));
  or_tmp_626 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_630 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_693_nl <= (VEC_LOOP_j_sva_11_0(3)) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_692_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_691_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1138_nl <= MUX_s_1_2_2(or_692_nl, or_691_nl, fsm_output(0));
  mux_tmp_1139 <= MUX_s_1_2_2(or_693_nl, mux_1138_nl, fsm_output(5));
  or_709_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_708_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1148_nl <= MUX_s_1_2_2(or_709_nl, or_708_nl, fsm_output(0));
  or_707_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1149_nl <= MUX_s_1_2_2(mux_1148_nl, or_707_nl, fsm_output(5));
  or_705_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1150 <= MUX_s_1_2_2(mux_1149_nl, or_705_nl, fsm_output(4));
  or_712_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_710_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1152 <= MUX_s_1_2_2(or_712_nl, or_710_nl, fsm_output(5));
  or_tmp_728 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_731 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_792_nl <= (VEC_LOOP_j_sva_11_0(3)) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_791_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_790_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1205_nl <= MUX_s_1_2_2(or_791_nl, or_790_nl, fsm_output(0));
  mux_tmp_1206 <= MUX_s_1_2_2(or_792_nl, mux_1205_nl, fsm_output(5));
  or_800_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_799_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1209_nl <= MUX_s_1_2_2(or_800_nl, or_799_nl, fsm_output(0));
  or_798_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1210_nl <= MUX_s_1_2_2(mux_1209_nl, or_798_nl, fsm_output(5));
  or_796_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_tmp_1211 <= MUX_s_1_2_2(mux_1210_nl, or_796_nl, fsm_output(4));
  or_804_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_802_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1212 <= MUX_s_1_2_2(or_804_nl, or_802_nl, fsm_output(5));
  or_tmp_839 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_843 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_906_nl <= (VEC_LOOP_j_sva_11_0(3)) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_905_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_904_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1282_nl <= MUX_s_1_2_2(or_905_nl, or_904_nl, fsm_output(0));
  mux_tmp_1283 <= MUX_s_1_2_2(or_906_nl, mux_1282_nl, fsm_output(5));
  or_922_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_921_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1292_nl <= MUX_s_1_2_2(or_922_nl, or_921_nl, fsm_output(0));
  nand_433_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0011"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_1293_nl <= MUX_s_1_2_2(mux_1292_nl, nand_433_nl, fsm_output(5));
  or_918_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1294 <= MUX_s_1_2_2(mux_1293_nl, or_918_nl, fsm_output(4));
  or_925_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_923_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1296 <= MUX_s_1_2_2(or_925_nl, or_923_nl, fsm_output(5));
  or_tmp_941 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_944 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1005_nl <= (VEC_LOOP_j_sva_11_0(3)) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1004_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1003_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1349_nl <= MUX_s_1_2_2(or_1004_nl, or_1003_nl, fsm_output(0));
  mux_tmp_1350 <= MUX_s_1_2_2(or_1005_nl, mux_1349_nl, fsm_output(5));
  or_1013_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1012_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1353_nl <= MUX_s_1_2_2(or_1013_nl, or_1012_nl, fsm_output(0));
  or_1011_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1354_nl <= MUX_s_1_2_2(mux_1353_nl, or_1011_nl, fsm_output(5));
  or_1009_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1355 <= MUX_s_1_2_2(mux_1354_nl, or_1009_nl, fsm_output(4));
  or_1017_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1015_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1356 <= MUX_s_1_2_2(or_1017_nl, or_1015_nl, fsm_output(5));
  or_tmp_1052 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_1056 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1119_nl <= (VEC_LOOP_j_sva_11_0(3)) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1118_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1117_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1426_nl <= MUX_s_1_2_2(or_1118_nl, or_1117_nl, fsm_output(0));
  mux_tmp_1427 <= MUX_s_1_2_2(or_1119_nl, mux_1426_nl, fsm_output(5));
  or_1135_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1134_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1436_nl <= MUX_s_1_2_2(or_1135_nl, or_1134_nl, fsm_output(0));
  nand_432_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0101"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_1437_nl <= MUX_s_1_2_2(mux_1436_nl, nand_432_nl, fsm_output(5));
  or_1131_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1438 <= MUX_s_1_2_2(mux_1437_nl, or_1131_nl, fsm_output(4));
  or_1138_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1136_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1440 <= MUX_s_1_2_2(or_1138_nl, or_1136_nl, fsm_output(5));
  or_tmp_1154 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_1157 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1218_nl <= (VEC_LOOP_j_sva_11_0(3)) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1217_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1216_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1493_nl <= MUX_s_1_2_2(or_1217_nl, or_1216_nl, fsm_output(0));
  mux_tmp_1494 <= MUX_s_1_2_2(or_1218_nl, mux_1493_nl, fsm_output(5));
  or_1226_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1225_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1497_nl <= MUX_s_1_2_2(or_1226_nl, or_1225_nl, fsm_output(0));
  nand_431_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0110"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_1498_nl <= MUX_s_1_2_2(mux_1497_nl, nand_431_nl, fsm_output(5));
  or_1222_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_tmp_1499 <= MUX_s_1_2_2(mux_1498_nl, or_1222_nl, fsm_output(4));
  or_1230_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1228_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1500 <= MUX_s_1_2_2(or_1230_nl, or_1228_nl, fsm_output(5));
  or_tmp_1265 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_1269 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1332_nl <= (VEC_LOOP_j_sva_11_0(3)) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1331_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1330_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1570_nl <= MUX_s_1_2_2(or_1331_nl, or_1330_nl, fsm_output(0));
  mux_tmp_1571 <= MUX_s_1_2_2(or_1332_nl, mux_1570_nl, fsm_output(5));
  or_1348_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1347_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1580_nl <= MUX_s_1_2_2(or_1348_nl, or_1347_nl, fsm_output(0));
  nand_430_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_1581_nl <= MUX_s_1_2_2(mux_1580_nl, nand_430_nl, fsm_output(5));
  or_1344_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1582 <= MUX_s_1_2_2(mux_1581_nl, or_1344_nl, fsm_output(4));
  nand_418_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  or_1349_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1584 <= MUX_s_1_2_2(nand_418_nl, or_1349_nl, fsm_output(5));
  or_tmp_1367 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_1370 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1431_nl <= (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1430_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1429_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1637_nl <= MUX_s_1_2_2(or_1430_nl, or_1429_nl, fsm_output(0));
  mux_tmp_1638 <= MUX_s_1_2_2(or_1431_nl, mux_1637_nl, fsm_output(5));
  or_1439_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1438_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1641_nl <= MUX_s_1_2_2(or_1439_nl, or_1438_nl, fsm_output(0));
  or_1437_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1642_nl <= MUX_s_1_2_2(mux_1641_nl, or_1437_nl, fsm_output(5));
  or_1435_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1643 <= MUX_s_1_2_2(mux_1642_nl, or_1435_nl, fsm_output(4));
  or_1443_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1441_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1644 <= MUX_s_1_2_2(or_1443_nl, or_1441_nl, fsm_output(5));
  or_tmp_1478 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_1482 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1545_nl <= (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1544_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1543_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1714_nl <= MUX_s_1_2_2(or_1544_nl, or_1543_nl, fsm_output(0));
  mux_tmp_1715 <= MUX_s_1_2_2(or_1545_nl, mux_1714_nl, fsm_output(5));
  or_1561_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1560_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1724_nl <= MUX_s_1_2_2(or_1561_nl, or_1560_nl, fsm_output(0));
  nand_429_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1001"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_1725_nl <= MUX_s_1_2_2(mux_1724_nl, nand_429_nl, fsm_output(5));
  or_1557_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1726 <= MUX_s_1_2_2(mux_1725_nl, or_1557_nl, fsm_output(4));
  or_1564_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1562_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1728 <= MUX_s_1_2_2(or_1564_nl, or_1562_nl, fsm_output(5));
  or_tmp_1580 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_1583 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1644_nl <= (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1643_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1642_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1781_nl <= MUX_s_1_2_2(or_1643_nl, or_1642_nl, fsm_output(0));
  mux_tmp_1782 <= MUX_s_1_2_2(or_1644_nl, mux_1781_nl, fsm_output(5));
  or_1652_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1651_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1785_nl <= MUX_s_1_2_2(or_1652_nl, or_1651_nl, fsm_output(0));
  nand_428_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1010"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_1786_nl <= MUX_s_1_2_2(mux_1785_nl, nand_428_nl, fsm_output(5));
  or_1648_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_tmp_1787 <= MUX_s_1_2_2(mux_1786_nl, or_1648_nl, fsm_output(4));
  or_1656_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1654_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1788 <= MUX_s_1_2_2(or_1656_nl, or_1654_nl, fsm_output(5));
  or_tmp_1691 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_1695 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1758_nl <= (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1757_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1756_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_1858_nl <= MUX_s_1_2_2(or_1757_nl, or_1756_nl, fsm_output(0));
  mux_tmp_1859 <= MUX_s_1_2_2(or_1758_nl, mux_1858_nl, fsm_output(5));
  or_1774_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1773_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_1868_nl <= MUX_s_1_2_2(or_1774_nl, or_1773_nl, fsm_output(0));
  nand_427_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_1869_nl <= MUX_s_1_2_2(mux_1868_nl, nand_427_nl, fsm_output(5));
  or_1770_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_1870 <= MUX_s_1_2_2(mux_1869_nl, or_1770_nl, fsm_output(4));
  nand_416_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  or_1775_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_1872 <= MUX_s_1_2_2(nand_416_nl, or_1775_nl, fsm_output(5));
  or_1853_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(10));
  or_1852_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)) OR (fsm_output(9)) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  mux_1922_nl <= MUX_s_1_2_2(or_1853_nl, or_1852_nl, fsm_output(0));
  or_tmp_1797 <= (fsm_output(5)) OR mux_1922_nl;
  not_tmp_378 <= NOT((fsm_output(6)) AND (fsm_output(10)));
  nor_874_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(4))) OR (fsm_output(9)) OR
      (fsm_output(3)) OR not_tmp_378);
  nor_875_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)) OR (NOT((fsm_output(9)) AND (fsm_output(3)) AND (fsm_output(6))
      AND (fsm_output(10)))));
  mux_1926_nl <= MUX_s_1_2_2(nor_874_nl, nor_875_nl, fsm_output(0));
  nand_73_nl <= NOT((fsm_output(5)) AND mux_1926_nl);
  or_1856_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(4)) OR (fsm_output(9)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_1855_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)) OR (NOT (fsm_output(9))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (fsm_output(10));
  mux_1925_nl <= MUX_s_1_2_2(or_1856_nl, or_1855_nl, fsm_output(0));
  or_1857_nl <= (fsm_output(5)) OR mux_1925_nl;
  mux_tmp_1927 <= MUX_s_1_2_2(nand_73_nl, or_1857_nl, fsm_output(8));
  nor_872_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(4)) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(10)));
  nor_873_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(4)) OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(10))));
  mux_1929_nl <= MUX_s_1_2_2(nor_872_nl, nor_873_nl, fsm_output(0));
  nand_tmp_74 <= NOT((fsm_output(5)) AND mux_1929_nl);
  or_tmp_1811 <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(4)))
      OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(10));
  or_tmp_1812 <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(4)) OR (NOT (fsm_output(9)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  not_tmp_381 <= NOT((fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(10)));
  or_tmp_1821 <= (fsm_output(4)) OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  or_tmp_1907 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_1911 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_1974_nl <= (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_1973_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1972_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_2003_nl <= MUX_s_1_2_2(or_1973_nl, or_1972_nl, fsm_output(0));
  mux_tmp_2004 <= MUX_s_1_2_2(or_1974_nl, mux_2003_nl, fsm_output(5));
  or_1990_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_1989_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_2013_nl <= MUX_s_1_2_2(or_1990_nl, or_1989_nl, fsm_output(0));
  nand_426_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_2014_nl <= MUX_s_1_2_2(mux_2013_nl, nand_426_nl, fsm_output(5));
  or_1986_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_2015 <= MUX_s_1_2_2(mux_2014_nl, or_1986_nl, fsm_output(4));
  nand_414_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  or_1991_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_2017 <= MUX_s_1_2_2(nand_414_nl, or_1991_nl, fsm_output(5));
  or_tmp_2009 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_2012 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_2073_nl <= (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_2072_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_2071_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_2070_nl <= MUX_s_1_2_2(or_2072_nl, or_2071_nl, fsm_output(0));
  mux_tmp_2071 <= MUX_s_1_2_2(or_2073_nl, mux_2070_nl, fsm_output(5));
  or_2081_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  or_2080_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(8))) OR (fsm_output(10));
  mux_2074_nl <= MUX_s_1_2_2(or_2081_nl, or_2080_nl, fsm_output(0));
  nand_425_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_2075_nl <= MUX_s_1_2_2(mux_2074_nl, nand_425_nl, fsm_output(5));
  or_2077_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR
      (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_tmp_2076 <= MUX_s_1_2_2(mux_2075_nl, or_2077_nl, fsm_output(4));
  nand_412_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  or_2083_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_2077 <= MUX_s_1_2_2(nand_412_nl, or_2083_nl, fsm_output(5));
  or_tmp_2120 <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_2124 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_2187_nl <= (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  nand_291_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (fsm_output(3)) AND (NOT (fsm_output(6)))
      AND (fsm_output(9)) AND (fsm_output(8)) AND (NOT (fsm_output(10))));
  or_2185_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_2147_nl <= MUX_s_1_2_2(nand_291_nl, or_2185_nl, fsm_output(0));
  mux_tmp_2148 <= MUX_s_1_2_2(or_2187_nl, mux_2147_nl, fsm_output(5));
  nand_288_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (VEC_LOOP_j_sva_11_0(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT
      (fsm_output(9))) AND (fsm_output(8)) AND (NOT (fsm_output(10))));
  nand_289_nl <= NOT((NOT (fsm_output(3))) AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(6)) AND (fsm_output(9))
      AND (fsm_output(8)) AND (NOT (fsm_output(10))));
  mux_2157_nl <= MUX_s_1_2_2(nand_288_nl, nand_289_nl, fsm_output(0));
  nand_424_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_2158_nl <= MUX_s_1_2_2(mux_2157_nl, nand_424_nl, fsm_output(5));
  or_2199_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_tmp_2159 <= MUX_s_1_2_2(mux_2158_nl, or_2199_nl, fsm_output(4));
  nand_410_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  or_2204_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(6)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_2161 <= MUX_s_1_2_2(nand_410_nl, or_2204_nl, fsm_output(5));
  and_dcpl_260 <= and_dcpl_124 AND and_dcpl_100 AND and_dcpl_98;
  nor_784_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  or_tmp_2220 <= nor_784_cse OR (NOT (fsm_output(3))) OR (fsm_output(10));
  or_tmp_2223 <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(10));
  or_tmp_2225 <= (NOT(and_573_cse OR (fsm_output(3)))) OR (fsm_output(10));
  or_tmp_2230 <= and_573_cse OR (fsm_output(3)) OR (fsm_output(10));
  or_tmp_2233 <= ((fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(1))) OR (fsm_output(10));
  mux_tmp_2218 <= MUX_s_1_2_2((NOT or_tmp_2233), or_tmp_21, fsm_output(6));
  mux_tmp_2220 <= MUX_s_1_2_2(and_dcpl_102, nor_tmp_6, fsm_output(6));
  mux_tmp_2223 <= MUX_s_1_2_2((NOT nor_tmp_9), or_tmp_2233, fsm_output(6));
  or_tmp_2237 <= NOT((fsm_output(6)) AND (fsm_output(1)) AND (fsm_output(3)) AND
      (NOT (fsm_output(10))));
  or_tmp_2238 <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(10));
  mux_tmp_2239 <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), fsm_output(3));
  mux_2240_nl <= MUX_s_1_2_2(and_dcpl_101, mux_tmp_2239, or_2348_cse);
  nand_tmp_92 <= NOT((fsm_output(6)) AND (NOT mux_2240_nl));
  nor_tmp_286 <= or_2898_cse AND (fsm_output(10));
  or_tmp_2246 <= (fsm_output(6)) OR (NOT (fsm_output(3))) OR (fsm_output(10));
  or_tmp_2248 <= (or_2348_cse AND (fsm_output(3))) OR (fsm_output(10));
  not_tmp_426 <= NOT((fsm_output(6)) AND or_tmp_2248);
  nor_tmp_288 <= ((fsm_output(3)) OR (fsm_output(1))) AND (fsm_output(10));
  and_tmp_10 <= (fsm_output(6)) AND nor_tmp_288;
  mux_tmp_2250 <= MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, or_2348_cse);
  mux_tmp_2251 <= MUX_s_1_2_2(and_dcpl_101, mux_tmp_2239, fsm_output(1));
  mux_tmp_2254 <= MUX_s_1_2_2(and_dcpl_101, mux_tmp_2239, and_573_cse);
  or_tmp_2253 <= ((fsm_output(3)) AND (fsm_output(1))) OR (fsm_output(10));
  or_tmp_2255 <= (fsm_output(6)) OR or_tmp_2253;
  mux_tmp_2265 <= MUX_s_1_2_2(and_dcpl_109, (fsm_output(10)), fsm_output(6));
  nor_tmp_291 <= or_2348_cse AND (fsm_output(3)) AND (fsm_output(10));
  or_tmp_2257 <= (fsm_output(6)) OR or_tmp_2248;
  nor_tmp_295 <= or_2902_cse AND (fsm_output(10));
  mux_tmp_2285 <= MUX_s_1_2_2((NOT nor_tmp_288), (fsm_output(10)), fsm_output(6));
  mux_2289_nl <= MUX_s_1_2_2(and_dcpl_101, or_tmp_2230, fsm_output(6));
  mux_tmp_2290 <= MUX_s_1_2_2(not_tmp_378, mux_2289_nl, fsm_output(7));
  or_tmp_2260 <= (fsm_output(3)) OR (NOT (fsm_output(10)));
  or_tmp_2263 <= (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  nand_tmp_93 <= NOT((fsm_output(6)) AND (NOT or_tmp_2230));
  or_tmp_2266 <= (fsm_output(1)) OR (NOT mux_tmp_2239);
  mux_tmp_2309 <= MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, fsm_output(1));
  mux_2310_nl <= MUX_s_1_2_2(mux_tmp_2309, (NOT or_tmp_2266), fsm_output(0));
  or_tmp_2267 <= (fsm_output(6)) OR mux_2310_nl;
  or_tmp_2269 <= (NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(3))))
      OR (fsm_output(10));
  nand_tmp_95 <= NOT((fsm_output(6)) AND (NOT or_tmp_2269));
  or_tmp_2271 <= (NOT((fsm_output(1)) OR (fsm_output(3)))) OR (fsm_output(10));
  nand_tmp_96 <= NOT((fsm_output(6)) AND (NOT or_tmp_2253));
  or_tmp_2275 <= (NOT((fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1)))) OR
      (fsm_output(10));
  or_tmp_2276 <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(10));
  or_tmp_2277 <= (fsm_output(0)) OR (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(10));
  mux_tmp_2327 <= MUX_s_1_2_2(or_tmp_2277, nor_tmp_291, fsm_output(6));
  or_tmp_2280 <= (fsm_output(6)) OR (NOT or_tmp_2220);
  or_tmp_2281 <= (fsm_output(6)) OR and_dcpl_110;
  or_tmp_2282 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(10));
  or_tmp_2289 <= nor_784_cse OR (fsm_output(3)) OR (NOT (fsm_output(10)));
  not_tmp_463 <= NOT((fsm_output(6)) AND or_tmp_2289);
  mux_tmp_2349 <= MUX_s_1_2_2((NOT or_tmp_2248), or_tmp_21, fsm_output(6));
  and_tmp_16 <= (fsm_output(6)) AND or_tmp_2282;
  or_tmp_2293 <= (fsm_output(6)) OR (NOT nor_tmp_295);
  mux_tmp_2362 <= MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, and_573_cse);
  nor_tmp_300 <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(3)) AND (fsm_output(10));
  or_tmp_2327 <= NOT((fsm_output(5)) AND (fsm_output(8)) AND (fsm_output(6)) AND
      (NOT (fsm_output(10))));
  or_tmp_2329 <= (fsm_output(5)) OR (fsm_output(8)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_tmp_2331 <= (fsm_output(5)) OR (fsm_output(8)) OR (NOT (fsm_output(6)));
  or_tmp_2333 <= (NOT (fsm_output(8))) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_tmp_2334 <= (NOT (fsm_output(8))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_tmp_2400 <= MUX_s_1_2_2(or_tmp_2334, or_tmp_2333, fsm_output(5));
  mux_tmp_2401 <= MUX_s_1_2_2(or_tmp_4, or_tmp_14, fsm_output(8));
  mux_tmp_2402 <= MUX_s_1_2_2(mux_tmp_2401, or_tmp_2333, fsm_output(5));
  or_tmp_2335 <= (fsm_output(5)) OR mux_tmp_2401;
  or_2393_nl <= (fsm_output(8)) OR not_tmp_378;
  mux_tmp_2406 <= MUX_s_1_2_2(or_2393_nl, or_tmp_2334, fsm_output(5));
  or_tmp_2338 <= (fsm_output(5)) OR (fsm_output(8)) OR not_tmp_378;
  nand_tmp_105 <= NOT((fsm_output(5)) AND (NOT mux_tmp_2401));
  mux_tmp_2423 <= MUX_s_1_2_2(or_tmp_2334, mux_tmp_917, fsm_output(5));
  nor_tmp_307 <= (fsm_output(8)) AND (fsm_output(6)) AND (fsm_output(10));
  mux_tmp_2425 <= MUX_s_1_2_2((NOT (fsm_output(6))), or_tmp_434, fsm_output(8));
  mux_tmp_2426 <= MUX_s_1_2_2((NOT mux_tmp_2425), nor_tmp_307, fsm_output(5));
  or_tmp_2342 <= (fsm_output(5)) OR mux_tmp_2425;
  mux_2427_nl <= MUX_s_1_2_2(not_tmp_378, or_tmp_434, fsm_output(8));
  or_tmp_2343 <= (fsm_output(5)) OR mux_2427_nl;
  mux_2433_itm <= MUX_s_1_2_2(or_tmp_4, (fsm_output(6)), fsm_output(8));
  mux_2435_itm <= MUX_s_1_2_2(or_tmp_4, or_tmp_434, fsm_output(8));
  mux_tmp_2436 <= MUX_s_1_2_2((NOT mux_2435_itm), nor_tmp_307, fsm_output(5));
  nand_tmp_107 <= NOT((fsm_output(5)) AND (NOT mux_2433_itm));
  nand_tmp_108 <= NOT((fsm_output(5)) AND (NOT mux_2435_itm));
  or_2415_cse <= (fsm_output(9)) OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  mux_tmp_2466 <= MUX_s_1_2_2(or_tmp_195, or_2415_cse, fsm_output(1));
  or_2409_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(1))) OR (fsm_output(9))
      OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_2463_cse <= MUX_s_1_2_2(or_2409_nl, or_2824_cse, fsm_output(0));
  or_2425_nl <= (fsm_output(5)) OR (fsm_output(2)) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (fsm_output(4)) OR (fsm_output(10));
  or_2424_nl <= (fsm_output(2)) OR (fsm_output(0)) OR nand_226_cse;
  mux_2470_nl <= MUX_s_1_2_2(or_529_cse, or_2826_cse, fsm_output(0));
  mux_2471_nl <= MUX_s_1_2_2(mux_2470_nl, or_2839_cse, fsm_output(2));
  mux_2472_nl <= MUX_s_1_2_2(or_2424_nl, mux_2471_nl, fsm_output(5));
  mux_2473_nl <= MUX_s_1_2_2(or_2425_nl, mux_2472_nl, fsm_output(6));
  or_2419_nl <= (fsm_output(3)) OR mux_tmp_2466;
  mux_2469_nl <= MUX_s_1_2_2(or_2419_nl, or_529_cse, fsm_output(0));
  or_3285_nl <= (NOT (fsm_output(6))) OR (fsm_output(5)) OR (NOT (fsm_output(2)))
      OR mux_2469_nl;
  mux_2474_nl <= MUX_s_1_2_2(mux_2473_nl, or_3285_nl, fsm_output(7));
  nand_111_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_2466));
  mux_2467_nl <= MUX_s_1_2_2(or_2824_cse, nand_111_nl, fsm_output(0));
  or_2417_nl <= (fsm_output(6)) OR (NOT (fsm_output(5))) OR (fsm_output(2)) OR mux_2467_nl;
  mux_2464_nl <= MUX_s_1_2_2(or_2819_cse, mux_2463_cse, fsm_output(2));
  or_2412_nl <= (fsm_output(5)) OR mux_2464_nl;
  nor_756_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(1)) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_757_nl <= NOT((fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(9)) OR nand_398_cse);
  mux_2462_nl <= MUX_s_1_2_2(nor_756_nl, nor_757_nl, fsm_output(0));
  nand_110_nl <= NOT((fsm_output(5)) AND (fsm_output(2)) AND mux_2462_nl);
  mux_2465_nl <= MUX_s_1_2_2(or_2412_nl, nand_110_nl, fsm_output(6));
  mux_2468_nl <= MUX_s_1_2_2(or_2417_nl, mux_2465_nl, fsm_output(7));
  mux_2475_itm <= MUX_s_1_2_2(mux_2474_nl, mux_2468_nl, fsm_output(8));
  nor_743_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_744_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(4)) OR (fsm_output(10)));
  mux_2486_nl <= MUX_s_1_2_2(nor_743_nl, nor_744_nl, fsm_output(5));
  or_3233_nl <= (NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  or_3232_nl <= (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_34;
  mux_3706_nl <= MUX_s_1_2_2(or_3233_nl, or_3232_nl, fsm_output(2));
  nor_745_nl <= NOT((fsm_output(5)) OR mux_3706_nl);
  mux_2487_nl <= MUX_s_1_2_2(mux_2486_nl, nor_745_nl, fsm_output(6));
  or_2441_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  or_2439_nl <= (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(8)) OR nand_398_cse;
  mux_2483_nl <= MUX_s_1_2_2(or_2441_nl, or_2439_nl, fsm_output(2));
  nor_746_nl <= NOT((fsm_output(5)) OR mux_2483_nl);
  nor_1285_nl <= NOT((fsm_output(7)) OR (fsm_output(3)) OR (NOT (fsm_output(8)))
      OR (fsm_output(4)) OR (fsm_output(9)) OR (fsm_output(10)));
  nor_1286_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(8))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (fsm_output(10)));
  mux_89_nl <= MUX_s_1_2_2(nor_1285_nl, nor_1286_nl, fsm_output(2));
  and_558_nl <= (fsm_output(5)) AND mux_89_nl;
  mux_2484_nl <= MUX_s_1_2_2(nor_746_nl, and_558_nl, fsm_output(6));
  mux_2488_nl <= MUX_s_1_2_2(mux_2487_nl, mux_2484_nl, fsm_output(1));
  nor_750_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_34);
  nor_1278_nl <= NOT((fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(4))
      OR (fsm_output(9)) OR (NOT (fsm_output(10))));
  mux_2478_nl <= MUX_s_1_2_2(nor_750_nl, nor_1278_nl, fsm_output(2));
  mux_2479_nl <= MUX_s_1_2_2(nor_1276_cse, mux_2478_nl, fsm_output(5));
  mux_2480_nl <= MUX_s_1_2_2(mux_2479_nl, nor_1279_cse, fsm_output(6));
  nor_1280_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(8)))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (fsm_output(10)));
  nor_1281_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(3)) OR (NOT (fsm_output(8)))
      OR (fsm_output(4)) OR (fsm_output(9)) OR (fsm_output(10)));
  mux_93_nl <= MUX_s_1_2_2(nor_1280_nl, nor_1281_nl, fsm_output(2));
  mux_94_nl <= MUX_s_1_2_2(mux_93_nl, nor_544_cse, fsm_output(5));
  and_796_nl <= (fsm_output(6)) AND mux_94_nl;
  mux_2481_nl <= MUX_s_1_2_2(mux_2480_nl, and_796_nl, fsm_output(1));
  not_tmp_519 <= MUX_s_1_2_2(mux_2488_nl, mux_2481_nl, fsm_output(0));
  and_dcpl_264 <= NOT((fsm_output(10)) OR (fsm_output(6)));
  mux_2490_nl <= MUX_s_1_2_2((NOT (fsm_output(3))), (fsm_output(3)), fsm_output(1));
  or_463_nl <= (NOT (fsm_output(1))) OR (fsm_output(3));
  mux_2491_nl <= MUX_s_1_2_2(mux_2490_nl, or_463_nl, fsm_output(0));
  mux_2492_nl <= MUX_s_1_2_2(mux_2491_nl, (fsm_output(3)), fsm_output(2));
  and_dcpl_266 <= (NOT mux_2492_nl) AND and_dcpl_264 AND (NOT (fsm_output(7))) AND
      (NOT (fsm_output(5))) AND (NOT (fsm_output(8))) AND and_dcpl;
  and_dcpl_268 <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  nor_741_nl <= NOT((fsm_output(5)) OR (NOT((fsm_output(0)) AND (fsm_output(3)))));
  nor_742_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(3)));
  mux_2496_nl <= MUX_s_1_2_2(nor_741_nl, nor_742_nl, fsm_output(4));
  and_dcpl_273 <= mux_2496_nl AND and_dcpl_26 AND and_dcpl_268 AND (NOT (fsm_output(2)))
      AND nor_610_cse;
  mux_tmp_2502 <= MUX_s_1_2_2(and_dcpl_101, mux_tmp_2239, fsm_output(2));
  not_tmp_529 <= NOT(and_459_cse OR (fsm_output(10)));
  nor_tmp_330 <= (and_573_cse OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")))
      AND (fsm_output(10));
  or_2468_nl <= (or_2385_cse AND (fsm_output(3))) OR (fsm_output(10));
  mux_tmp_2508 <= MUX_s_1_2_2(nor_tmp_330, or_2468_nl, fsm_output(9));
  or_tmp_2416 <= and_458_cse OR (fsm_output(10));
  or_tmp_2419 <= and_440_cse OR (fsm_output(10));
  mux_tmp_2519 <= MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, fsm_output(2));
  mux_tmp_2523 <= MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, fsm_output(2));
  mux_tmp_2525 <= MUX_s_1_2_2(mux_tmp_2502, mux_tmp_2519, fsm_output(1));
  nor_tmp_338 <= or_2894_cse AND (fsm_output(10));
  or_3280_cse <= and_573_cse OR (fsm_output(2));
  or_tmp_2429 <= (or_3280_cse AND (fsm_output(3))) OR (fsm_output(10));
  or_3279_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  nor_tmp_342 <= or_3279_cse AND (fsm_output(10));
  or_2489_nl <= (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(10));
  mux_tmp_2549 <= MUX_s_1_2_2(or_tmp_2429, or_2489_nl, fsm_output(9));
  mux_tmp_2650 <= MUX_s_1_2_2(nor_601_cse, and_816_cse, fsm_output(7));
  and_dcpl_279 <= and_dcpl_40 AND and_dcpl_30;
  and_dcpl_281 <= and_dcpl_103 AND and_dcpl_116;
  mux_tmp_2687 <= MUX_s_1_2_2((NOT and_dcpl_240), nor_tmp_6, fsm_output(6));
  or_tmp_2474 <= (fsm_output(6)) OR or_tmp_2275;
  mux_tmp_2696 <= MUX_s_1_2_2(and_dcpl_101, or_tmp_21, fsm_output(6));
  nand_117_nl <= NOT((fsm_output(6)) AND (NOT or_tmp_2248));
  mux_tmp_2698 <= MUX_s_1_2_2((NOT (fsm_output(6))), nand_117_nl, fsm_output(7));
  nor_719_nl <= NOT((fsm_output(6)) OR (NOT or_tmp_2230));
  mux_tmp_2701 <= MUX_s_1_2_2(nor_719_nl, or_tmp_4, fsm_output(7));
  or_tmp_2479 <= (fsm_output(6)) OR and_dcpl_101;
  nand_tmp_119 <= NOT((fsm_output(6)) AND (NOT nor_tmp_300));
  or_tmp_2483 <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3)) OR (NOT (fsm_output(10)));
  and_dcpl_283 <= and_dcpl_128 AND and_dcpl_100 AND and_dcpl_116;
  and_dcpl_305 <= and_dcpl_2 AND and_dcpl;
  or_2556_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(4))
      OR (fsm_output(10));
  or_2555_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_2746_cse <= MUX_s_1_2_2(or_2556_nl, or_2555_nl, fsm_output(2));
  nor_702_nl <= NOT((fsm_output(1)) OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR
      (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_704_nl <= NOT((fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  mux_2753_nl <= MUX_s_1_2_2(nor_539_cse, nor_704_nl, fsm_output(1));
  mux_2754_nl <= MUX_s_1_2_2(nor_702_nl, mux_2753_nl, fsm_output(5));
  nor_705_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(7))) OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(4))
      OR (fsm_output(10)));
  mux_2755_nl <= MUX_s_1_2_2(mux_2754_nl, nor_705_nl, fsm_output(6));
  nor_706_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(1)) OR (fsm_output(2)) OR
      (NOT (fsm_output(7))) OR (fsm_output(9)) OR not_tmp_34);
  nor_707_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(7)) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(4))) OR
      (fsm_output(10)));
  nor_708_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_1296_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  mux_2750_nl <= MUX_s_1_2_2(nor_708_nl, nor_1296_nl, fsm_output(1));
  mux_2751_nl <= MUX_s_1_2_2(nor_707_nl, mux_2750_nl, fsm_output(5));
  mux_2752_nl <= MUX_s_1_2_2(nor_706_nl, mux_2751_nl, fsm_output(6));
  mux_2756_nl <= MUX_s_1_2_2(mux_2755_nl, mux_2752_nl, fsm_output(3));
  nor_710_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(4)))
      OR (fsm_output(10)));
  nor_711_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(7)) OR
      (fsm_output(9)) OR not_tmp_34);
  nor_712_nl <= NOT((fsm_output(1)) OR mux_2746_cse);
  mux_2747_nl <= MUX_s_1_2_2(nor_711_nl, nor_712_nl, fsm_output(5));
  mux_2748_nl <= MUX_s_1_2_2(nor_710_nl, mux_2747_nl, fsm_output(6));
  or_53_nl <= (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(4))
      OR (NOT (fsm_output(10)));
  or_51_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 7)/=STD_LOGIC_VECTOR'("100")) OR nand_398_cse;
  mux_74_nl <= MUX_s_1_2_2(or_53_nl, or_51_nl, fsm_output(2));
  or_2553_nl <= (fsm_output(1)) OR mux_74_nl;
  nand_120_nl <= NOT((fsm_output(1)) AND mux_71_cse);
  mux_2745_nl <= MUX_s_1_2_2(or_2553_nl, nand_120_nl, fsm_output(5));
  nor_713_nl <= NOT((fsm_output(6)) OR mux_2745_nl);
  mux_2749_nl <= MUX_s_1_2_2(mux_2748_nl, nor_713_nl, fsm_output(3));
  not_tmp_596 <= MUX_s_1_2_2(mux_2756_nl, mux_2749_nl, fsm_output(0));
  or_tmp_2516 <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(4)) OR (fsm_output(10));
  or_2578_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR nand_398_cse;
  mux_tmp_2758 <= MUX_s_1_2_2(or_2578_nl, or_tmp_2516, fsm_output(9));
  mux_tmp_2788 <= MUX_s_1_2_2(or_tmp_2238, (fsm_output(10)), fsm_output(6));
  mux_tmp_2790 <= MUX_s_1_2_2(or_tmp_21, or_tmp_237, fsm_output(6));
  or_2621_nl <= (fsm_output(0)) OR (NOT and_dcpl_240);
  mux_tmp_2796 <= MUX_s_1_2_2(or_2621_nl, mux_tmp_2309, fsm_output(6));
  mux_2799_nl <= MUX_s_1_2_2(nor_tmp_6, mux_tmp_2239, fsm_output(1));
  mux_tmp_2800 <= MUX_s_1_2_2(and_dcpl_240, mux_2799_nl, fsm_output(0));
  mux_tmp_2813 <= MUX_s_1_2_2(or_tmp_2277, or_tmp_2230, fsm_output(6));
  or_207_nl <= (fsm_output(4)) OR (NOT (fsm_output(10)));
  mux_2871_nl <= MUX_s_1_2_2(or_tmp_178, or_207_nl, fsm_output(1));
  or_tmp_2594 <= (fsm_output(3)) OR (fsm_output(9)) OR mux_2871_nl;
  nor_672_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR
      nand_398_cse);
  nor_673_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR
      nand_398_cse);
  mux_2878_nl <= MUX_s_1_2_2(nor_672_nl, nor_673_nl, fsm_output(0));
  mux_2879_nl <= MUX_s_1_2_2(mux_2878_nl, and_464_cse, fsm_output(2));
  and_503_nl <= (NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01"))))
      AND mux_2879_nl;
  or_2662_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR nand_398_cse;
  or_2659_nl <= (fsm_output(0)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(1))
      OR (fsm_output(4)) OR (fsm_output(10));
  mux_2876_nl <= MUX_s_1_2_2(or_2839_cse, or_2659_nl, fsm_output(2));
  mux_2877_nl <= MUX_s_1_2_2(or_2662_nl, mux_2876_nl, fsm_output(5));
  nor_674_nl <= NOT((fsm_output(6)) OR mux_2877_nl);
  mux_2880_nl <= MUX_s_1_2_2(and_503_nl, nor_674_nl, fsm_output(7));
  mux_2873_nl <= MUX_s_1_2_2(or_tmp_2594, or_529_cse, fsm_output(0));
  nor_675_nl <= NOT((fsm_output(5)) OR (fsm_output(2)) OR mux_2873_nl);
  mux_2872_nl <= MUX_s_1_2_2(or_525_cse, or_tmp_2594, fsm_output(0));
  and_505_nl <= (fsm_output(5)) AND (fsm_output(2)) AND (NOT mux_2872_nl);
  mux_2874_nl <= MUX_s_1_2_2(nor_675_nl, and_505_nl, fsm_output(6));
  or_2647_nl <= (fsm_output(0)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  mux_2870_nl <= MUX_s_1_2_2(mux_2463_cse, or_2647_nl, fsm_output(2));
  nor_676_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10"))
      OR mux_2870_nl);
  mux_2875_nl <= MUX_s_1_2_2(mux_2874_nl, nor_676_nl, fsm_output(7));
  not_tmp_634 <= MUX_s_1_2_2(mux_2880_nl, mux_2875_nl, fsm_output(8));
  or_tmp_2631 <= (fsm_output(2)) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(7)))
      OR (fsm_output(4)) OR (fsm_output(10));
  nor_654_nl <= NOT((NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(8))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  nor_655_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(8)) OR (fsm_output(7)) OR
      (fsm_output(4)) OR (fsm_output(10)));
  nor_656_nl <= NOT((fsm_output(2)) OR (fsm_output(8)) OR (fsm_output(7)) OR (NOT
      (fsm_output(4))) OR (fsm_output(10)));
  mux_2899_nl <= MUX_s_1_2_2(nor_655_nl, nor_656_nl, fsm_output(9));
  mux_2900_nl <= MUX_s_1_2_2(nor_654_nl, mux_2899_nl, fsm_output(1));
  and_498_nl <= (fsm_output(6)) AND mux_2900_nl;
  nor_657_nl <= NOT((fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(8))
      OR nand_240_cse);
  and_499_nl <= (fsm_output(1)) AND (fsm_output(9)) AND (fsm_output(2)) AND (fsm_output(8))
      AND (fsm_output(7)) AND (NOT (fsm_output(4))) AND (NOT (fsm_output(10)));
  mux_2898_nl <= MUX_s_1_2_2(nor_657_nl, and_499_nl, fsm_output(6));
  mux_2901_nl <= MUX_s_1_2_2(and_498_nl, mux_2898_nl, fsm_output(5));
  or_2699_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (fsm_output(7))
      OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_2896_nl <= MUX_s_1_2_2(or_tmp_2631, or_2699_nl, fsm_output(9));
  nor_658_nl <= NOT((fsm_output(6)) OR (fsm_output(1)) OR mux_2896_nl);
  nor_659_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(9)) OR (NOT (fsm_output(2)))
      OR (fsm_output(8)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_660_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(2)) OR
      (NOT (fsm_output(8))) OR (fsm_output(7)) OR nand_398_cse);
  mux_2895_nl <= MUX_s_1_2_2(nor_659_nl, nor_660_nl, fsm_output(6));
  mux_2897_nl <= MUX_s_1_2_2(nor_658_nl, mux_2895_nl, fsm_output(5));
  mux_2902_nl <= MUX_s_1_2_2(mux_2901_nl, mux_2897_nl, fsm_output(3));
  or_2693_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (fsm_output(7))
      OR nand_398_cse;
  mux_2892_nl <= MUX_s_1_2_2(or_2693_nl, or_tmp_2631, fsm_output(9));
  nor_661_nl <= NOT((fsm_output(6)) OR (fsm_output(1)) OR mux_2892_nl);
  nor_662_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(8))) OR (fsm_output(7)) OR
      (fsm_output(4)) OR (fsm_output(10)));
  nor_663_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(8)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  mux_2891_nl <= MUX_s_1_2_2(nor_662_nl, nor_663_nl, fsm_output(9));
  and_500_nl <= (NOT((fsm_output(6)) OR (NOT (fsm_output(1))))) AND mux_2891_nl;
  mux_2893_nl <= MUX_s_1_2_2(nor_661_nl, and_500_nl, fsm_output(5));
  nor_664_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(1))) OR (fsm_output(9))
      OR mux_3498_cse);
  nor_665_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(1)) OR (fsm_output(9)) OR
      (NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(7))) OR
      (fsm_output(4)) OR (fsm_output(10)));
  mux_2890_nl <= MUX_s_1_2_2(nor_664_nl, nor_665_nl, fsm_output(5));
  mux_2894_nl <= MUX_s_1_2_2(mux_2893_nl, mux_2890_nl, fsm_output(3));
  not_tmp_646 <= MUX_s_1_2_2(mux_2902_nl, mux_2894_nl, fsm_output(0));
  or_248_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 9)/=STD_LOGIC_VECTOR'("10"));
  mux_523_nl <= MUX_s_1_2_2(or_248_nl, and_816_cse, fsm_output(4));
  or_tmp_2649 <= (fsm_output(8)) OR mux_523_nl;
  nand_tmp_136 <= (fsm_output(8)) OR (NOT (fsm_output(4))) OR and_816_cse;
  mux_tmp_2905 <= MUX_s_1_2_2(nand_tmp_136, or_tmp_2649, fsm_output(1));
  nand_tmp_137 <= NOT((fsm_output(4)) AND (NOT mux_726_cse));
  mux_tmp_2907 <= MUX_s_1_2_2(nand_tmp_137, or_tmp_182, fsm_output(8));
  or_tmp_2652 <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(10)));
  or_tmp_2653 <= (fsm_output(4)) OR and_816_cse;
  mux_tmp_2911 <= MUX_s_1_2_2(and_816_cse, or_tmp_187, fsm_output(4));
  mux_tmp_2912 <= MUX_s_1_2_2(mux_tmp_2911, or_tmp_2652, fsm_output(8));
  mux_2910_nl <= MUX_s_1_2_2(or_tmp_2653, or_tmp_2652, fsm_output(8));
  mux_tmp_2913 <= MUX_s_1_2_2(mux_tmp_2912, mux_2910_nl, fsm_output(1));
  mux_tmp_2919 <= MUX_s_1_2_2(or_tmp_179, nand_tmp_137, fsm_output(8));
  mux_2920_nl <= MUX_s_1_2_2(or_tmp_187, (NOT and_816_cse), fsm_output(4));
  mux_tmp_2921 <= MUX_s_1_2_2(mux_2920_nl, mux_tmp_2911, fsm_output(8));
  mux_tmp_2930 <= MUX_s_1_2_2(or_tmp_2652, or_tmp_179, fsm_output(8));
  or_tmp_2659 <= (fsm_output(8)) OR mux_tmp_2911;
  or_tmp_2663 <= (fsm_output(8)) OR (NOT or_tmp_2653);
  mux_520_nl <= MUX_s_1_2_2(mux_726_cse, and_816_cse, fsm_output(4));
  nand_tmp_140 <= NOT((fsm_output(8)) AND (NOT mux_520_nl));
  or_tmp_2707 <= (fsm_output(7)) OR (NOT((fsm_output(2)) AND (fsm_output(4)) AND
      (fsm_output(10))));
  and_dcpl_332 <= and_dcpl_128 AND and_dcpl_117 AND and_dcpl_116;
  nor_627_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_628_nl <= NOT((fsm_output(9)) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  mux_3168_nl <= MUX_s_1_2_2(nor_627_nl, nor_628_nl, fsm_output(1));
  nand_tmp_148 <= NOT((fsm_output(3)) AND mux_3168_nl);
  or_2886_nl <= (or_2894_cse AND (fsm_output(4))) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("000"));
  mux_3213_nl <= MUX_s_1_2_2(or_2951_cse, or_2886_nl, fsm_output(5));
  or_3260_nl <= (fsm_output(10)) OR mux_3213_nl;
  or_2882_nl <= (or_2348_cse AND (fsm_output(4))) OR CONV_SL_1_1(fsm_output(8 DOWNTO
      6)/=STD_LOGIC_VECTOR'("000"));
  mux_3212_nl <= MUX_s_1_2_2(or_2951_cse, or_2882_nl, and_459_cse);
  nand_220_nl <= NOT((fsm_output(10)) AND ((fsm_output(5)) OR mux_3212_nl));
  not_tmp_708 <= MUX_s_1_2_2(or_3260_nl, nand_220_nl, fsm_output(9));
  nor_tmp_445 <= or_2935_cse AND (fsm_output(9));
  mux_tmp_3219 <= MUX_s_1_2_2((NOT (fsm_output(9))), (fsm_output(9)), or_2935_cse);
  or_2905_nl <= (fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3));
  mux_3235_nl <= MUX_s_1_2_2(or_2520_cse, or_2905_nl, fsm_output(5));
  or_2904_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_3236 <= MUX_s_1_2_2(mux_3235_nl, or_2904_nl, fsm_output(2));
  or_tmp_2849 <= nor_1316_cse OR (fsm_output(9));
  mux_tmp_3244 <= MUX_s_1_2_2((NOT (fsm_output(9))), (fsm_output(9)), or_2951_cse);
  nor_tmp_456 <= CONV_SL_1_1(fsm_output(9 DOWNTO 7)=STD_LOGIC_VECTOR'("111"));
  mux_tmp_3256 <= MUX_s_1_2_2(nor_610_cse, nor_tmp_116, fsm_output(7));
  not_tmp_728 <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 7)/=STD_LOGIC_VECTOR'("000")));
  or_tmp_2864 <= (NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 6)/=STD_LOGIC_VECTOR'("0000"))))
      OR (fsm_output(10));
  mux_tmp_3269 <= MUX_s_1_2_2(and_dcpl_264, (fsm_output(10)), fsm_output(7));
  nor_tmp_461 <= (and_450_cse OR CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00")))
      AND (fsm_output(10));
  mux_3279_nl <= MUX_s_1_2_2(mux_tmp_741, and_754_cse, fsm_output(7));
  and_436_nl <= (CONV_SL_1_1(fsm_output(9 DOWNTO 7)/=STD_LOGIC_VECTOR'("000"))) AND
      (fsm_output(10));
  mux_tmp_3280 <= MUX_s_1_2_2(mux_3279_nl, and_436_nl, fsm_output(6));
  mux_tmp_3281 <= MUX_s_1_2_2(mux_tmp_741, and_754_cse, or_2520_cse);
  nand_tmp_157 <= NOT((fsm_output(8)) AND nand_376_cse);
  mux_tmp_3323 <= MUX_s_1_2_2(or_tmp_179, mux_tmp_374, fsm_output(8));
  mux_3350_nl <= MUX_s_1_2_2(mux_tmp_381, mux_tmp_3323, fsm_output(1));
  mux_3351_nl <= MUX_s_1_2_2(mux_382_cse, mux_3350_nl, fsm_output(0));
  mux_3352_nl <= MUX_s_1_2_2(nand_tmp_12, mux_3351_nl, fsm_output(6));
  mux_3353_nl <= MUX_s_1_2_2(mux_3352_nl, mux_3557_cse, fsm_output(5));
  mux_3354_nl <= MUX_s_1_2_2(mux_3353_nl, mux_3555_cse, fsm_output(7));
  mux_3368_nl <= MUX_s_1_2_2(mux_3575_cse, mux_3354_nl, fsm_output(3));
  mux_3369_itm <= MUX_s_1_2_2(mux_3368_nl, mux_3551_cse, fsm_output(2));
  mux_3380_nl <= MUX_s_1_2_2(nor_1276_cse, mux_3603_cse, fsm_output(5));
  mux_3381_nl <= MUX_s_1_2_2(mux_3380_nl, nor_1279_cse, fsm_output(6));
  nor_591_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10)));
  nor_1295_nl <= NOT((fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  mux_3377_nl <= MUX_s_1_2_2(nor_591_nl, nor_1295_nl, fsm_output(3));
  mux_3378_nl <= MUX_s_1_2_2(mux_3377_nl, nor_544_cse, fsm_output(5));
  and_417_nl <= (fsm_output(6)) AND mux_3378_nl;
  mux_3382_nl <= MUX_s_1_2_2(mux_3381_nl, and_417_nl, fsm_output(1));
  nor_594_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(8)) OR
      (fsm_output(4)) OR (NOT (fsm_output(10))));
  nor_595_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 7)/=STD_LOGIC_VECTOR'("100"))
      OR nand_398_cse);
  mux_3374_nl <= MUX_s_1_2_2(nor_594_nl, nor_595_nl, fsm_output(2));
  and_418_nl <= nor_515_cse AND mux_3374_nl;
  nor_596_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(3)) OR mux_2746_cse);
  mux_3375_nl <= MUX_s_1_2_2(and_418_nl, nor_596_nl, fsm_output(6));
  nor_1287_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(9)) OR (fsm_output(10)));
  and_419_nl <= (fsm_output(3)) AND mux_71_cse;
  mux_3371_nl <= MUX_s_1_2_2(nor_1287_nl, and_419_nl, fsm_output(5));
  mux_3372_nl <= MUX_s_1_2_2(mux_3371_nl, nor_545_cse, fsm_output(6));
  mux_3376_nl <= MUX_s_1_2_2(mux_3375_nl, mux_3372_nl, fsm_output(1));
  not_tmp_762 <= MUX_s_1_2_2(mux_3382_nl, mux_3376_nl, fsm_output(0));
  or_3007_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  or_3006_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_tmp_3386 <= MUX_s_1_2_2(or_3007_nl, or_3006_nl, fsm_output(5));
  mux_3406_nl <= MUX_s_1_2_2(or_tmp_178, or_tmp_179, fsm_output(8));
  or_3037_nl <= (NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(7)) OR mux_3406_nl;
  mux_3407_nl <= MUX_s_1_2_2(or_3016_cse, or_3037_nl, fsm_output(5));
  mux_3408_nl <= MUX_s_1_2_2(or_3018_cse, mux_3407_nl, fsm_output(0));
  nor_573_nl <= NOT((fsm_output(6)) OR mux_3408_nl);
  mux_3409_nl <= MUX_s_1_2_2(nor_573_nl, mux_3392_cse, fsm_output(3));
  not_tmp_776 <= MUX_s_1_2_2(mux_3409_nl, mux_3388_cse, fsm_output(9));
  mux_tmp_3418 <= MUX_s_1_2_2(or_tmp_118, or_154_cse, fsm_output(5));
  mux_3421_nl <= MUX_s_1_2_2(or_tmp_179, or_tmp_178, fsm_output(8));
  mux_tmp_3422 <= MUX_s_1_2_2(mux_3421_nl, or_tmp_118, fsm_output(5));
  mux_tmp_3426 <= MUX_s_1_2_2((NOT and_491_cse), or_tmp_179, fsm_output(8));
  mux_tmp_3430 <= MUX_s_1_2_2(or_tmp_118, or_tmp_191, fsm_output(5));
  mux_tmp_3436 <= MUX_s_1_2_2(or_154_cse, or_tmp_110, fsm_output(5));
  nand_tmp_167 <= NOT((fsm_output(8)) AND (NOT and_491_cse));
  mux_tmp_3449 <= MUX_s_1_2_2(nand_tmp_167, or_tmp_191, fsm_output(5));
  mux_tmp_3450 <= MUX_s_1_2_2((NOT (fsm_output(8))), or_tmp_150, fsm_output(5));
  mux_tmp_3452 <= MUX_s_1_2_2((NOT (fsm_output(8))), mux_tmp_3426, fsm_output(5));
  mux_tmp_3456 <= MUX_s_1_2_2((NOT (fsm_output(4))), and_491_cse, fsm_output(8));
  mux_tmp_3458 <= MUX_s_1_2_2((NOT and_491_cse), and_491_cse, fsm_output(8));
  mux_tmp_3459 <= MUX_s_1_2_2((NOT or_tmp_191), mux_tmp_3458, fsm_output(5));
  mux_tmp_3467 <= MUX_s_1_2_2(not_tmp_34, nand_tmp_167, fsm_output(5));
  nor_568_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(10))));
  mux_tmp_3468 <= MUX_s_1_2_2(nor_568_nl, and_491_cse, fsm_output(8));
  mux_tmp_3471 <= MUX_s_1_2_2(mux_tmp_3468, (fsm_output(8)), fsm_output(5));
  and_tmp_36 <= (fsm_output(8)) AND or_tmp_179;
  or_tmp_3025 <= (fsm_output(6)) OR (fsm_output(5)) OR (NOT (fsm_output(3))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  mux_3613_nl <= MUX_s_1_2_2(and_dcpl_109, (fsm_output(10)), fsm_output(1));
  or_tmp_3107 <= (fsm_output(6)) OR (NOT mux_3613_nl);
  STAGE_LOOP_i_3_0_sva_mx0c1 <= and_dcpl_111 AND and_dcpl_106;
  and_540_cse <= or_2348_cse AND (fsm_output(2));
  nor_738_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  VEC_LOOP_j_sva_11_0_mx0c1 <= and_dcpl_110 AND and_dcpl_127 AND and_dcpl_106;
  nor_724_nl <= NOT((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(10)));
  mux_2662_nl <= MUX_s_1_2_2(nor_601_cse, nor_724_nl, fsm_output(3));
  and_521_nl <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(9)) AND (fsm_output(10));
  mux_2661_nl <= MUX_s_1_2_2(and_521_nl, and_816_cse, or_3279_cse);
  mux_2663_nl <= MUX_s_1_2_2(mux_2662_nl, mux_2661_nl, fsm_output(7));
  or_2522_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("000"));
  mux_2664_nl <= MUX_s_1_2_2(mux_2663_nl, and_815_cse, or_2522_nl);
  modExp_result_sva_mx0c0 <= MUX_s_1_2_2(mux_2664_nl, and_816_cse, fsm_output(8));
  STAGE_LOOP_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(STAGE_LOOP_i_3_0_sva_2(3
      DOWNTO 1)) + SIGNED'( "011"), 3));
  STAGE_LOOP_acc_itm_2_1 <= STAGE_LOOP_acc_nl(2);
  and_305_m1c <= and_dcpl_128 AND and_dcpl_108 AND and_dcpl_279;
  and_307_m1c <= and_dcpl_156 AND and_dcpl_162 AND and_dcpl_139;
  and_309_m1c <= and_dcpl_102 AND and_dcpl_173 AND and_dcpl_245;
  and_312_m1c <= and_dcpl_128 AND and_dcpl_162 AND and_dcpl_22 AND and_dcpl;
  and_315_m1c <= and_dcpl_124 AND and_dcpl_117 AND and_dcpl_46 AND and_dcpl_50;
  and_317_m1c <= and_dcpl_102 AND and_dcpl_127 AND and_dcpl_172;
  and_320_m1c <= and_dcpl_102 AND and_dcpl_204 AND and_dcpl_2 AND and_472_cse;
  and_322_m1c <= and_dcpl_125 AND and_dcpl_154 AND and_472_cse;
  and_324_m1c <= and_dcpl_140 AND and_dcpl_145 AND and_472_cse;
  and_327_m1c <= and_dcpl_223 AND and_dcpl_100 AND and_dcpl_305;
  and_329_m1c <= and_dcpl_215 AND and_dcpl_108 AND and_dcpl_98;
  and_331_m1c <= and_dcpl_240 AND and_dcpl_162 AND and_dcpl_305;
  and_334_m1c <= and_dcpl_110 AND and_dcpl_173 AND and_dcpl_154 AND and_dcpl_30;
  and_336_m1c <= and_dcpl_215 AND and_dcpl_127 AND and_dcpl_239;
  and_339_m1c <= and_dcpl_215 AND and_dcpl_117 AND and_dcpl_40 AND and_472_cse;
  and_139_nl <= and_dcpl_129 AND and_dcpl_98;
  or_533_nl <= (fsm_output(2)) OR (NOT((fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(9))
      AND (fsm_output(3)) AND (fsm_output(4)) AND (fsm_output(10))));
  or_531_nl <= (NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(4))
      OR (NOT (fsm_output(10)));
  mux_1041_nl <= MUX_s_1_2_2(or_531_nl, or_529_cse, fsm_output(0));
  or_532_nl <= (fsm_output(2)) OR mux_1041_nl;
  mux_1042_nl <= MUX_s_1_2_2(or_533_nl, or_532_nl, fsm_output(5));
  nor_1194_nl <= NOT((fsm_output(6)) OR mux_1042_nl);
  or_527_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (NOT (fsm_output(9))) OR (fsm_output(3))
      OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  or_524_nl <= (fsm_output(9)) OR (fsm_output(3)) OR (NOT (fsm_output(4))) OR (fsm_output(10));
  or_523_nl <= (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  mux_1037_nl <= MUX_s_1_2_2(or_524_nl, or_523_nl, fsm_output(1));
  mux_1038_nl <= MUX_s_1_2_2(or_525_cse, mux_1037_nl, fsm_output(0));
  mux_1039_nl <= MUX_s_1_2_2(or_527_nl, mux_1038_nl, fsm_output(2));
  nor_1195_nl <= NOT((fsm_output(5)) OR mux_1039_nl);
  nor_1196_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(9)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_1197_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (fsm_output(3))
      OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  mux_1035_nl <= MUX_s_1_2_2(nor_1196_nl, nor_1197_nl, fsm_output(0));
  nor_1198_nl <= NOT((fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(9)) OR (NOT
      (fsm_output(3))) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  mux_1036_nl <= MUX_s_1_2_2(mux_1035_nl, nor_1198_nl, fsm_output(2));
  and_660_nl <= (fsm_output(5)) AND mux_1036_nl;
  mux_1040_nl <= MUX_s_1_2_2(nor_1195_nl, and_660_nl, fsm_output(6));
  mux_1043_nl <= MUX_s_1_2_2(nor_1194_nl, mux_1040_nl, fsm_output(7));
  or_516_nl <= (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(3)) OR nand_398_cse;
  mux_1032_nl <= MUX_s_1_2_2(or_tmp_453, or_516_nl, fsm_output(0));
  or_514_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(9))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(4))) OR (fsm_output(10));
  mux_1033_nl <= MUX_s_1_2_2(mux_1032_nl, or_514_nl, fsm_output(2));
  nor_1199_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1033_nl);
  or_512_nl <= (NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(3)) OR nand_398_cse;
  mux_1030_nl <= MUX_s_1_2_2(or_512_nl, or_tmp_453, fsm_output(0));
  and_661_nl <= (fsm_output(5)) AND (fsm_output(2)) AND (NOT mux_1030_nl);
  nor_1200_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(2))) OR (fsm_output(0))
      OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(4))
      OR (fsm_output(10)));
  mux_1031_nl <= MUX_s_1_2_2(and_661_nl, nor_1200_nl, fsm_output(6));
  mux_1034_nl <= MUX_s_1_2_2(nor_1199_nl, mux_1031_nl, fsm_output(7));
  mux_1044_nl <= MUX_s_1_2_2(mux_1043_nl, mux_1034_nl, fsm_output(8));
  and_145_nl <= not_tmp_240 AND and_dcpl_101 AND (fsm_output(1)) AND (fsm_output(7))
      AND (fsm_output(2)) AND nor_610_cse;
  nor_1191_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(2))) OR (fsm_output(5))
      OR (fsm_output(7)) OR (fsm_output(0)) OR (fsm_output(1)));
  nor_1192_nl <= NOT((fsm_output(8)) OR (fsm_output(2)) OR (NOT((fsm_output(5)) AND
      (fsm_output(7)) AND (fsm_output(0)) AND (fsm_output(1)))));
  mux_1046_nl <= MUX_s_1_2_2(nor_1191_nl, nor_1192_nl, fsm_output(4));
  and_153_nl <= mux_1046_nl AND and_dcpl_123 AND (fsm_output(6)) AND (NOT (fsm_output(9)));
  nor_1189_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(0)));
  nor_1190_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT (fsm_output(0))));
  mux_1047_nl <= MUX_s_1_2_2(nor_1189_nl, nor_1190_nl, fsm_output(4));
  and_162_nl <= mux_1047_nl AND and_dcpl_101 AND (NOT (fsm_output(1))) AND (fsm_output(5))
      AND (NOT (fsm_output(2))) AND and_dcpl_148;
  nor_1187_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (fsm_output(1)));
  nor_1188_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(7))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(1))));
  mux_1048_nl <= MUX_s_1_2_2(nor_1187_nl, nor_1188_nl, fsm_output(9));
  and_170_nl <= mux_1048_nl AND and_dcpl_101 AND and_dcpl_21;
  and_179_nl <= mux_tmp_1049 AND and_dcpl_124 AND (NOT (fsm_output(7))) AND (fsm_output(5))
      AND (NOT (fsm_output(2))) AND and_dcpl_165;
  nor_1185_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(0))
      OR (fsm_output(1)) OR (fsm_output(3)));
  nor_1186_nl <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (NOT((fsm_output(0)) AND
      (fsm_output(1)) AND (fsm_output(3)))));
  mux_1050_nl <= MUX_s_1_2_2(nor_1185_nl, nor_1186_nl, fsm_output(2));
  and_188_nl <= mux_1050_nl AND (NOT (fsm_output(10))) AND (fsm_output(7)) AND (NOT
      (fsm_output(8))) AND and_dcpl_50;
  nor_1183_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(0))));
  nor_1184_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7)))
      OR (fsm_output(0)));
  mux_1051_nl <= MUX_s_1_2_2(nor_1183_nl, nor_1184_nl, fsm_output(4));
  and_197_nl <= mux_1051_nl AND (NOT (fsm_output(10))) AND (NOT (fsm_output(3)))
      AND (NOT (fsm_output(1))) AND (fsm_output(6)) AND (fsm_output(2)) AND (fsm_output(9));
  nor_1181_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(6))
      OR (fsm_output(0)) OR (NOT (fsm_output(1))));
  nor_1182_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(0))) OR (fsm_output(1)));
  mux_1052_nl <= MUX_s_1_2_2(nor_1181_nl, nor_1182_nl, fsm_output(4));
  and_205_nl <= mux_1052_nl AND and_dcpl_123 AND (NOT (fsm_output(2))) AND (fsm_output(8))
      AND (fsm_output(9));
  nor_1179_nl <= NOT((fsm_output(4)) OR (fsm_output(8)) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT((fsm_output(0)) AND (fsm_output(10)))));
  nor_1180_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(7))) OR (fsm_output(0)) OR (fsm_output(10)));
  mux_1053_nl <= MUX_s_1_2_2(nor_1179_nl, nor_1180_nl, fsm_output(9));
  and_211_nl <= mux_1053_nl AND (fsm_output(3)) AND (fsm_output(1)) AND (NOT (fsm_output(6)))
      AND (fsm_output(2));
  nor_1177_nl <= NOT((fsm_output(2)) OR (fsm_output(6)) OR nand_237_cse);
  nor_1178_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(6))) OR (fsm_output(0))
      OR (fsm_output(1)));
  mux_1054_nl <= MUX_s_1_2_2(nor_1177_nl, nor_1178_nl, fsm_output(4));
  and_220_nl <= mux_1054_nl AND (fsm_output(10)) AND (NOT (fsm_output(3))) AND (NOT
      (fsm_output(7))) AND (fsm_output(5)) AND nor_610_cse;
  and_231_nl <= mux_tmp_1049 AND and_dcpl_215 AND (fsm_output(7)) AND (NOT (fsm_output(5)))
      AND (NOT (fsm_output(2))) AND nor_610_cse;
  nor_1175_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(0))) OR (fsm_output(1)));
  nor_1176_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(7)) OR (fsm_output(6))
      OR (fsm_output(0)) OR (NOT (fsm_output(1))));
  mux_1055_nl <= MUX_s_1_2_2(nor_1175_nl, nor_1176_nl, fsm_output(4));
  and_238_nl <= mux_1055_nl AND nor_tmp_6 AND (fsm_output(5)) AND (fsm_output(2))
      AND (NOT (fsm_output(9)));
  and_817_nl <= (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(6))) AND
      (fsm_output(0));
  nor_1174_nl <= NOT((fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(6)))
      OR (fsm_output(0)));
  mux_1056_nl <= MUX_s_1_2_2(and_817_nl, nor_1174_nl, fsm_output(4));
  and_246_nl <= mux_1056_nl AND (fsm_output(10)) AND (NOT (fsm_output(3))) AND (fsm_output(1))
      AND (NOT (fsm_output(2))) AND and_dcpl_148;
  and_657_nl <= (fsm_output(4)) AND (fsm_output(8)) AND (fsm_output(2)) AND (fsm_output(5))
      AND (fsm_output(7)) AND (fsm_output(0)) AND (fsm_output(1)) AND (NOT (fsm_output(3)));
  nor_1172_nl <= NOT((fsm_output(4)) OR (fsm_output(8)) OR (fsm_output(2)) OR (fsm_output(5))
      OR (fsm_output(7)) OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT (fsm_output(3))));
  mux_1057_nl <= MUX_s_1_2_2(and_657_nl, nor_1172_nl, fsm_output(9));
  and_253_nl <= mux_1057_nl AND and_dcpl_243;
  and_261_nl <= not_tmp_240 AND nor_tmp_6 AND (NOT (fsm_output(1))) AND (NOT (fsm_output(7)))
      AND (fsm_output(2)) AND and_dcpl_165;
  vec_rsc_0_0_i_adra_d_pff <= MUX1HOT_v_8_19_2(COMP_LOOP_acc_psp_sva_1, (z_out_7(12
      DOWNTO 5)), COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_12_1_1_sva(11 DOWNTO
      4)), (COMP_LOOP_acc_1_cse_2_sva(11 DOWNTO 4)), (COMP_LOOP_acc_11_psp_sva(10
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_4_sva(11 DOWNTO 4)), (COMP_LOOP_acc_13_psp_sva(9
      DOWNTO 2)), (COMP_LOOP_acc_1_cse_6_sva(11 DOWNTO 4)), (COMP_LOOP_acc_14_psp_sva(10
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_8_sva(11 DOWNTO 4)), (COMP_LOOP_acc_16_psp_sva(8
      DOWNTO 1)), (COMP_LOOP_acc_1_cse_10_sva(11 DOWNTO 4)), (COMP_LOOP_acc_17_psp_sva(10
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_12_sva(11 DOWNTO 4)), (COMP_LOOP_acc_19_psp_sva(9
      DOWNTO 2)), (COMP_LOOP_acc_1_cse_14_sva(11 DOWNTO 4)), (COMP_LOOP_acc_20_psp_sva(10
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_sva(11 DOWNTO 4)), STD_LOGIC_VECTOR'( and_dcpl_119
      & COMP_LOOP_or_32_cse & and_139_nl & mux_1044_nl & and_145_nl & and_153_nl
      & and_162_nl & and_170_nl & and_179_nl & and_188_nl & and_197_nl & and_205_nl
      & and_211_nl & and_220_nl & and_231_nl & and_238_nl & and_246_nl & and_253_nl
      & and_261_nl));
  vec_rsc_0_0_i_da_d_pff <= modulo_result_mux_1_cse;
  or_624_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR
      (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1093_nl <= MUX_s_1_2_2(or_624_nl, or_622_cse, fsm_output(5));
  mux_1094_nl <= MUX_s_1_2_2(mux_1093_nl, or_621_cse, fsm_output(4));
  or_615_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1090_nl <= MUX_s_1_2_2(or_617_cse, or_615_nl, fsm_output(5));
  mux_1091_nl <= MUX_s_1_2_2(mux_1090_nl, mux_tmp_1068, fsm_output(4));
  mux_1095_nl <= MUX_s_1_2_2(mux_1094_nl, mux_1091_nl, fsm_output(7));
  mux_1089_nl <= MUX_s_1_2_2(mux_tmp_1067, mux_1088_cse, fsm_output(7));
  mux_1096_nl <= MUX_s_1_2_2(mux_1095_nl, mux_1089_nl, fsm_output(2));
  or_605_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1082_nl <= MUX_s_1_2_2(or_607_cse, or_605_nl, fsm_output(5));
  mux_1083_nl <= MUX_s_1_2_2(or_609_cse, mux_1082_nl, fsm_output(4));
  mux_1081_nl <= MUX_s_1_2_2(mux_tmp_1062, nand_25_cse, fsm_output(4));
  mux_1084_nl <= MUX_s_1_2_2(mux_1083_nl, mux_1081_nl, fsm_output(7));
  or_602_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1076_nl <= MUX_s_1_2_2(or_602_nl, or_601_cse, fsm_output(0));
  mux_1077_nl <= MUX_s_1_2_2(mux_1076_nl, or_tmp_515, fsm_output(5));
  mux_1078_nl <= MUX_s_1_2_2(or_tmp_518, mux_1077_nl, fsm_output(4));
  or_597_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1074_nl <= MUX_s_1_2_2(mux_1073_cse, or_597_nl, fsm_output(5));
  mux_1075_nl <= MUX_s_1_2_2(mux_1074_nl, or_596_cse, fsm_output(4));
  mux_1079_nl <= MUX_s_1_2_2(mux_1078_nl, mux_1075_nl, fsm_output(7));
  mux_1085_nl <= MUX_s_1_2_2(mux_1084_nl, mux_1079_nl, fsm_output(2));
  mux_1097_nl <= MUX_s_1_2_2(mux_1096_nl, mux_1085_nl, fsm_output(1));
  or_594_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_592_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1069_nl <= MUX_s_1_2_2(or_592_nl, mux_tmp_1068, fsm_output(4));
  mux_1070_nl <= MUX_s_1_2_2(or_594_nl, mux_1069_nl, fsm_output(7));
  or_588_nl <= (fsm_output(7)) OR mux_tmp_1067;
  mux_1071_nl <= MUX_s_1_2_2(mux_1070_nl, or_588_nl, fsm_output(2));
  or_581_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_580_nl <= (fsm_output(4)) OR mux_tmp_1062;
  mux_1063_nl <= MUX_s_1_2_2(or_581_nl, or_580_nl, fsm_output(7));
  or_573_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1058_nl <= MUX_s_1_2_2(or_573_nl, or_tmp_515, fsm_output(5));
  mux_1059_nl <= MUX_s_1_2_2(or_tmp_518, mux_1058_nl, fsm_output(4));
  or_570_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1060_nl <= MUX_s_1_2_2(mux_1059_nl, or_570_nl, fsm_output(7));
  mux_1064_nl <= MUX_s_1_2_2(mux_1063_nl, mux_1060_nl, fsm_output(2));
  mux_1072_nl <= MUX_s_1_2_2(mux_1071_nl, mux_1064_nl, fsm_output(1));
  or_569_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  mux_1098_nl <= MUX_s_1_2_2(mux_1097_nl, mux_1072_nl, or_569_nl);
  vec_rsc_0_0_i_wea_d_pff <= NOT mux_1098_nl;
  nor_1148_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_642_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_1147_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1149_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1125_nl <= MUX_s_1_2_2(nor_1148_cse, nor_1149_nl, fsm_output(0));
  mux_1126_nl <= MUX_s_1_2_2(nor_1147_nl, mux_1125_nl, fsm_output(8));
  and_654_nl <= nor_223_cse AND mux_1126_nl;
  or_670_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_669_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1123_nl <= MUX_s_1_2_2(or_670_nl, or_669_nl, fsm_output(0));
  nor_1150_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1123_nl);
  nor_1151_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_1152_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1122_nl <= MUX_s_1_2_2(nor_1151_nl, nor_1152_nl, fsm_output(7));
  mux_1124_nl <= MUX_s_1_2_2(nor_1150_nl, mux_1122_nl, fsm_output(6));
  mux_1127_nl <= MUX_s_1_2_2(and_654_nl, mux_1124_nl, fsm_output(5));
  nor_1153_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_661_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_659_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1118_nl <= MUX_s_1_2_2(or_661_nl, or_659_nl, fsm_output(0));
  nor_1154_nl <= NOT((fsm_output(8)) OR mux_1118_nl);
  nor_1155_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1119_nl <= MUX_s_1_2_2(nor_1154_nl, nor_1155_nl, fsm_output(7));
  mux_1120_nl <= MUX_s_1_2_2(nor_1153_nl, mux_1119_nl, fsm_output(6));
  nor_1156_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_1157_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR
      (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1158_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1115_nl <= MUX_s_1_2_2(nor_1158_nl, nor_1148_cse, fsm_output(0));
  mux_1116_nl <= MUX_s_1_2_2(nor_1157_nl, mux_1115_nl, fsm_output(8));
  and_655_nl <= (fsm_output(7)) AND mux_1116_nl;
  mux_1117_nl <= MUX_s_1_2_2(nor_1156_nl, and_655_nl, fsm_output(6));
  mux_1121_nl <= MUX_s_1_2_2(mux_1120_nl, mux_1117_nl, fsm_output(5));
  mux_1128_nl <= MUX_s_1_2_2(mux_1127_nl, mux_1121_nl, fsm_output(2));
  or_650_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_649_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1111_nl <= MUX_s_1_2_2(or_650_nl, or_649_nl, fsm_output(0));
  or_648_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_646_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (VEC_LOOP_j_sva_11_0(2)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  mux_1110_nl <= MUX_s_1_2_2(or_648_nl, or_646_nl, fsm_output(0));
  mux_1112_nl <= MUX_s_1_2_2(mux_1111_nl, mux_1110_nl, fsm_output(8));
  nor_1160_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1112_nl);
  nor_1161_nl <= NOT((fsm_output(8)) OR (VEC_LOOP_j_sva_11_0(3)) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_641_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1107_nl <= MUX_s_1_2_2(or_642_cse, or_641_nl, fsm_output(0));
  nor_1162_nl <= NOT((fsm_output(8)) OR mux_1107_nl);
  mux_1108_nl <= MUX_s_1_2_2(nor_1161_nl, nor_1162_nl, fsm_output(7));
  nor_1163_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_1164_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1106_nl <= MUX_s_1_2_2(nor_1163_nl, nor_1164_nl, fsm_output(7));
  mux_1109_nl <= MUX_s_1_2_2(mux_1108_nl, mux_1106_nl, fsm_output(6));
  mux_1113_nl <= MUX_s_1_2_2(nor_1160_nl, mux_1109_nl, fsm_output(5));
  or_635_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_633_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1102_nl <= MUX_s_1_2_2(or_633_nl, or_642_cse, fsm_output(0));
  mux_1103_nl <= MUX_s_1_2_2(or_635_nl, mux_1102_nl, fsm_output(8));
  or_630_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1104_nl <= MUX_s_1_2_2(mux_1103_nl, or_630_nl, fsm_output(7));
  nor_1165_nl <= NOT((fsm_output(6)) OR mux_1104_nl);
  nor_1166_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1167_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1168_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1099_nl <= MUX_s_1_2_2(nor_1167_nl, nor_1168_nl, fsm_output(0));
  mux_1100_nl <= MUX_s_1_2_2(nor_1166_nl, mux_1099_nl, fsm_output(8));
  and_656_nl <= (fsm_output(7)) AND mux_1100_nl;
  nor_1169_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1101_nl <= MUX_s_1_2_2(and_656_nl, nor_1169_nl, fsm_output(6));
  mux_1105_nl <= MUX_s_1_2_2(nor_1165_nl, mux_1101_nl, fsm_output(5));
  mux_1114_nl <= MUX_s_1_2_2(mux_1113_nl, mux_1105_nl, fsm_output(2));
  vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1128_nl, mux_1114_nl,
      fsm_output(4));
  or_730_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_728_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("000")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1166_nl <= MUX_s_1_2_2(or_728_nl, mux_tmp_1152, fsm_output(4));
  mux_1167_nl <= MUX_s_1_2_2(or_730_nl, mux_1166_nl, fsm_output(7));
  or_727_nl <= (fsm_output(7)) OR mux_tmp_1150;
  mux_1168_nl <= MUX_s_1_2_2(mux_1167_nl, or_727_nl, fsm_output(2));
  or_726_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_725_nl <= (fsm_output(4)) OR mux_tmp_1139;
  mux_1164_nl <= MUX_s_1_2_2(or_726_nl, or_725_nl, fsm_output(7));
  or_724_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1161_nl <= MUX_s_1_2_2(or_724_nl, or_tmp_626, fsm_output(5));
  mux_1162_nl <= MUX_s_1_2_2(or_tmp_630, mux_1161_nl, fsm_output(4));
  or_723_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1163_nl <= MUX_s_1_2_2(mux_1162_nl, or_723_nl, fsm_output(7));
  mux_1165_nl <= MUX_s_1_2_2(mux_1164_nl, mux_1163_nl, fsm_output(2));
  mux_1169_nl <= MUX_s_1_2_2(mux_1168_nl, mux_1165_nl, fsm_output(1));
  or_722_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1156_nl <= MUX_s_1_2_2(or_722_nl, or_622_cse, fsm_output(5));
  mux_1157_nl <= MUX_s_1_2_2(mux_1156_nl, or_621_cse, fsm_output(4));
  or_713_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(3)) OR
      (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1153_nl <= MUX_s_1_2_2(or_617_cse, or_713_nl, fsm_output(5));
  mux_1154_nl <= MUX_s_1_2_2(mux_1153_nl, mux_tmp_1152, fsm_output(4));
  mux_1158_nl <= MUX_s_1_2_2(mux_1157_nl, mux_1154_nl, fsm_output(7));
  mux_1151_nl <= MUX_s_1_2_2(mux_tmp_1150, mux_1088_cse, fsm_output(7));
  mux_1159_nl <= MUX_s_1_2_2(mux_1158_nl, mux_1151_nl, fsm_output(2));
  or_694_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1141_nl <= MUX_s_1_2_2(or_607_cse, or_694_nl, fsm_output(5));
  mux_1142_nl <= MUX_s_1_2_2(or_609_cse, mux_1141_nl, fsm_output(4));
  mux_1140_nl <= MUX_s_1_2_2(mux_tmp_1139, nand_25_cse, fsm_output(4));
  mux_1143_nl <= MUX_s_1_2_2(mux_1142_nl, mux_1140_nl, fsm_output(7));
  or_685_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1133_nl <= MUX_s_1_2_2(or_685_nl, or_601_cse, fsm_output(0));
  mux_1134_nl <= MUX_s_1_2_2(mux_1133_nl, or_tmp_626, fsm_output(5));
  mux_1135_nl <= MUX_s_1_2_2(or_tmp_630, mux_1134_nl, fsm_output(4));
  or_678_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1131_nl <= MUX_s_1_2_2(mux_1073_cse, or_678_nl, fsm_output(5));
  mux_1132_nl <= MUX_s_1_2_2(mux_1131_nl, or_596_cse, fsm_output(4));
  mux_1136_nl <= MUX_s_1_2_2(mux_1135_nl, mux_1132_nl, fsm_output(7));
  mux_1144_nl <= MUX_s_1_2_2(mux_1143_nl, mux_1136_nl, fsm_output(2));
  mux_1160_nl <= MUX_s_1_2_2(mux_1159_nl, mux_1144_nl, fsm_output(1));
  nor_224_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")));
  mux_1170_nl <= MUX_s_1_2_2(mux_1169_nl, mux_1160_nl, nor_224_nl);
  vec_rsc_0_1_i_wea_d_pff <= NOT mux_1170_nl;
  nor_1123_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_748_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_1122_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1124_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1197_nl <= MUX_s_1_2_2(nor_1123_cse, nor_1124_nl, fsm_output(0));
  mux_1198_nl <= MUX_s_1_2_2(nor_1122_nl, mux_1197_nl, fsm_output(8));
  and_651_nl <= nor_223_cse AND mux_1198_nl;
  or_776_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_775_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1195_nl <= MUX_s_1_2_2(or_776_nl, or_775_nl, fsm_output(0));
  nor_1125_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1195_nl);
  nor_1126_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_1127_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1194_nl <= MUX_s_1_2_2(nor_1126_nl, nor_1127_nl, fsm_output(7));
  mux_1196_nl <= MUX_s_1_2_2(nor_1125_nl, mux_1194_nl, fsm_output(6));
  mux_1199_nl <= MUX_s_1_2_2(and_651_nl, mux_1196_nl, fsm_output(5));
  nor_1128_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_767_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_765_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1190_nl <= MUX_s_1_2_2(or_767_nl, or_765_nl, fsm_output(0));
  nor_1129_nl <= NOT((fsm_output(8)) OR mux_1190_nl);
  nor_1130_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1191_nl <= MUX_s_1_2_2(nor_1129_nl, nor_1130_nl, fsm_output(7));
  mux_1192_nl <= MUX_s_1_2_2(nor_1128_nl, mux_1191_nl, fsm_output(6));
  nor_1131_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_1132_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR
      (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1133_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1187_nl <= MUX_s_1_2_2(nor_1133_nl, nor_1123_cse, fsm_output(0));
  mux_1188_nl <= MUX_s_1_2_2(nor_1132_nl, mux_1187_nl, fsm_output(8));
  and_652_nl <= (fsm_output(7)) AND mux_1188_nl;
  mux_1189_nl <= MUX_s_1_2_2(nor_1131_nl, and_652_nl, fsm_output(6));
  mux_1193_nl <= MUX_s_1_2_2(mux_1192_nl, mux_1189_nl, fsm_output(5));
  mux_1200_nl <= MUX_s_1_2_2(mux_1199_nl, mux_1193_nl, fsm_output(2));
  or_756_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_755_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1183_nl <= MUX_s_1_2_2(or_756_nl, or_755_nl, fsm_output(0));
  or_754_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_752_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (VEC_LOOP_j_sva_11_0(2)) OR (NOT
      (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1182_nl <= MUX_s_1_2_2(or_754_nl, or_752_nl, fsm_output(0));
  mux_1184_nl <= MUX_s_1_2_2(mux_1183_nl, mux_1182_nl, fsm_output(8));
  nor_1135_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1184_nl);
  nor_1136_nl <= NOT((fsm_output(8)) OR (VEC_LOOP_j_sva_11_0(3)) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_747_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1179_nl <= MUX_s_1_2_2(or_748_cse, or_747_nl, fsm_output(0));
  nor_1137_nl <= NOT((fsm_output(8)) OR mux_1179_nl);
  mux_1180_nl <= MUX_s_1_2_2(nor_1136_nl, nor_1137_nl, fsm_output(7));
  nor_1138_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_1139_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1178_nl <= MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, fsm_output(7));
  mux_1181_nl <= MUX_s_1_2_2(mux_1180_nl, mux_1178_nl, fsm_output(6));
  mux_1185_nl <= MUX_s_1_2_2(nor_1135_nl, mux_1181_nl, fsm_output(5));
  or_741_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_739_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1174_nl <= MUX_s_1_2_2(or_739_nl, or_748_cse, fsm_output(0));
  mux_1175_nl <= MUX_s_1_2_2(or_741_nl, mux_1174_nl, fsm_output(8));
  or_736_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1176_nl <= MUX_s_1_2_2(mux_1175_nl, or_736_nl, fsm_output(7));
  nor_1140_nl <= NOT((fsm_output(6)) OR mux_1176_nl);
  nor_1141_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1142_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1143_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1171_nl <= MUX_s_1_2_2(nor_1142_nl, nor_1143_nl, fsm_output(0));
  mux_1172_nl <= MUX_s_1_2_2(nor_1141_nl, mux_1171_nl, fsm_output(8));
  and_653_nl <= (fsm_output(7)) AND mux_1172_nl;
  nor_1144_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1173_nl <= MUX_s_1_2_2(and_653_nl, nor_1144_nl, fsm_output(6));
  mux_1177_nl <= MUX_s_1_2_2(nor_1140_nl, mux_1173_nl, fsm_output(5));
  mux_1186_nl <= MUX_s_1_2_2(mux_1185_nl, mux_1177_nl, fsm_output(2));
  vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1200_nl, mux_1186_nl,
      fsm_output(4));
  or_837_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR
      (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1237_nl <= MUX_s_1_2_2(or_837_nl, or_622_cse, fsm_output(5));
  mux_1238_nl <= MUX_s_1_2_2(mux_1237_nl, or_621_cse, fsm_output(4));
  or_828_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1234_nl <= MUX_s_1_2_2(or_617_cse, or_828_nl, fsm_output(5));
  mux_1235_nl <= MUX_s_1_2_2(mux_1234_nl, mux_tmp_1212, fsm_output(4));
  mux_1239_nl <= MUX_s_1_2_2(mux_1238_nl, mux_1235_nl, fsm_output(7));
  mux_1233_nl <= MUX_s_1_2_2(mux_tmp_1211, mux_1088_cse, fsm_output(7));
  mux_1240_nl <= MUX_s_1_2_2(mux_1239_nl, mux_1233_nl, fsm_output(2));
  or_818_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1226_nl <= MUX_s_1_2_2(or_607_cse, or_818_nl, fsm_output(5));
  mux_1227_nl <= MUX_s_1_2_2(or_609_cse, mux_1226_nl, fsm_output(4));
  mux_1225_nl <= MUX_s_1_2_2(mux_tmp_1206, nand_25_cse, fsm_output(4));
  mux_1228_nl <= MUX_s_1_2_2(mux_1227_nl, mux_1225_nl, fsm_output(7));
  or_815_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1220_nl <= MUX_s_1_2_2(or_815_nl, or_601_cse, fsm_output(0));
  mux_1221_nl <= MUX_s_1_2_2(mux_1220_nl, or_tmp_728, fsm_output(5));
  mux_1222_nl <= MUX_s_1_2_2(or_tmp_731, mux_1221_nl, fsm_output(4));
  or_810_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1218_nl <= MUX_s_1_2_2(mux_1073_cse, or_810_nl, fsm_output(5));
  mux_1219_nl <= MUX_s_1_2_2(mux_1218_nl, or_596_cse, fsm_output(4));
  mux_1223_nl <= MUX_s_1_2_2(mux_1222_nl, mux_1219_nl, fsm_output(7));
  mux_1229_nl <= MUX_s_1_2_2(mux_1228_nl, mux_1223_nl, fsm_output(2));
  mux_1241_nl <= MUX_s_1_2_2(mux_1240_nl, mux_1229_nl, fsm_output(1));
  or_807_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_805_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1213_nl <= MUX_s_1_2_2(or_805_nl, mux_tmp_1212, fsm_output(4));
  mux_1214_nl <= MUX_s_1_2_2(or_807_nl, mux_1213_nl, fsm_output(7));
  or_801_nl <= (fsm_output(7)) OR mux_tmp_1211;
  mux_1215_nl <= MUX_s_1_2_2(mux_1214_nl, or_801_nl, fsm_output(2));
  or_794_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_793_nl <= (fsm_output(4)) OR mux_tmp_1206;
  mux_1207_nl <= MUX_s_1_2_2(or_794_nl, or_793_nl, fsm_output(7));
  or_786_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1202_nl <= MUX_s_1_2_2(or_786_nl, or_tmp_728, fsm_output(5));
  mux_1203_nl <= MUX_s_1_2_2(or_tmp_731, mux_1202_nl, fsm_output(4));
  or_783_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1204_nl <= MUX_s_1_2_2(mux_1203_nl, or_783_nl, fsm_output(7));
  mux_1208_nl <= MUX_s_1_2_2(mux_1207_nl, mux_1204_nl, fsm_output(2));
  mux_1216_nl <= MUX_s_1_2_2(mux_1215_nl, mux_1208_nl, fsm_output(1));
  or_782_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  mux_1242_nl <= MUX_s_1_2_2(mux_1241_nl, mux_1216_nl, or_782_nl);
  vec_rsc_0_2_i_wea_d_pff <= NOT mux_1242_nl;
  nor_1098_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_855_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_1097_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1099_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1269_nl <= MUX_s_1_2_2(nor_1098_cse, nor_1099_nl, fsm_output(0));
  mux_1270_nl <= MUX_s_1_2_2(nor_1097_nl, mux_1269_nl, fsm_output(8));
  and_648_nl <= nor_223_cse AND mux_1270_nl;
  or_883_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_882_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1267_nl <= MUX_s_1_2_2(or_883_nl, or_882_nl, fsm_output(0));
  nor_1100_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1267_nl);
  nor_1101_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_1102_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1266_nl <= MUX_s_1_2_2(nor_1101_nl, nor_1102_nl, fsm_output(7));
  mux_1268_nl <= MUX_s_1_2_2(nor_1100_nl, mux_1266_nl, fsm_output(6));
  mux_1271_nl <= MUX_s_1_2_2(and_648_nl, mux_1268_nl, fsm_output(5));
  nor_1103_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_874_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_872_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1262_nl <= MUX_s_1_2_2(or_874_nl, or_872_nl, fsm_output(0));
  nor_1104_nl <= NOT((fsm_output(8)) OR mux_1262_nl);
  nor_1105_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1263_nl <= MUX_s_1_2_2(nor_1104_nl, nor_1105_nl, fsm_output(7));
  mux_1264_nl <= MUX_s_1_2_2(nor_1103_nl, mux_1263_nl, fsm_output(6));
  nor_1106_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_1107_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1108_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1259_nl <= MUX_s_1_2_2(nor_1108_nl, nor_1098_cse, fsm_output(0));
  mux_1260_nl <= MUX_s_1_2_2(nor_1107_nl, mux_1259_nl, fsm_output(8));
  and_649_nl <= (fsm_output(7)) AND mux_1260_nl;
  mux_1261_nl <= MUX_s_1_2_2(nor_1106_nl, and_649_nl, fsm_output(6));
  mux_1265_nl <= MUX_s_1_2_2(mux_1264_nl, mux_1261_nl, fsm_output(5));
  mux_1272_nl <= MUX_s_1_2_2(mux_1271_nl, mux_1265_nl, fsm_output(2));
  or_863_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_862_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1255_nl <= MUX_s_1_2_2(or_863_nl, or_862_nl, fsm_output(0));
  or_861_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_859_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (VEC_LOOP_j_sva_11_0(2)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  mux_1254_nl <= MUX_s_1_2_2(or_861_nl, or_859_nl, fsm_output(0));
  mux_1256_nl <= MUX_s_1_2_2(mux_1255_nl, mux_1254_nl, fsm_output(8));
  nor_1110_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1256_nl);
  nor_1111_nl <= NOT((fsm_output(8)) OR (VEC_LOOP_j_sva_11_0(3)) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_854_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1251_nl <= MUX_s_1_2_2(or_855_cse, or_854_nl, fsm_output(0));
  nor_1112_nl <= NOT((fsm_output(8)) OR mux_1251_nl);
  mux_1252_nl <= MUX_s_1_2_2(nor_1111_nl, nor_1112_nl, fsm_output(7));
  nor_1113_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_1114_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1250_nl <= MUX_s_1_2_2(nor_1113_nl, nor_1114_nl, fsm_output(7));
  mux_1253_nl <= MUX_s_1_2_2(mux_1252_nl, mux_1250_nl, fsm_output(6));
  mux_1257_nl <= MUX_s_1_2_2(nor_1110_nl, mux_1253_nl, fsm_output(5));
  or_848_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_846_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1246_nl <= MUX_s_1_2_2(or_846_nl, or_855_cse, fsm_output(0));
  mux_1247_nl <= MUX_s_1_2_2(or_848_nl, mux_1246_nl, fsm_output(8));
  or_843_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1248_nl <= MUX_s_1_2_2(mux_1247_nl, or_843_nl, fsm_output(7));
  nor_1115_nl <= NOT((fsm_output(6)) OR mux_1248_nl);
  nor_1116_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1117_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1118_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1243_nl <= MUX_s_1_2_2(nor_1117_nl, nor_1118_nl, fsm_output(0));
  mux_1244_nl <= MUX_s_1_2_2(nor_1116_nl, mux_1243_nl, fsm_output(8));
  and_650_nl <= (fsm_output(7)) AND mux_1244_nl;
  nor_1119_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1245_nl <= MUX_s_1_2_2(and_650_nl, nor_1119_nl, fsm_output(6));
  mux_1249_nl <= MUX_s_1_2_2(nor_1115_nl, mux_1245_nl, fsm_output(5));
  mux_1258_nl <= MUX_s_1_2_2(mux_1257_nl, mux_1249_nl, fsm_output(2));
  vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1272_nl, mux_1258_nl,
      fsm_output(4));
  or_943_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_941_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1310_nl <= MUX_s_1_2_2(or_941_nl, mux_tmp_1296, fsm_output(4));
  mux_1311_nl <= MUX_s_1_2_2(or_943_nl, mux_1310_nl, fsm_output(7));
  or_940_nl <= (fsm_output(7)) OR mux_tmp_1294;
  mux_1312_nl <= MUX_s_1_2_2(mux_1311_nl, or_940_nl, fsm_output(2));
  or_939_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_938_nl <= (fsm_output(4)) OR mux_tmp_1283;
  mux_1308_nl <= MUX_s_1_2_2(or_939_nl, or_938_nl, fsm_output(7));
  or_937_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1305_nl <= MUX_s_1_2_2(or_937_nl, or_tmp_839, fsm_output(5));
  mux_1306_nl <= MUX_s_1_2_2(or_tmp_843, mux_1305_nl, fsm_output(4));
  or_936_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1307_nl <= MUX_s_1_2_2(mux_1306_nl, or_936_nl, fsm_output(7));
  mux_1309_nl <= MUX_s_1_2_2(mux_1308_nl, mux_1307_nl, fsm_output(2));
  mux_1313_nl <= MUX_s_1_2_2(mux_1312_nl, mux_1309_nl, fsm_output(1));
  or_935_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1300_nl <= MUX_s_1_2_2(or_935_nl, or_622_cse, fsm_output(5));
  mux_1301_nl <= MUX_s_1_2_2(mux_1300_nl, or_621_cse, fsm_output(4));
  or_926_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(3)) OR
      (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1297_nl <= MUX_s_1_2_2(or_617_cse, or_926_nl, fsm_output(5));
  mux_1298_nl <= MUX_s_1_2_2(mux_1297_nl, mux_tmp_1296, fsm_output(4));
  mux_1302_nl <= MUX_s_1_2_2(mux_1301_nl, mux_1298_nl, fsm_output(7));
  mux_1295_nl <= MUX_s_1_2_2(mux_tmp_1294, mux_1088_cse, fsm_output(7));
  mux_1303_nl <= MUX_s_1_2_2(mux_1302_nl, mux_1295_nl, fsm_output(2));
  or_907_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1285_nl <= MUX_s_1_2_2(or_607_cse, or_907_nl, fsm_output(5));
  mux_1286_nl <= MUX_s_1_2_2(or_609_cse, mux_1285_nl, fsm_output(4));
  mux_1284_nl <= MUX_s_1_2_2(mux_tmp_1283, nand_25_cse, fsm_output(4));
  mux_1287_nl <= MUX_s_1_2_2(mux_1286_nl, mux_1284_nl, fsm_output(7));
  or_898_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1277_nl <= MUX_s_1_2_2(or_898_nl, or_601_cse, fsm_output(0));
  mux_1278_nl <= MUX_s_1_2_2(mux_1277_nl, or_tmp_839, fsm_output(5));
  mux_1279_nl <= MUX_s_1_2_2(or_tmp_843, mux_1278_nl, fsm_output(4));
  or_891_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1275_nl <= MUX_s_1_2_2(mux_1073_cse, or_891_nl, fsm_output(5));
  mux_1276_nl <= MUX_s_1_2_2(mux_1275_nl, or_596_cse, fsm_output(4));
  mux_1280_nl <= MUX_s_1_2_2(mux_1279_nl, mux_1276_nl, fsm_output(7));
  mux_1288_nl <= MUX_s_1_2_2(mux_1287_nl, mux_1280_nl, fsm_output(2));
  mux_1304_nl <= MUX_s_1_2_2(mux_1303_nl, mux_1288_nl, fsm_output(1));
  nor_231_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")));
  mux_1314_nl <= MUX_s_1_2_2(mux_1313_nl, mux_1304_nl, nor_231_nl);
  vec_rsc_0_3_i_wea_d_pff <= NOT mux_1314_nl;
  nor_1073_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_961_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_1072_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1074_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1341_nl <= MUX_s_1_2_2(nor_1073_cse, nor_1074_nl, fsm_output(0));
  mux_1342_nl <= MUX_s_1_2_2(nor_1072_nl, mux_1341_nl, fsm_output(8));
  and_645_nl <= nor_223_cse AND mux_1342_nl;
  or_989_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_988_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1339_nl <= MUX_s_1_2_2(or_989_nl, or_988_nl, fsm_output(0));
  nor_1075_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1339_nl);
  nor_1076_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_1077_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1338_nl <= MUX_s_1_2_2(nor_1076_nl, nor_1077_nl, fsm_output(7));
  mux_1340_nl <= MUX_s_1_2_2(nor_1075_nl, mux_1338_nl, fsm_output(6));
  mux_1343_nl <= MUX_s_1_2_2(and_645_nl, mux_1340_nl, fsm_output(5));
  nor_1078_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_980_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_978_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1334_nl <= MUX_s_1_2_2(or_980_nl, or_978_nl, fsm_output(0));
  nor_1079_nl <= NOT((fsm_output(8)) OR mux_1334_nl);
  nor_1080_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1335_nl <= MUX_s_1_2_2(nor_1079_nl, nor_1080_nl, fsm_output(7));
  mux_1336_nl <= MUX_s_1_2_2(nor_1078_nl, mux_1335_nl, fsm_output(6));
  nor_1081_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_1082_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1083_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1331_nl <= MUX_s_1_2_2(nor_1083_nl, nor_1073_cse, fsm_output(0));
  mux_1332_nl <= MUX_s_1_2_2(nor_1082_nl, mux_1331_nl, fsm_output(8));
  and_646_nl <= (fsm_output(7)) AND mux_1332_nl;
  mux_1333_nl <= MUX_s_1_2_2(nor_1081_nl, and_646_nl, fsm_output(6));
  mux_1337_nl <= MUX_s_1_2_2(mux_1336_nl, mux_1333_nl, fsm_output(5));
  mux_1344_nl <= MUX_s_1_2_2(mux_1343_nl, mux_1337_nl, fsm_output(2));
  or_969_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_968_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1327_nl <= MUX_s_1_2_2(or_969_nl, or_968_nl, fsm_output(0));
  or_967_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_965_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (VEC_LOOP_j_sva_11_0(2)) OR (NOT
      (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1326_nl <= MUX_s_1_2_2(or_967_nl, or_965_nl, fsm_output(0));
  mux_1328_nl <= MUX_s_1_2_2(mux_1327_nl, mux_1326_nl, fsm_output(8));
  nor_1085_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1328_nl);
  nor_1086_nl <= NOT((fsm_output(8)) OR (VEC_LOOP_j_sva_11_0(3)) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_960_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1323_nl <= MUX_s_1_2_2(or_961_cse, or_960_nl, fsm_output(0));
  nor_1087_nl <= NOT((fsm_output(8)) OR mux_1323_nl);
  mux_1324_nl <= MUX_s_1_2_2(nor_1086_nl, nor_1087_nl, fsm_output(7));
  nor_1088_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_1089_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1322_nl <= MUX_s_1_2_2(nor_1088_nl, nor_1089_nl, fsm_output(7));
  mux_1325_nl <= MUX_s_1_2_2(mux_1324_nl, mux_1322_nl, fsm_output(6));
  mux_1329_nl <= MUX_s_1_2_2(nor_1085_nl, mux_1325_nl, fsm_output(5));
  or_954_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_952_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1318_nl <= MUX_s_1_2_2(or_952_nl, or_961_cse, fsm_output(0));
  mux_1319_nl <= MUX_s_1_2_2(or_954_nl, mux_1318_nl, fsm_output(8));
  or_949_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1320_nl <= MUX_s_1_2_2(mux_1319_nl, or_949_nl, fsm_output(7));
  nor_1090_nl <= NOT((fsm_output(6)) OR mux_1320_nl);
  nor_1091_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1092_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1093_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1315_nl <= MUX_s_1_2_2(nor_1092_nl, nor_1093_nl, fsm_output(0));
  mux_1316_nl <= MUX_s_1_2_2(nor_1091_nl, mux_1315_nl, fsm_output(8));
  and_647_nl <= (fsm_output(7)) AND mux_1316_nl;
  nor_1094_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1317_nl <= MUX_s_1_2_2(and_647_nl, nor_1094_nl, fsm_output(6));
  mux_1321_nl <= MUX_s_1_2_2(nor_1090_nl, mux_1317_nl, fsm_output(5));
  mux_1330_nl <= MUX_s_1_2_2(mux_1329_nl, mux_1321_nl, fsm_output(2));
  vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1344_nl, mux_1330_nl,
      fsm_output(4));
  or_1050_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR
      (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1381_nl <= MUX_s_1_2_2(or_1050_nl, or_622_cse, fsm_output(5));
  mux_1382_nl <= MUX_s_1_2_2(mux_1381_nl, or_621_cse, fsm_output(4));
  or_1041_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1378_nl <= MUX_s_1_2_2(or_617_cse, or_1041_nl, fsm_output(5));
  mux_1379_nl <= MUX_s_1_2_2(mux_1378_nl, mux_tmp_1356, fsm_output(4));
  mux_1383_nl <= MUX_s_1_2_2(mux_1382_nl, mux_1379_nl, fsm_output(7));
  mux_1377_nl <= MUX_s_1_2_2(mux_tmp_1355, mux_1088_cse, fsm_output(7));
  mux_1384_nl <= MUX_s_1_2_2(mux_1383_nl, mux_1377_nl, fsm_output(2));
  or_1031_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1370_nl <= MUX_s_1_2_2(or_607_cse, or_1031_nl, fsm_output(5));
  mux_1371_nl <= MUX_s_1_2_2(or_609_cse, mux_1370_nl, fsm_output(4));
  mux_1369_nl <= MUX_s_1_2_2(mux_tmp_1350, nand_25_cse, fsm_output(4));
  mux_1372_nl <= MUX_s_1_2_2(mux_1371_nl, mux_1369_nl, fsm_output(7));
  or_1028_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1364_nl <= MUX_s_1_2_2(or_1028_nl, or_601_cse, fsm_output(0));
  mux_1365_nl <= MUX_s_1_2_2(mux_1364_nl, or_tmp_941, fsm_output(5));
  mux_1366_nl <= MUX_s_1_2_2(or_tmp_944, mux_1365_nl, fsm_output(4));
  or_1023_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1362_nl <= MUX_s_1_2_2(mux_1073_cse, or_1023_nl, fsm_output(5));
  mux_1363_nl <= MUX_s_1_2_2(mux_1362_nl, or_596_cse, fsm_output(4));
  mux_1367_nl <= MUX_s_1_2_2(mux_1366_nl, mux_1363_nl, fsm_output(7));
  mux_1373_nl <= MUX_s_1_2_2(mux_1372_nl, mux_1367_nl, fsm_output(2));
  mux_1385_nl <= MUX_s_1_2_2(mux_1384_nl, mux_1373_nl, fsm_output(1));
  or_1020_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_1018_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1357_nl <= MUX_s_1_2_2(or_1018_nl, mux_tmp_1356, fsm_output(4));
  mux_1358_nl <= MUX_s_1_2_2(or_1020_nl, mux_1357_nl, fsm_output(7));
  or_1014_nl <= (fsm_output(7)) OR mux_tmp_1355;
  mux_1359_nl <= MUX_s_1_2_2(mux_1358_nl, or_1014_nl, fsm_output(2));
  or_1007_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_1006_nl <= (fsm_output(4)) OR mux_tmp_1350;
  mux_1351_nl <= MUX_s_1_2_2(or_1007_nl, or_1006_nl, fsm_output(7));
  or_999_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1346_nl <= MUX_s_1_2_2(or_999_nl, or_tmp_941, fsm_output(5));
  mux_1347_nl <= MUX_s_1_2_2(or_tmp_944, mux_1346_nl, fsm_output(4));
  or_996_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1348_nl <= MUX_s_1_2_2(mux_1347_nl, or_996_nl, fsm_output(7));
  mux_1352_nl <= MUX_s_1_2_2(mux_1351_nl, mux_1348_nl, fsm_output(2));
  mux_1360_nl <= MUX_s_1_2_2(mux_1359_nl, mux_1352_nl, fsm_output(1));
  or_995_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"));
  mux_1386_nl <= MUX_s_1_2_2(mux_1385_nl, mux_1360_nl, or_995_nl);
  vec_rsc_0_4_i_wea_d_pff <= NOT mux_1386_nl;
  nor_1048_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1068_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_1047_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1049_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1413_nl <= MUX_s_1_2_2(nor_1048_cse, nor_1049_nl, fsm_output(0));
  mux_1414_nl <= MUX_s_1_2_2(nor_1047_nl, mux_1413_nl, fsm_output(8));
  and_642_nl <= nor_223_cse AND mux_1414_nl;
  or_1096_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1095_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1411_nl <= MUX_s_1_2_2(or_1096_nl, or_1095_nl, fsm_output(0));
  nor_1050_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1411_nl);
  nor_1051_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_1052_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1410_nl <= MUX_s_1_2_2(nor_1051_nl, nor_1052_nl, fsm_output(7));
  mux_1412_nl <= MUX_s_1_2_2(nor_1050_nl, mux_1410_nl, fsm_output(6));
  mux_1415_nl <= MUX_s_1_2_2(and_642_nl, mux_1412_nl, fsm_output(5));
  nor_1053_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_1087_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1085_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1406_nl <= MUX_s_1_2_2(or_1087_nl, or_1085_nl, fsm_output(0));
  nor_1054_nl <= NOT((fsm_output(8)) OR mux_1406_nl);
  nor_1055_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1407_nl <= MUX_s_1_2_2(nor_1054_nl, nor_1055_nl, fsm_output(7));
  mux_1408_nl <= MUX_s_1_2_2(nor_1053_nl, mux_1407_nl, fsm_output(6));
  nor_1056_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_1057_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR
      (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1058_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1403_nl <= MUX_s_1_2_2(nor_1058_nl, nor_1048_cse, fsm_output(0));
  mux_1404_nl <= MUX_s_1_2_2(nor_1057_nl, mux_1403_nl, fsm_output(8));
  and_643_nl <= (fsm_output(7)) AND mux_1404_nl;
  mux_1405_nl <= MUX_s_1_2_2(nor_1056_nl, and_643_nl, fsm_output(6));
  mux_1409_nl <= MUX_s_1_2_2(mux_1408_nl, mux_1405_nl, fsm_output(5));
  mux_1416_nl <= MUX_s_1_2_2(mux_1415_nl, mux_1409_nl, fsm_output(2));
  or_1076_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1075_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1399_nl <= MUX_s_1_2_2(or_1076_nl, or_1075_nl, fsm_output(0));
  or_1074_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1072_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (VEC_LOOP_j_sva_11_0(2))) OR
      (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  mux_1398_nl <= MUX_s_1_2_2(or_1074_nl, or_1072_nl, fsm_output(0));
  mux_1400_nl <= MUX_s_1_2_2(mux_1399_nl, mux_1398_nl, fsm_output(8));
  nor_1060_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1400_nl);
  nor_1061_nl <= NOT((fsm_output(8)) OR (VEC_LOOP_j_sva_11_0(3)) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1067_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1395_nl <= MUX_s_1_2_2(or_1068_cse, or_1067_nl, fsm_output(0));
  nor_1062_nl <= NOT((fsm_output(8)) OR mux_1395_nl);
  mux_1396_nl <= MUX_s_1_2_2(nor_1061_nl, nor_1062_nl, fsm_output(7));
  nor_1063_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_1064_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1394_nl <= MUX_s_1_2_2(nor_1063_nl, nor_1064_nl, fsm_output(7));
  mux_1397_nl <= MUX_s_1_2_2(mux_1396_nl, mux_1394_nl, fsm_output(6));
  mux_1401_nl <= MUX_s_1_2_2(nor_1060_nl, mux_1397_nl, fsm_output(5));
  or_1061_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1059_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1390_nl <= MUX_s_1_2_2(or_1059_nl, or_1068_cse, fsm_output(0));
  mux_1391_nl <= MUX_s_1_2_2(or_1061_nl, mux_1390_nl, fsm_output(8));
  or_1056_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1392_nl <= MUX_s_1_2_2(mux_1391_nl, or_1056_nl, fsm_output(7));
  nor_1065_nl <= NOT((fsm_output(6)) OR mux_1392_nl);
  nor_1066_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1067_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1068_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1387_nl <= MUX_s_1_2_2(nor_1067_nl, nor_1068_nl, fsm_output(0));
  mux_1388_nl <= MUX_s_1_2_2(nor_1066_nl, mux_1387_nl, fsm_output(8));
  and_644_nl <= (fsm_output(7)) AND mux_1388_nl;
  nor_1069_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1389_nl <= MUX_s_1_2_2(and_644_nl, nor_1069_nl, fsm_output(6));
  mux_1393_nl <= MUX_s_1_2_2(nor_1065_nl, mux_1389_nl, fsm_output(5));
  mux_1402_nl <= MUX_s_1_2_2(mux_1401_nl, mux_1393_nl, fsm_output(2));
  vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1416_nl, mux_1402_nl,
      fsm_output(4));
  or_1156_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_1154_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1454_nl <= MUX_s_1_2_2(or_1154_nl, mux_tmp_1440, fsm_output(4));
  mux_1455_nl <= MUX_s_1_2_2(or_1156_nl, mux_1454_nl, fsm_output(7));
  or_1153_nl <= (fsm_output(7)) OR mux_tmp_1438;
  mux_1456_nl <= MUX_s_1_2_2(mux_1455_nl, or_1153_nl, fsm_output(2));
  or_1152_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_1151_nl <= (fsm_output(4)) OR mux_tmp_1427;
  mux_1452_nl <= MUX_s_1_2_2(or_1152_nl, or_1151_nl, fsm_output(7));
  or_1150_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1449_nl <= MUX_s_1_2_2(or_1150_nl, or_tmp_1052, fsm_output(5));
  mux_1450_nl <= MUX_s_1_2_2(or_tmp_1056, mux_1449_nl, fsm_output(4));
  or_1149_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1451_nl <= MUX_s_1_2_2(mux_1450_nl, or_1149_nl, fsm_output(7));
  mux_1453_nl <= MUX_s_1_2_2(mux_1452_nl, mux_1451_nl, fsm_output(2));
  mux_1457_nl <= MUX_s_1_2_2(mux_1456_nl, mux_1453_nl, fsm_output(1));
  or_1148_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1444_nl <= MUX_s_1_2_2(or_1148_nl, or_622_cse, fsm_output(5));
  mux_1445_nl <= MUX_s_1_2_2(mux_1444_nl, or_621_cse, fsm_output(4));
  or_1139_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(3)) OR
      (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1441_nl <= MUX_s_1_2_2(or_617_cse, or_1139_nl, fsm_output(5));
  mux_1442_nl <= MUX_s_1_2_2(mux_1441_nl, mux_tmp_1440, fsm_output(4));
  mux_1446_nl <= MUX_s_1_2_2(mux_1445_nl, mux_1442_nl, fsm_output(7));
  mux_1439_nl <= MUX_s_1_2_2(mux_tmp_1438, mux_1088_cse, fsm_output(7));
  mux_1447_nl <= MUX_s_1_2_2(mux_1446_nl, mux_1439_nl, fsm_output(2));
  or_1120_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1429_nl <= MUX_s_1_2_2(or_607_cse, or_1120_nl, fsm_output(5));
  mux_1430_nl <= MUX_s_1_2_2(or_609_cse, mux_1429_nl, fsm_output(4));
  mux_1428_nl <= MUX_s_1_2_2(mux_tmp_1427, nand_25_cse, fsm_output(4));
  mux_1431_nl <= MUX_s_1_2_2(mux_1430_nl, mux_1428_nl, fsm_output(7));
  or_1111_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1421_nl <= MUX_s_1_2_2(or_1111_nl, or_601_cse, fsm_output(0));
  mux_1422_nl <= MUX_s_1_2_2(mux_1421_nl, or_tmp_1052, fsm_output(5));
  mux_1423_nl <= MUX_s_1_2_2(or_tmp_1056, mux_1422_nl, fsm_output(4));
  or_1104_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1419_nl <= MUX_s_1_2_2(mux_1073_cse, or_1104_nl, fsm_output(5));
  mux_1420_nl <= MUX_s_1_2_2(mux_1419_nl, or_596_cse, fsm_output(4));
  mux_1424_nl <= MUX_s_1_2_2(mux_1423_nl, mux_1420_nl, fsm_output(7));
  mux_1432_nl <= MUX_s_1_2_2(mux_1431_nl, mux_1424_nl, fsm_output(2));
  mux_1448_nl <= MUX_s_1_2_2(mux_1447_nl, mux_1432_nl, fsm_output(1));
  nor_238_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")));
  mux_1458_nl <= MUX_s_1_2_2(mux_1457_nl, mux_1448_nl, nor_238_nl);
  vec_rsc_0_5_i_wea_d_pff <= NOT mux_1458_nl;
  nor_1023_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1174_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_1022_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1024_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1485_nl <= MUX_s_1_2_2(nor_1023_cse, nor_1024_nl, fsm_output(0));
  mux_1486_nl <= MUX_s_1_2_2(nor_1022_nl, mux_1485_nl, fsm_output(8));
  and_639_nl <= nor_223_cse AND mux_1486_nl;
  or_1202_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1201_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1483_nl <= MUX_s_1_2_2(or_1202_nl, or_1201_nl, fsm_output(0));
  nor_1025_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1483_nl);
  nor_1026_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_1027_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1482_nl <= MUX_s_1_2_2(nor_1026_nl, nor_1027_nl, fsm_output(7));
  mux_1484_nl <= MUX_s_1_2_2(nor_1025_nl, mux_1482_nl, fsm_output(6));
  mux_1487_nl <= MUX_s_1_2_2(and_639_nl, mux_1484_nl, fsm_output(5));
  nor_1028_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_1193_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1191_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1478_nl <= MUX_s_1_2_2(or_1193_nl, or_1191_nl, fsm_output(0));
  nor_1029_nl <= NOT((fsm_output(8)) OR mux_1478_nl);
  nor_1030_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1479_nl <= MUX_s_1_2_2(nor_1029_nl, nor_1030_nl, fsm_output(7));
  mux_1480_nl <= MUX_s_1_2_2(nor_1028_nl, mux_1479_nl, fsm_output(6));
  nor_1031_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_1032_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR
      (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1033_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1475_nl <= MUX_s_1_2_2(nor_1033_nl, nor_1023_cse, fsm_output(0));
  mux_1476_nl <= MUX_s_1_2_2(nor_1032_nl, mux_1475_nl, fsm_output(8));
  and_640_nl <= (fsm_output(7)) AND mux_1476_nl;
  mux_1477_nl <= MUX_s_1_2_2(nor_1031_nl, and_640_nl, fsm_output(6));
  mux_1481_nl <= MUX_s_1_2_2(mux_1480_nl, mux_1477_nl, fsm_output(5));
  mux_1488_nl <= MUX_s_1_2_2(mux_1487_nl, mux_1481_nl, fsm_output(2));
  or_1182_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1181_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1471_nl <= MUX_s_1_2_2(or_1182_nl, or_1181_nl, fsm_output(0));
  or_1180_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1178_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (VEC_LOOP_j_sva_11_0(2))) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1470_nl <= MUX_s_1_2_2(or_1180_nl, or_1178_nl, fsm_output(0));
  mux_1472_nl <= MUX_s_1_2_2(mux_1471_nl, mux_1470_nl, fsm_output(8));
  nor_1035_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1472_nl);
  nor_1036_nl <= NOT((fsm_output(8)) OR (VEC_LOOP_j_sva_11_0(3)) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1173_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1467_nl <= MUX_s_1_2_2(or_1174_cse, or_1173_nl, fsm_output(0));
  nor_1037_nl <= NOT((fsm_output(8)) OR mux_1467_nl);
  mux_1468_nl <= MUX_s_1_2_2(nor_1036_nl, nor_1037_nl, fsm_output(7));
  nor_1038_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_1039_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1466_nl <= MUX_s_1_2_2(nor_1038_nl, nor_1039_nl, fsm_output(7));
  mux_1469_nl <= MUX_s_1_2_2(mux_1468_nl, mux_1466_nl, fsm_output(6));
  mux_1473_nl <= MUX_s_1_2_2(nor_1035_nl, mux_1469_nl, fsm_output(5));
  or_1167_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1165_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1462_nl <= MUX_s_1_2_2(or_1165_nl, or_1174_cse, fsm_output(0));
  mux_1463_nl <= MUX_s_1_2_2(or_1167_nl, mux_1462_nl, fsm_output(8));
  or_1162_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1464_nl <= MUX_s_1_2_2(mux_1463_nl, or_1162_nl, fsm_output(7));
  nor_1040_nl <= NOT((fsm_output(6)) OR mux_1464_nl);
  nor_1041_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1042_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1043_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1459_nl <= MUX_s_1_2_2(nor_1042_nl, nor_1043_nl, fsm_output(0));
  mux_1460_nl <= MUX_s_1_2_2(nor_1041_nl, mux_1459_nl, fsm_output(8));
  and_641_nl <= (fsm_output(7)) AND mux_1460_nl;
  nor_1044_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1461_nl <= MUX_s_1_2_2(and_641_nl, nor_1044_nl, fsm_output(6));
  mux_1465_nl <= MUX_s_1_2_2(nor_1040_nl, mux_1461_nl, fsm_output(5));
  mux_1474_nl <= MUX_s_1_2_2(mux_1473_nl, mux_1465_nl, fsm_output(2));
  vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1488_nl, mux_1474_nl,
      fsm_output(4));
  or_1263_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR
      (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1525_nl <= MUX_s_1_2_2(or_1263_nl, or_622_cse, fsm_output(5));
  mux_1526_nl <= MUX_s_1_2_2(mux_1525_nl, or_621_cse, fsm_output(4));
  or_1254_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1522_nl <= MUX_s_1_2_2(or_617_cse, or_1254_nl, fsm_output(5));
  mux_1523_nl <= MUX_s_1_2_2(mux_1522_nl, mux_tmp_1500, fsm_output(4));
  mux_1527_nl <= MUX_s_1_2_2(mux_1526_nl, mux_1523_nl, fsm_output(7));
  mux_1521_nl <= MUX_s_1_2_2(mux_tmp_1499, mux_1088_cse, fsm_output(7));
  mux_1528_nl <= MUX_s_1_2_2(mux_1527_nl, mux_1521_nl, fsm_output(2));
  or_1244_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1514_nl <= MUX_s_1_2_2(or_607_cse, or_1244_nl, fsm_output(5));
  mux_1515_nl <= MUX_s_1_2_2(or_609_cse, mux_1514_nl, fsm_output(4));
  mux_1513_nl <= MUX_s_1_2_2(mux_tmp_1494, nand_25_cse, fsm_output(4));
  mux_1516_nl <= MUX_s_1_2_2(mux_1515_nl, mux_1513_nl, fsm_output(7));
  or_1241_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1508_nl <= MUX_s_1_2_2(or_1241_nl, or_601_cse, fsm_output(0));
  mux_1509_nl <= MUX_s_1_2_2(mux_1508_nl, or_tmp_1154, fsm_output(5));
  mux_1510_nl <= MUX_s_1_2_2(or_tmp_1157, mux_1509_nl, fsm_output(4));
  or_1236_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1506_nl <= MUX_s_1_2_2(mux_1073_cse, or_1236_nl, fsm_output(5));
  mux_1507_nl <= MUX_s_1_2_2(mux_1506_nl, or_596_cse, fsm_output(4));
  mux_1511_nl <= MUX_s_1_2_2(mux_1510_nl, mux_1507_nl, fsm_output(7));
  mux_1517_nl <= MUX_s_1_2_2(mux_1516_nl, mux_1511_nl, fsm_output(2));
  mux_1529_nl <= MUX_s_1_2_2(mux_1528_nl, mux_1517_nl, fsm_output(1));
  or_1233_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_1231_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1501_nl <= MUX_s_1_2_2(or_1231_nl, mux_tmp_1500, fsm_output(4));
  mux_1502_nl <= MUX_s_1_2_2(or_1233_nl, mux_1501_nl, fsm_output(7));
  or_1227_nl <= (fsm_output(7)) OR mux_tmp_1499;
  mux_1503_nl <= MUX_s_1_2_2(mux_1502_nl, or_1227_nl, fsm_output(2));
  or_1220_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_1219_nl <= (fsm_output(4)) OR mux_tmp_1494;
  mux_1495_nl <= MUX_s_1_2_2(or_1220_nl, or_1219_nl, fsm_output(7));
  or_1212_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1490_nl <= MUX_s_1_2_2(or_1212_nl, or_tmp_1154, fsm_output(5));
  mux_1491_nl <= MUX_s_1_2_2(or_tmp_1157, mux_1490_nl, fsm_output(4));
  or_1209_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1492_nl <= MUX_s_1_2_2(mux_1491_nl, or_1209_nl, fsm_output(7));
  mux_1496_nl <= MUX_s_1_2_2(mux_1495_nl, mux_1492_nl, fsm_output(2));
  mux_1504_nl <= MUX_s_1_2_2(mux_1503_nl, mux_1496_nl, fsm_output(1));
  or_1208_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"));
  mux_1530_nl <= MUX_s_1_2_2(mux_1529_nl, mux_1504_nl, or_1208_nl);
  vec_rsc_0_6_i_wea_d_pff <= NOT mux_1530_nl;
  nor_998_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1281_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_997_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_999_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1557_nl <= MUX_s_1_2_2(nor_998_cse, nor_999_nl, fsm_output(0));
  mux_1558_nl <= MUX_s_1_2_2(nor_997_nl, mux_1557_nl, fsm_output(8));
  and_636_nl <= nor_223_cse AND mux_1558_nl;
  or_1309_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1308_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1555_nl <= MUX_s_1_2_2(or_1309_nl, or_1308_nl, fsm_output(0));
  nor_1000_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1555_nl);
  nor_1001_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_1002_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1554_nl <= MUX_s_1_2_2(nor_1001_nl, nor_1002_nl, fsm_output(7));
  mux_1556_nl <= MUX_s_1_2_2(nor_1000_nl, mux_1554_nl, fsm_output(6));
  mux_1559_nl <= MUX_s_1_2_2(and_636_nl, mux_1556_nl, fsm_output(5));
  nor_1003_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("011")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_1300_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1298_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1550_nl <= MUX_s_1_2_2(or_1300_nl, or_1298_nl, fsm_output(0));
  nor_1004_nl <= NOT((fsm_output(8)) OR mux_1550_nl);
  nor_1005_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1551_nl <= MUX_s_1_2_2(nor_1004_nl, nor_1005_nl, fsm_output(7));
  mux_1552_nl <= MUX_s_1_2_2(nor_1003_nl, mux_1551_nl, fsm_output(6));
  nor_1006_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_1007_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_1008_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1547_nl <= MUX_s_1_2_2(nor_1008_nl, nor_998_cse, fsm_output(0));
  mux_1548_nl <= MUX_s_1_2_2(nor_1007_nl, mux_1547_nl, fsm_output(8));
  and_637_nl <= (fsm_output(7)) AND mux_1548_nl;
  mux_1549_nl <= MUX_s_1_2_2(nor_1006_nl, and_637_nl, fsm_output(6));
  mux_1553_nl <= MUX_s_1_2_2(mux_1552_nl, mux_1549_nl, fsm_output(5));
  mux_1560_nl <= MUX_s_1_2_2(mux_1559_nl, mux_1553_nl, fsm_output(2));
  or_1289_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1288_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1543_nl <= MUX_s_1_2_2(or_1289_nl, or_1288_nl, fsm_output(0));
  or_1287_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1285_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (VEC_LOOP_j_sva_11_0(2))) OR
      (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT
      (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1542_nl <= MUX_s_1_2_2(or_1287_nl, or_1285_nl, fsm_output(0));
  mux_1544_nl <= MUX_s_1_2_2(mux_1543_nl, mux_1542_nl, fsm_output(8));
  nor_1010_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1544_nl);
  nor_1011_nl <= NOT((fsm_output(8)) OR (VEC_LOOP_j_sva_11_0(3)) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1280_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1539_nl <= MUX_s_1_2_2(or_1281_cse, or_1280_nl, fsm_output(0));
  nor_1012_nl <= NOT((fsm_output(8)) OR mux_1539_nl);
  mux_1540_nl <= MUX_s_1_2_2(nor_1011_nl, nor_1012_nl, fsm_output(7));
  nor_1013_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_1014_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1538_nl <= MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, fsm_output(7));
  mux_1541_nl <= MUX_s_1_2_2(mux_1540_nl, mux_1538_nl, fsm_output(6));
  mux_1545_nl <= MUX_s_1_2_2(nor_1010_nl, mux_1541_nl, fsm_output(5));
  or_1274_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1272_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1534_nl <= MUX_s_1_2_2(or_1272_nl, or_1281_cse, fsm_output(0));
  mux_1535_nl <= MUX_s_1_2_2(or_1274_nl, mux_1534_nl, fsm_output(8));
  or_1269_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1536_nl <= MUX_s_1_2_2(mux_1535_nl, or_1269_nl, fsm_output(7));
  nor_1015_nl <= NOT((fsm_output(6)) OR mux_1536_nl);
  nor_1016_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1017_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_1018_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1531_nl <= MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, fsm_output(0));
  mux_1532_nl <= MUX_s_1_2_2(nor_1016_nl, mux_1531_nl, fsm_output(8));
  and_638_nl <= (fsm_output(7)) AND mux_1532_nl;
  nor_1019_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1533_nl <= MUX_s_1_2_2(and_638_nl, nor_1019_nl, fsm_output(6));
  mux_1537_nl <= MUX_s_1_2_2(nor_1015_nl, mux_1533_nl, fsm_output(5));
  mux_1546_nl <= MUX_s_1_2_2(mux_1545_nl, mux_1537_nl, fsm_output(2));
  vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1560_nl, mux_1546_nl,
      fsm_output(4));
  or_1369_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_1367_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("011")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1598_nl <= MUX_s_1_2_2(or_1367_nl, mux_tmp_1584, fsm_output(4));
  mux_1599_nl <= MUX_s_1_2_2(or_1369_nl, mux_1598_nl, fsm_output(7));
  or_1366_nl <= (fsm_output(7)) OR mux_tmp_1582;
  mux_1600_nl <= MUX_s_1_2_2(mux_1599_nl, or_1366_nl, fsm_output(2));
  nand_336_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  or_1364_nl <= (fsm_output(4)) OR mux_tmp_1571;
  mux_1596_nl <= MUX_s_1_2_2(nand_336_nl, or_1364_nl, fsm_output(7));
  or_1363_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1593_nl <= MUX_s_1_2_2(or_1363_nl, or_tmp_1265, fsm_output(5));
  mux_1594_nl <= MUX_s_1_2_2(or_tmp_1269, mux_1593_nl, fsm_output(4));
  or_1362_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1595_nl <= MUX_s_1_2_2(mux_1594_nl, or_1362_nl, fsm_output(7));
  mux_1597_nl <= MUX_s_1_2_2(mux_1596_nl, mux_1595_nl, fsm_output(2));
  mux_1601_nl <= MUX_s_1_2_2(mux_1600_nl, mux_1597_nl, fsm_output(1));
  or_1361_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1588_nl <= MUX_s_1_2_2(or_1361_nl, or_622_cse, fsm_output(5));
  mux_1589_nl <= MUX_s_1_2_2(mux_1588_nl, or_621_cse, fsm_output(4));
  or_1352_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(3)) OR
      (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1585_nl <= MUX_s_1_2_2(or_617_cse, or_1352_nl, fsm_output(5));
  mux_1586_nl <= MUX_s_1_2_2(mux_1585_nl, mux_tmp_1584, fsm_output(4));
  mux_1590_nl <= MUX_s_1_2_2(mux_1589_nl, mux_1586_nl, fsm_output(7));
  mux_1583_nl <= MUX_s_1_2_2(mux_tmp_1582, mux_1088_cse, fsm_output(7));
  mux_1591_nl <= MUX_s_1_2_2(mux_1590_nl, mux_1583_nl, fsm_output(2));
  nand_338_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  mux_1573_nl <= MUX_s_1_2_2(or_607_cse, nand_338_nl, fsm_output(5));
  mux_1574_nl <= MUX_s_1_2_2(or_609_cse, mux_1573_nl, fsm_output(4));
  mux_1572_nl <= MUX_s_1_2_2(mux_tmp_1571, nand_25_cse, fsm_output(4));
  mux_1575_nl <= MUX_s_1_2_2(mux_1574_nl, mux_1572_nl, fsm_output(7));
  or_1324_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1565_nl <= MUX_s_1_2_2(or_1324_nl, or_601_cse, fsm_output(0));
  mux_1566_nl <= MUX_s_1_2_2(mux_1565_nl, or_tmp_1265, fsm_output(5));
  mux_1567_nl <= MUX_s_1_2_2(or_tmp_1269, mux_1566_nl, fsm_output(4));
  or_1317_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1563_nl <= MUX_s_1_2_2(mux_1073_cse, or_1317_nl, fsm_output(5));
  mux_1564_nl <= MUX_s_1_2_2(mux_1563_nl, or_596_cse, fsm_output(4));
  mux_1568_nl <= MUX_s_1_2_2(mux_1567_nl, mux_1564_nl, fsm_output(7));
  mux_1576_nl <= MUX_s_1_2_2(mux_1575_nl, mux_1568_nl, fsm_output(2));
  mux_1592_nl <= MUX_s_1_2_2(mux_1591_nl, mux_1576_nl, fsm_output(1));
  and_635_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
  mux_1602_nl <= MUX_s_1_2_2(mux_1601_nl, mux_1592_nl, and_635_nl);
  vec_rsc_0_7_i_wea_d_pff <= NOT mux_1602_nl;
  nor_975_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1387_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_974_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_976_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1629_nl <= MUX_s_1_2_2(nor_975_cse, nor_976_nl, fsm_output(0));
  mux_1630_nl <= MUX_s_1_2_2(nor_974_nl, mux_1629_nl, fsm_output(8));
  and_630_nl <= nor_223_cse AND mux_1630_nl;
  nand_333_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10))));
  or_1414_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1627_nl <= MUX_s_1_2_2(nand_333_nl, or_1414_nl, fsm_output(0));
  nor_977_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1627_nl);
  nor_978_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_979_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1626_nl <= MUX_s_1_2_2(nor_978_nl, nor_979_nl, fsm_output(7));
  mux_1628_nl <= MUX_s_1_2_2(nor_977_nl, mux_1626_nl, fsm_output(6));
  mux_1631_nl <= MUX_s_1_2_2(and_630_nl, mux_1628_nl, fsm_output(5));
  and_631_nl <= (fsm_output(7)) AND (NOT (fsm_output(8))) AND (fsm_output(0)) AND
      (VEC_LOOP_j_sva_11_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("011")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3))
      AND (fsm_output(9)) AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  or_1406_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1404_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1622_nl <= MUX_s_1_2_2(or_1406_nl, or_1404_nl, fsm_output(0));
  nor_980_nl <= NOT((fsm_output(8)) OR mux_1622_nl);
  nor_981_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1623_nl <= MUX_s_1_2_2(nor_980_nl, nor_981_nl, fsm_output(7));
  mux_1624_nl <= MUX_s_1_2_2(and_631_nl, mux_1623_nl, fsm_output(6));
  nor_982_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  and_828_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(0)) AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (VEC_LOOP_j_sva_11_0(1)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(1))) AND (fsm_output(10));
  nor_984_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1619_nl <= MUX_s_1_2_2(nor_984_nl, nor_975_cse, fsm_output(0));
  mux_1620_nl <= MUX_s_1_2_2(and_828_nl, mux_1619_nl, fsm_output(8));
  and_632_nl <= (fsm_output(7)) AND mux_1620_nl;
  mux_1621_nl <= MUX_s_1_2_2(nor_982_nl, and_632_nl, fsm_output(6));
  mux_1625_nl <= MUX_s_1_2_2(mux_1624_nl, mux_1621_nl, fsm_output(5));
  mux_1632_nl <= MUX_s_1_2_2(mux_1631_nl, mux_1625_nl, fsm_output(2));
  or_1395_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1394_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1615_nl <= MUX_s_1_2_2(or_1395_nl, or_1394_nl, fsm_output(0));
  or_1393_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1391_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR (NOT (VEC_LOOP_j_sva_11_0(2))) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1614_nl <= MUX_s_1_2_2(or_1393_nl, or_1391_nl, fsm_output(0));
  mux_1616_nl <= MUX_s_1_2_2(mux_1615_nl, mux_1614_nl, fsm_output(8));
  nor_986_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1616_nl);
  nor_987_nl <= NOT((fsm_output(8)) OR (VEC_LOOP_j_sva_11_0(3)) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1386_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1611_nl <= MUX_s_1_2_2(or_1387_cse, or_1386_nl, fsm_output(0));
  nor_988_nl <= NOT((fsm_output(8)) OR mux_1611_nl);
  mux_1612_nl <= MUX_s_1_2_2(nor_987_nl, nor_988_nl, fsm_output(7));
  nor_989_nl <= NOT((NOT((fsm_output(8)) AND (fsm_output(0)) AND (fsm_output(3))
      AND CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("0111")) AND (NOT (fsm_output(9)))))
      OR not_tmp_260);
  nor_990_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1610_nl <= MUX_s_1_2_2(nor_989_nl, nor_990_nl, fsm_output(7));
  mux_1613_nl <= MUX_s_1_2_2(mux_1612_nl, mux_1610_nl, fsm_output(6));
  mux_1617_nl <= MUX_s_1_2_2(nor_986_nl, mux_1613_nl, fsm_output(5));
  nand_417_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(0))) AND (fsm_output(3))
      AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (fsm_output(10)));
  or_1378_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1606_nl <= MUX_s_1_2_2(or_1378_nl, or_1387_cse, fsm_output(0));
  mux_1607_nl <= MUX_s_1_2_2(nand_417_nl, mux_1606_nl, fsm_output(8));
  or_1375_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1608_nl <= MUX_s_1_2_2(mux_1607_nl, or_1375_nl, fsm_output(7));
  nor_991_nl <= NOT((fsm_output(6)) OR mux_1608_nl);
  nor_992_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  and_634_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  nor_993_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1603_nl <= MUX_s_1_2_2(and_634_nl, nor_993_nl, fsm_output(0));
  mux_1604_nl <= MUX_s_1_2_2(nor_992_nl, mux_1603_nl, fsm_output(8));
  and_633_nl <= (fsm_output(7)) AND mux_1604_nl;
  nor_994_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1605_nl <= MUX_s_1_2_2(and_633_nl, nor_994_nl, fsm_output(6));
  mux_1609_nl <= MUX_s_1_2_2(nor_991_nl, mux_1605_nl, fsm_output(5));
  mux_1618_nl <= MUX_s_1_2_2(mux_1617_nl, mux_1609_nl, fsm_output(2));
  vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1632_nl, mux_1618_nl,
      fsm_output(4));
  or_1476_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR
      (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1669_nl <= MUX_s_1_2_2(or_1476_nl, or_622_cse, fsm_output(5));
  mux_1670_nl <= MUX_s_1_2_2(mux_1669_nl, or_621_cse, fsm_output(4));
  or_1467_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1666_nl <= MUX_s_1_2_2(or_617_cse, or_1467_nl, fsm_output(5));
  mux_1667_nl <= MUX_s_1_2_2(mux_1666_nl, mux_tmp_1644, fsm_output(4));
  mux_1671_nl <= MUX_s_1_2_2(mux_1670_nl, mux_1667_nl, fsm_output(7));
  mux_1665_nl <= MUX_s_1_2_2(mux_tmp_1643, mux_1088_cse, fsm_output(7));
  mux_1672_nl <= MUX_s_1_2_2(mux_1671_nl, mux_1665_nl, fsm_output(2));
  or_1457_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1658_nl <= MUX_s_1_2_2(or_607_cse, or_1457_nl, fsm_output(5));
  mux_1659_nl <= MUX_s_1_2_2(or_609_cse, mux_1658_nl, fsm_output(4));
  mux_1657_nl <= MUX_s_1_2_2(mux_tmp_1638, nand_25_cse, fsm_output(4));
  mux_1660_nl <= MUX_s_1_2_2(mux_1659_nl, mux_1657_nl, fsm_output(7));
  or_1454_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1652_nl <= MUX_s_1_2_2(or_1454_nl, or_601_cse, fsm_output(0));
  mux_1653_nl <= MUX_s_1_2_2(mux_1652_nl, or_tmp_1367, fsm_output(5));
  mux_1654_nl <= MUX_s_1_2_2(or_tmp_1370, mux_1653_nl, fsm_output(4));
  or_1449_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1650_nl <= MUX_s_1_2_2(mux_1073_cse, or_1449_nl, fsm_output(5));
  mux_1651_nl <= MUX_s_1_2_2(mux_1650_nl, or_596_cse, fsm_output(4));
  mux_1655_nl <= MUX_s_1_2_2(mux_1654_nl, mux_1651_nl, fsm_output(7));
  mux_1661_nl <= MUX_s_1_2_2(mux_1660_nl, mux_1655_nl, fsm_output(2));
  mux_1673_nl <= MUX_s_1_2_2(mux_1672_nl, mux_1661_nl, fsm_output(1));
  or_1446_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_1444_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1645_nl <= MUX_s_1_2_2(or_1444_nl, mux_tmp_1644, fsm_output(4));
  mux_1646_nl <= MUX_s_1_2_2(or_1446_nl, mux_1645_nl, fsm_output(7));
  or_1440_nl <= (fsm_output(7)) OR mux_tmp_1643;
  mux_1647_nl <= MUX_s_1_2_2(mux_1646_nl, or_1440_nl, fsm_output(2));
  or_1433_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_1432_nl <= (fsm_output(4)) OR mux_tmp_1638;
  mux_1639_nl <= MUX_s_1_2_2(or_1433_nl, or_1432_nl, fsm_output(7));
  or_1425_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1634_nl <= MUX_s_1_2_2(or_1425_nl, or_tmp_1367, fsm_output(5));
  mux_1635_nl <= MUX_s_1_2_2(or_tmp_1370, mux_1634_nl, fsm_output(4));
  or_1422_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1636_nl <= MUX_s_1_2_2(mux_1635_nl, or_1422_nl, fsm_output(7));
  mux_1640_nl <= MUX_s_1_2_2(mux_1639_nl, mux_1636_nl, fsm_output(2));
  mux_1648_nl <= MUX_s_1_2_2(mux_1647_nl, mux_1640_nl, fsm_output(1));
  or_1421_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  mux_1674_nl <= MUX_s_1_2_2(mux_1673_nl, mux_1648_nl, or_1421_nl);
  vec_rsc_0_8_i_wea_d_pff <= NOT mux_1674_nl;
  nor_950_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1494_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_949_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_951_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1701_nl <= MUX_s_1_2_2(nor_950_cse, nor_951_nl, fsm_output(0));
  mux_1702_nl <= MUX_s_1_2_2(nor_949_nl, mux_1701_nl, fsm_output(8));
  and_627_nl <= nor_223_cse AND mux_1702_nl;
  or_1522_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1521_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1699_nl <= MUX_s_1_2_2(or_1522_nl, or_1521_nl, fsm_output(0));
  nor_952_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1699_nl);
  nor_953_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_954_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1698_nl <= MUX_s_1_2_2(nor_953_nl, nor_954_nl, fsm_output(7));
  mux_1700_nl <= MUX_s_1_2_2(nor_952_nl, mux_1698_nl, fsm_output(6));
  mux_1703_nl <= MUX_s_1_2_2(and_627_nl, mux_1700_nl, fsm_output(5));
  nor_955_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_1513_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1511_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1694_nl <= MUX_s_1_2_2(or_1513_nl, or_1511_nl, fsm_output(0));
  nor_956_nl <= NOT((fsm_output(8)) OR mux_1694_nl);
  nor_957_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1695_nl <= MUX_s_1_2_2(nor_956_nl, nor_957_nl, fsm_output(7));
  mux_1696_nl <= MUX_s_1_2_2(nor_955_nl, mux_1695_nl, fsm_output(6));
  nor_958_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_959_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR
      (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_960_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1691_nl <= MUX_s_1_2_2(nor_960_nl, nor_950_cse, fsm_output(0));
  mux_1692_nl <= MUX_s_1_2_2(nor_959_nl, mux_1691_nl, fsm_output(8));
  and_628_nl <= (fsm_output(7)) AND mux_1692_nl;
  mux_1693_nl <= MUX_s_1_2_2(nor_958_nl, and_628_nl, fsm_output(6));
  mux_1697_nl <= MUX_s_1_2_2(mux_1696_nl, mux_1693_nl, fsm_output(5));
  mux_1704_nl <= MUX_s_1_2_2(mux_1703_nl, mux_1697_nl, fsm_output(2));
  or_1502_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1501_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1687_nl <= MUX_s_1_2_2(or_1502_nl, or_1501_nl, fsm_output(0));
  or_1500_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1498_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (VEC_LOOP_j_sva_11_0(2)) OR
      (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  mux_1686_nl <= MUX_s_1_2_2(or_1500_nl, or_1498_nl, fsm_output(0));
  mux_1688_nl <= MUX_s_1_2_2(mux_1687_nl, mux_1686_nl, fsm_output(8));
  nor_962_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1688_nl);
  nor_963_nl <= NOT((fsm_output(8)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1493_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1683_nl <= MUX_s_1_2_2(or_1494_cse, or_1493_nl, fsm_output(0));
  nor_964_nl <= NOT((fsm_output(8)) OR mux_1683_nl);
  mux_1684_nl <= MUX_s_1_2_2(nor_963_nl, nor_964_nl, fsm_output(7));
  nor_965_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_966_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1682_nl <= MUX_s_1_2_2(nor_965_nl, nor_966_nl, fsm_output(7));
  mux_1685_nl <= MUX_s_1_2_2(mux_1684_nl, mux_1682_nl, fsm_output(6));
  mux_1689_nl <= MUX_s_1_2_2(nor_962_nl, mux_1685_nl, fsm_output(5));
  or_1487_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1485_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1678_nl <= MUX_s_1_2_2(or_1485_nl, or_1494_cse, fsm_output(0));
  mux_1679_nl <= MUX_s_1_2_2(or_1487_nl, mux_1678_nl, fsm_output(8));
  or_1482_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1680_nl <= MUX_s_1_2_2(mux_1679_nl, or_1482_nl, fsm_output(7));
  nor_967_nl <= NOT((fsm_output(6)) OR mux_1680_nl);
  nor_968_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_969_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_970_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1675_nl <= MUX_s_1_2_2(nor_969_nl, nor_970_nl, fsm_output(0));
  mux_1676_nl <= MUX_s_1_2_2(nor_968_nl, mux_1675_nl, fsm_output(8));
  and_629_nl <= (fsm_output(7)) AND mux_1676_nl;
  nor_971_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1677_nl <= MUX_s_1_2_2(and_629_nl, nor_971_nl, fsm_output(6));
  mux_1681_nl <= MUX_s_1_2_2(nor_967_nl, mux_1677_nl, fsm_output(5));
  mux_1690_nl <= MUX_s_1_2_2(mux_1689_nl, mux_1681_nl, fsm_output(2));
  vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1704_nl, mux_1690_nl,
      fsm_output(4));
  or_1582_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_1580_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1742_nl <= MUX_s_1_2_2(or_1580_nl, mux_tmp_1728, fsm_output(4));
  mux_1743_nl <= MUX_s_1_2_2(or_1582_nl, mux_1742_nl, fsm_output(7));
  or_1579_nl <= (fsm_output(7)) OR mux_tmp_1726;
  mux_1744_nl <= MUX_s_1_2_2(mux_1743_nl, or_1579_nl, fsm_output(2));
  or_1578_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_1577_nl <= (fsm_output(4)) OR mux_tmp_1715;
  mux_1740_nl <= MUX_s_1_2_2(or_1578_nl, or_1577_nl, fsm_output(7));
  or_1576_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1737_nl <= MUX_s_1_2_2(or_1576_nl, or_tmp_1478, fsm_output(5));
  mux_1738_nl <= MUX_s_1_2_2(or_tmp_1482, mux_1737_nl, fsm_output(4));
  or_1575_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1739_nl <= MUX_s_1_2_2(mux_1738_nl, or_1575_nl, fsm_output(7));
  mux_1741_nl <= MUX_s_1_2_2(mux_1740_nl, mux_1739_nl, fsm_output(2));
  mux_1745_nl <= MUX_s_1_2_2(mux_1744_nl, mux_1741_nl, fsm_output(1));
  or_1574_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1732_nl <= MUX_s_1_2_2(or_1574_nl, or_622_cse, fsm_output(5));
  mux_1733_nl <= MUX_s_1_2_2(mux_1732_nl, or_621_cse, fsm_output(4));
  or_1565_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(3)) OR
      (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1729_nl <= MUX_s_1_2_2(or_617_cse, or_1565_nl, fsm_output(5));
  mux_1730_nl <= MUX_s_1_2_2(mux_1729_nl, mux_tmp_1728, fsm_output(4));
  mux_1734_nl <= MUX_s_1_2_2(mux_1733_nl, mux_1730_nl, fsm_output(7));
  mux_1727_nl <= MUX_s_1_2_2(mux_tmp_1726, mux_1088_cse, fsm_output(7));
  mux_1735_nl <= MUX_s_1_2_2(mux_1734_nl, mux_1727_nl, fsm_output(2));
  or_1546_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1717_nl <= MUX_s_1_2_2(or_607_cse, or_1546_nl, fsm_output(5));
  mux_1718_nl <= MUX_s_1_2_2(or_609_cse, mux_1717_nl, fsm_output(4));
  mux_1716_nl <= MUX_s_1_2_2(mux_tmp_1715, nand_25_cse, fsm_output(4));
  mux_1719_nl <= MUX_s_1_2_2(mux_1718_nl, mux_1716_nl, fsm_output(7));
  or_1537_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1709_nl <= MUX_s_1_2_2(or_1537_nl, or_601_cse, fsm_output(0));
  mux_1710_nl <= MUX_s_1_2_2(mux_1709_nl, or_tmp_1478, fsm_output(5));
  mux_1711_nl <= MUX_s_1_2_2(or_tmp_1482, mux_1710_nl, fsm_output(4));
  or_1530_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1707_nl <= MUX_s_1_2_2(mux_1073_cse, or_1530_nl, fsm_output(5));
  mux_1708_nl <= MUX_s_1_2_2(mux_1707_nl, or_596_cse, fsm_output(4));
  mux_1712_nl <= MUX_s_1_2_2(mux_1711_nl, mux_1708_nl, fsm_output(7));
  mux_1720_nl <= MUX_s_1_2_2(mux_1719_nl, mux_1712_nl, fsm_output(2));
  mux_1736_nl <= MUX_s_1_2_2(mux_1735_nl, mux_1720_nl, fsm_output(1));
  nor_252_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")));
  mux_1746_nl <= MUX_s_1_2_2(mux_1745_nl, mux_1736_nl, nor_252_nl);
  vec_rsc_0_9_i_wea_d_pff <= NOT mux_1746_nl;
  nor_925_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1600_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_924_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_926_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1773_nl <= MUX_s_1_2_2(nor_925_cse, nor_926_nl, fsm_output(0));
  mux_1774_nl <= MUX_s_1_2_2(nor_924_nl, mux_1773_nl, fsm_output(8));
  and_624_nl <= nor_223_cse AND mux_1774_nl;
  or_1628_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1627_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1771_nl <= MUX_s_1_2_2(or_1628_nl, or_1627_nl, fsm_output(0));
  nor_927_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1771_nl);
  nor_928_nl <= NOT((NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_929_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1770_nl <= MUX_s_1_2_2(nor_928_nl, nor_929_nl, fsm_output(7));
  mux_1772_nl <= MUX_s_1_2_2(nor_927_nl, mux_1770_nl, fsm_output(6));
  mux_1775_nl <= MUX_s_1_2_2(and_624_nl, mux_1772_nl, fsm_output(5));
  nor_930_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_1619_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1617_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1766_nl <= MUX_s_1_2_2(or_1619_nl, or_1617_nl, fsm_output(0));
  nor_931_nl <= NOT((fsm_output(8)) OR mux_1766_nl);
  nor_932_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1767_nl <= MUX_s_1_2_2(nor_931_nl, nor_932_nl, fsm_output(7));
  mux_1768_nl <= MUX_s_1_2_2(nor_930_nl, mux_1767_nl, fsm_output(6));
  nor_933_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_934_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR
      (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_935_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1763_nl <= MUX_s_1_2_2(nor_935_nl, nor_925_cse, fsm_output(0));
  mux_1764_nl <= MUX_s_1_2_2(nor_934_nl, mux_1763_nl, fsm_output(8));
  and_625_nl <= (fsm_output(7)) AND mux_1764_nl;
  mux_1765_nl <= MUX_s_1_2_2(nor_933_nl, and_625_nl, fsm_output(6));
  mux_1769_nl <= MUX_s_1_2_2(mux_1768_nl, mux_1765_nl, fsm_output(5));
  mux_1776_nl <= MUX_s_1_2_2(mux_1775_nl, mux_1769_nl, fsm_output(2));
  or_1608_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1607_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1759_nl <= MUX_s_1_2_2(or_1608_nl, or_1607_nl, fsm_output(0));
  or_1606_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1604_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (VEC_LOOP_j_sva_11_0(2)) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1758_nl <= MUX_s_1_2_2(or_1606_nl, or_1604_nl, fsm_output(0));
  mux_1760_nl <= MUX_s_1_2_2(mux_1759_nl, mux_1758_nl, fsm_output(8));
  nor_937_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1760_nl);
  nor_938_nl <= NOT((fsm_output(8)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1599_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1755_nl <= MUX_s_1_2_2(or_1600_cse, or_1599_nl, fsm_output(0));
  nor_939_nl <= NOT((fsm_output(8)) OR mux_1755_nl);
  mux_1756_nl <= MUX_s_1_2_2(nor_938_nl, nor_939_nl, fsm_output(7));
  nor_940_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_941_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1754_nl <= MUX_s_1_2_2(nor_940_nl, nor_941_nl, fsm_output(7));
  mux_1757_nl <= MUX_s_1_2_2(mux_1756_nl, mux_1754_nl, fsm_output(6));
  mux_1761_nl <= MUX_s_1_2_2(nor_937_nl, mux_1757_nl, fsm_output(5));
  or_1593_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1591_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1750_nl <= MUX_s_1_2_2(or_1591_nl, or_1600_cse, fsm_output(0));
  mux_1751_nl <= MUX_s_1_2_2(or_1593_nl, mux_1750_nl, fsm_output(8));
  or_1588_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1752_nl <= MUX_s_1_2_2(mux_1751_nl, or_1588_nl, fsm_output(7));
  nor_942_nl <= NOT((fsm_output(6)) OR mux_1752_nl);
  nor_943_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_944_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_945_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1747_nl <= MUX_s_1_2_2(nor_944_nl, nor_945_nl, fsm_output(0));
  mux_1748_nl <= MUX_s_1_2_2(nor_943_nl, mux_1747_nl, fsm_output(8));
  and_626_nl <= (fsm_output(7)) AND mux_1748_nl;
  nor_946_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1749_nl <= MUX_s_1_2_2(and_626_nl, nor_946_nl, fsm_output(6));
  mux_1753_nl <= MUX_s_1_2_2(nor_942_nl, mux_1749_nl, fsm_output(5));
  mux_1762_nl <= MUX_s_1_2_2(mux_1761_nl, mux_1753_nl, fsm_output(2));
  vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1776_nl, mux_1762_nl,
      fsm_output(4));
  or_1689_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT (fsm_output(3))) OR
      (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1813_nl <= MUX_s_1_2_2(or_1689_nl, or_622_cse, fsm_output(5));
  mux_1814_nl <= MUX_s_1_2_2(mux_1813_nl, or_621_cse, fsm_output(4));
  or_1680_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1810_nl <= MUX_s_1_2_2(or_617_cse, or_1680_nl, fsm_output(5));
  mux_1811_nl <= MUX_s_1_2_2(mux_1810_nl, mux_tmp_1788, fsm_output(4));
  mux_1815_nl <= MUX_s_1_2_2(mux_1814_nl, mux_1811_nl, fsm_output(7));
  mux_1809_nl <= MUX_s_1_2_2(mux_tmp_1787, mux_1088_cse, fsm_output(7));
  mux_1816_nl <= MUX_s_1_2_2(mux_1815_nl, mux_1809_nl, fsm_output(2));
  or_1670_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1802_nl <= MUX_s_1_2_2(or_607_cse, or_1670_nl, fsm_output(5));
  mux_1803_nl <= MUX_s_1_2_2(or_609_cse, mux_1802_nl, fsm_output(4));
  mux_1801_nl <= MUX_s_1_2_2(mux_tmp_1782, nand_25_cse, fsm_output(4));
  mux_1804_nl <= MUX_s_1_2_2(mux_1803_nl, mux_1801_nl, fsm_output(7));
  or_1667_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1796_nl <= MUX_s_1_2_2(or_1667_nl, or_601_cse, fsm_output(0));
  mux_1797_nl <= MUX_s_1_2_2(mux_1796_nl, or_tmp_1580, fsm_output(5));
  mux_1798_nl <= MUX_s_1_2_2(or_tmp_1583, mux_1797_nl, fsm_output(4));
  or_1662_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1794_nl <= MUX_s_1_2_2(mux_1073_cse, or_1662_nl, fsm_output(5));
  mux_1795_nl <= MUX_s_1_2_2(mux_1794_nl, or_596_cse, fsm_output(4));
  mux_1799_nl <= MUX_s_1_2_2(mux_1798_nl, mux_1795_nl, fsm_output(7));
  mux_1805_nl <= MUX_s_1_2_2(mux_1804_nl, mux_1799_nl, fsm_output(2));
  mux_1817_nl <= MUX_s_1_2_2(mux_1816_nl, mux_1805_nl, fsm_output(1));
  or_1659_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_1657_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1789_nl <= MUX_s_1_2_2(or_1657_nl, mux_tmp_1788, fsm_output(4));
  mux_1790_nl <= MUX_s_1_2_2(or_1659_nl, mux_1789_nl, fsm_output(7));
  or_1653_nl <= (fsm_output(7)) OR mux_tmp_1787;
  mux_1791_nl <= MUX_s_1_2_2(mux_1790_nl, or_1653_nl, fsm_output(2));
  or_1646_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_1645_nl <= (fsm_output(4)) OR mux_tmp_1782;
  mux_1783_nl <= MUX_s_1_2_2(or_1646_nl, or_1645_nl, fsm_output(7));
  or_1638_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1778_nl <= MUX_s_1_2_2(or_1638_nl, or_tmp_1580, fsm_output(5));
  mux_1779_nl <= MUX_s_1_2_2(or_tmp_1583, mux_1778_nl, fsm_output(4));
  or_1635_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1780_nl <= MUX_s_1_2_2(mux_1779_nl, or_1635_nl, fsm_output(7));
  mux_1784_nl <= MUX_s_1_2_2(mux_1783_nl, mux_1780_nl, fsm_output(2));
  mux_1792_nl <= MUX_s_1_2_2(mux_1791_nl, mux_1784_nl, fsm_output(1));
  or_1634_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  mux_1818_nl <= MUX_s_1_2_2(mux_1817_nl, mux_1792_nl, or_1634_nl);
  vec_rsc_0_10_i_wea_d_pff <= NOT mux_1818_nl;
  nor_900_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1707_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_899_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_901_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1845_nl <= MUX_s_1_2_2(nor_900_cse, nor_901_nl, fsm_output(0));
  mux_1846_nl <= MUX_s_1_2_2(nor_899_nl, mux_1845_nl, fsm_output(8));
  and_621_nl <= nor_223_cse AND mux_1846_nl;
  or_1735_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1734_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1843_nl <= MUX_s_1_2_2(or_1735_nl, or_1734_nl, fsm_output(0));
  nor_902_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1843_nl);
  nor_903_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_904_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1842_nl <= MUX_s_1_2_2(nor_903_nl, nor_904_nl, fsm_output(7));
  mux_1844_nl <= MUX_s_1_2_2(nor_902_nl, mux_1842_nl, fsm_output(6));
  mux_1847_nl <= MUX_s_1_2_2(and_621_nl, mux_1844_nl, fsm_output(5));
  nor_905_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("101")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_1726_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1724_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1838_nl <= MUX_s_1_2_2(or_1726_nl, or_1724_nl, fsm_output(0));
  nor_906_nl <= NOT((fsm_output(8)) OR mux_1838_nl);
  nor_907_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1839_nl <= MUX_s_1_2_2(nor_906_nl, nor_907_nl, fsm_output(7));
  mux_1840_nl <= MUX_s_1_2_2(nor_905_nl, mux_1839_nl, fsm_output(6));
  nor_908_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_909_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_910_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1835_nl <= MUX_s_1_2_2(nor_910_nl, nor_900_cse, fsm_output(0));
  mux_1836_nl <= MUX_s_1_2_2(nor_909_nl, mux_1835_nl, fsm_output(8));
  and_622_nl <= (fsm_output(7)) AND mux_1836_nl;
  mux_1837_nl <= MUX_s_1_2_2(nor_908_nl, and_622_nl, fsm_output(6));
  mux_1841_nl <= MUX_s_1_2_2(mux_1840_nl, mux_1837_nl, fsm_output(5));
  mux_1848_nl <= MUX_s_1_2_2(mux_1847_nl, mux_1841_nl, fsm_output(2));
  or_1715_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1714_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1831_nl <= MUX_s_1_2_2(or_1715_nl, or_1714_nl, fsm_output(0));
  or_1713_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1711_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (VEC_LOOP_j_sva_11_0(2)) OR
      (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT
      (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1830_nl <= MUX_s_1_2_2(or_1713_nl, or_1711_nl, fsm_output(0));
  mux_1832_nl <= MUX_s_1_2_2(mux_1831_nl, mux_1830_nl, fsm_output(8));
  nor_912_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1832_nl);
  nor_913_nl <= NOT((fsm_output(8)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1706_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1827_nl <= MUX_s_1_2_2(or_1707_cse, or_1706_nl, fsm_output(0));
  nor_914_nl <= NOT((fsm_output(8)) OR mux_1827_nl);
  mux_1828_nl <= MUX_s_1_2_2(nor_913_nl, nor_914_nl, fsm_output(7));
  nor_915_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(9))
      OR not_tmp_260);
  nor_916_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1826_nl <= MUX_s_1_2_2(nor_915_nl, nor_916_nl, fsm_output(7));
  mux_1829_nl <= MUX_s_1_2_2(mux_1828_nl, mux_1826_nl, fsm_output(6));
  mux_1833_nl <= MUX_s_1_2_2(nor_912_nl, mux_1829_nl, fsm_output(5));
  or_1700_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1698_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1822_nl <= MUX_s_1_2_2(or_1698_nl, or_1707_cse, fsm_output(0));
  mux_1823_nl <= MUX_s_1_2_2(or_1700_nl, mux_1822_nl, fsm_output(8));
  or_1695_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1824_nl <= MUX_s_1_2_2(mux_1823_nl, or_1695_nl, fsm_output(7));
  nor_917_nl <= NOT((fsm_output(6)) OR mux_1824_nl);
  nor_918_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_919_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_920_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1819_nl <= MUX_s_1_2_2(nor_919_nl, nor_920_nl, fsm_output(0));
  mux_1820_nl <= MUX_s_1_2_2(nor_918_nl, mux_1819_nl, fsm_output(8));
  and_623_nl <= (fsm_output(7)) AND mux_1820_nl;
  nor_921_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1821_nl <= MUX_s_1_2_2(and_623_nl, nor_921_nl, fsm_output(6));
  mux_1825_nl <= MUX_s_1_2_2(nor_917_nl, mux_1821_nl, fsm_output(5));
  mux_1834_nl <= MUX_s_1_2_2(mux_1833_nl, mux_1825_nl, fsm_output(2));
  vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1848_nl, mux_1834_nl,
      fsm_output(4));
  or_1795_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_1793_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1886_nl <= MUX_s_1_2_2(or_1793_nl, mux_tmp_1872, fsm_output(4));
  mux_1887_nl <= MUX_s_1_2_2(or_1795_nl, mux_1886_nl, fsm_output(7));
  or_1792_nl <= (fsm_output(7)) OR mux_tmp_1870;
  mux_1888_nl <= MUX_s_1_2_2(mux_1887_nl, or_1792_nl, fsm_output(2));
  nand_319_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  or_1790_nl <= (fsm_output(4)) OR mux_tmp_1859;
  mux_1884_nl <= MUX_s_1_2_2(nand_319_nl, or_1790_nl, fsm_output(7));
  or_1789_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1881_nl <= MUX_s_1_2_2(or_1789_nl, or_tmp_1691, fsm_output(5));
  mux_1882_nl <= MUX_s_1_2_2(or_tmp_1695, mux_1881_nl, fsm_output(4));
  or_1788_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1883_nl <= MUX_s_1_2_2(mux_1882_nl, or_1788_nl, fsm_output(7));
  mux_1885_nl <= MUX_s_1_2_2(mux_1884_nl, mux_1883_nl, fsm_output(2));
  mux_1889_nl <= MUX_s_1_2_2(mux_1888_nl, mux_1885_nl, fsm_output(1));
  or_1787_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_1876_nl <= MUX_s_1_2_2(or_1787_nl, or_622_cse, fsm_output(5));
  mux_1877_nl <= MUX_s_1_2_2(mux_1876_nl, or_621_cse, fsm_output(4));
  or_1778_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(3)) OR
      (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_1873_nl <= MUX_s_1_2_2(or_617_cse, or_1778_nl, fsm_output(5));
  mux_1874_nl <= MUX_s_1_2_2(mux_1873_nl, mux_tmp_1872, fsm_output(4));
  mux_1878_nl <= MUX_s_1_2_2(mux_1877_nl, mux_1874_nl, fsm_output(7));
  mux_1871_nl <= MUX_s_1_2_2(mux_tmp_1870, mux_1088_cse, fsm_output(7));
  mux_1879_nl <= MUX_s_1_2_2(mux_1878_nl, mux_1871_nl, fsm_output(2));
  nand_321_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  mux_1861_nl <= MUX_s_1_2_2(or_607_cse, nand_321_nl, fsm_output(5));
  mux_1862_nl <= MUX_s_1_2_2(or_609_cse, mux_1861_nl, fsm_output(4));
  mux_1860_nl <= MUX_s_1_2_2(mux_tmp_1859, nand_25_cse, fsm_output(4));
  mux_1863_nl <= MUX_s_1_2_2(mux_1862_nl, mux_1860_nl, fsm_output(7));
  or_1750_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1853_nl <= MUX_s_1_2_2(or_1750_nl, or_601_cse, fsm_output(0));
  mux_1854_nl <= MUX_s_1_2_2(mux_1853_nl, or_tmp_1691, fsm_output(5));
  mux_1855_nl <= MUX_s_1_2_2(or_tmp_1695, mux_1854_nl, fsm_output(4));
  or_1743_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1851_nl <= MUX_s_1_2_2(mux_1073_cse, or_1743_nl, fsm_output(5));
  mux_1852_nl <= MUX_s_1_2_2(mux_1851_nl, or_596_cse, fsm_output(4));
  mux_1856_nl <= MUX_s_1_2_2(mux_1855_nl, mux_1852_nl, fsm_output(7));
  mux_1864_nl <= MUX_s_1_2_2(mux_1863_nl, mux_1856_nl, fsm_output(2));
  mux_1880_nl <= MUX_s_1_2_2(mux_1879_nl, mux_1864_nl, fsm_output(1));
  and_620_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  mux_1890_nl <= MUX_s_1_2_2(mux_1889_nl, mux_1880_nl, and_620_nl);
  vec_rsc_0_11_i_wea_d_pff <= NOT mux_1890_nl;
  nor_877_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1813_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_876_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_878_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1917_nl <= MUX_s_1_2_2(nor_877_cse, nor_878_nl, fsm_output(0));
  mux_1918_nl <= MUX_s_1_2_2(nor_876_nl, mux_1917_nl, fsm_output(8));
  and_615_nl <= nor_223_cse AND mux_1918_nl;
  nand_316_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10))));
  or_1840_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1915_nl <= MUX_s_1_2_2(nand_316_nl, or_1840_nl, fsm_output(0));
  nor_879_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1915_nl);
  nor_880_nl <= NOT((NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_881_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1914_nl <= MUX_s_1_2_2(nor_880_nl, nor_881_nl, fsm_output(7));
  mux_1916_nl <= MUX_s_1_2_2(nor_879_nl, mux_1914_nl, fsm_output(6));
  mux_1919_nl <= MUX_s_1_2_2(and_615_nl, mux_1916_nl, fsm_output(5));
  and_616_nl <= (fsm_output(7)) AND (NOT (fsm_output(8))) AND (fsm_output(0)) AND
      (VEC_LOOP_j_sva_11_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("101")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3))
      AND (fsm_output(9)) AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  or_1832_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1830_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1910_nl <= MUX_s_1_2_2(or_1832_nl, or_1830_nl, fsm_output(0));
  nor_882_nl <= NOT((fsm_output(8)) OR mux_1910_nl);
  nor_883_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1911_nl <= MUX_s_1_2_2(nor_882_nl, nor_883_nl, fsm_output(7));
  mux_1912_nl <= MUX_s_1_2_2(and_616_nl, mux_1911_nl, fsm_output(6));
  nor_884_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  and_827_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(0)) AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (VEC_LOOP_j_sva_11_0(1)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(1))) AND (fsm_output(10));
  nor_886_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1907_nl <= MUX_s_1_2_2(nor_886_nl, nor_877_cse, fsm_output(0));
  mux_1908_nl <= MUX_s_1_2_2(and_827_nl, mux_1907_nl, fsm_output(8));
  and_617_nl <= (fsm_output(7)) AND mux_1908_nl;
  mux_1909_nl <= MUX_s_1_2_2(nor_884_nl, and_617_nl, fsm_output(6));
  mux_1913_nl <= MUX_s_1_2_2(mux_1912_nl, mux_1909_nl, fsm_output(5));
  mux_1920_nl <= MUX_s_1_2_2(mux_1919_nl, mux_1913_nl, fsm_output(2));
  or_1821_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1820_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1903_nl <= MUX_s_1_2_2(or_1821_nl, or_1820_nl, fsm_output(0));
  or_1819_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1817_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (VEC_LOOP_j_sva_11_0(2)) OR
      (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1902_nl <= MUX_s_1_2_2(or_1819_nl, or_1817_nl, fsm_output(0));
  mux_1904_nl <= MUX_s_1_2_2(mux_1903_nl, mux_1902_nl, fsm_output(8));
  nor_888_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1904_nl);
  nor_889_nl <= NOT((fsm_output(8)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1812_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1899_nl <= MUX_s_1_2_2(or_1813_cse, or_1812_nl, fsm_output(0));
  nor_890_nl <= NOT((fsm_output(8)) OR mux_1899_nl);
  mux_1900_nl <= MUX_s_1_2_2(nor_889_nl, nor_890_nl, fsm_output(7));
  nor_891_nl <= NOT((NOT((fsm_output(8)) AND (fsm_output(0)) AND (fsm_output(3))
      AND CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1011")) AND (NOT (fsm_output(9)))))
      OR not_tmp_260);
  nor_892_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1898_nl <= MUX_s_1_2_2(nor_891_nl, nor_892_nl, fsm_output(7));
  mux_1901_nl <= MUX_s_1_2_2(mux_1900_nl, mux_1898_nl, fsm_output(6));
  mux_1905_nl <= MUX_s_1_2_2(nor_888_nl, mux_1901_nl, fsm_output(5));
  nand_415_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(0))) AND (fsm_output(3))
      AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (fsm_output(10)));
  or_1804_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1894_nl <= MUX_s_1_2_2(or_1804_nl, or_1813_cse, fsm_output(0));
  mux_1895_nl <= MUX_s_1_2_2(nand_415_nl, mux_1894_nl, fsm_output(8));
  or_1801_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1896_nl <= MUX_s_1_2_2(mux_1895_nl, or_1801_nl, fsm_output(7));
  nor_893_nl <= NOT((fsm_output(6)) OR mux_1896_nl);
  nor_894_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  and_619_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  nor_895_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1891_nl <= MUX_s_1_2_2(and_619_nl, nor_895_nl, fsm_output(0));
  mux_1892_nl <= MUX_s_1_2_2(nor_894_nl, mux_1891_nl, fsm_output(8));
  and_618_nl <= (fsm_output(7)) AND mux_1892_nl;
  nor_896_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1893_nl <= MUX_s_1_2_2(and_618_nl, nor_896_nl, fsm_output(6));
  mux_1897_nl <= MUX_s_1_2_2(nor_893_nl, mux_1893_nl, fsm_output(5));
  mux_1906_nl <= MUX_s_1_2_2(mux_1905_nl, mux_1897_nl, fsm_output(2));
  vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1920_nl, mux_1906_nl,
      fsm_output(4));
  or_1905_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(4)) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  or_1903_nl <= (NOT (fsm_output(0))) OR (fsm_output(4)) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_1958_nl <= MUX_s_1_2_2(or_1905_nl, or_1903_nl, fsm_output(5));
  nand_311_nl <= NOT((fsm_output(4)) AND (fsm_output(9)) AND (fsm_output(3)) AND
      (fsm_output(6)) AND (NOT (fsm_output(10))));
  or_1900_nl <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (fsm_output(3)) OR not_tmp_378;
  mux_1957_nl <= MUX_s_1_2_2(nand_311_nl, or_1900_nl, fsm_output(0));
  or_1902_nl <= (fsm_output(5)) OR mux_1957_nl;
  mux_1959_nl <= MUX_s_1_2_2(mux_1958_nl, or_1902_nl, fsm_output(8));
  or_1898_nl <= (fsm_output(4)) OR (NOT (fsm_output(9))) OR (fsm_output(3)) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  or_1896_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(4))) OR (fsm_output(9)) OR not_tmp_381;
  mux_1954_nl <= MUX_s_1_2_2(or_1898_nl, or_1896_nl, fsm_output(0));
  mux_1955_nl <= MUX_s_1_2_2(mux_1954_nl, or_tmp_1812, fsm_output(5));
  mux_1956_nl <= MUX_s_1_2_2(mux_1955_nl, or_tmp_1811, fsm_output(8));
  mux_1960_nl <= MUX_s_1_2_2(mux_1959_nl, mux_1956_nl, fsm_output(7));
  nand_437_nl <= NOT((fsm_output(0)) AND (fsm_output(4)) AND (fsm_output(9)) AND
      (fsm_output(3)) AND (NOT (fsm_output(6))) AND (fsm_output(10)));
  or_1891_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_1951_nl <= MUX_s_1_2_2(or_tmp_1821, or_1891_nl, fsm_output(0));
  mux_1952_nl <= MUX_s_1_2_2(nand_437_nl, mux_1951_nl, fsm_output(5));
  or_1894_nl <= (fsm_output(8)) OR mux_1952_nl;
  or_1890_nl <= (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (fsm_output(4)) OR (fsm_output(9))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(10));
  or_1889_nl <= (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_1888_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_1948_nl <= MUX_s_1_2_2(or_1889_nl, or_1888_nl, fsm_output(0));
  mux_1949_nl <= MUX_s_1_2_2(or_1890_nl, mux_1948_nl, fsm_output(5));
  mux_1950_nl <= MUX_s_1_2_2(mux_1949_nl, nand_tmp_74, fsm_output(8));
  mux_1953_nl <= MUX_s_1_2_2(or_1894_nl, mux_1950_nl, fsm_output(7));
  mux_1961_nl <= MUX_s_1_2_2(mux_1960_nl, mux_1953_nl, fsm_output(1));
  or_1887_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(4))) OR (fsm_output(9))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(10));
  or_1886_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(9)) OR not_tmp_381;
  mux_1944_nl <= MUX_s_1_2_2(or_1887_nl, or_1886_nl, fsm_output(5));
  or_1884_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(9)) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_1883_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_1943_nl <= MUX_s_1_2_2(or_1884_nl, or_1883_nl, fsm_output(5));
  mux_1945_nl <= MUX_s_1_2_2(mux_1944_nl, mux_1943_nl, fsm_output(8));
  mux_1946_nl <= MUX_s_1_2_2(mux_tmp_1927, mux_1945_nl, fsm_output(7));
  or_1882_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(4))) OR (fsm_output(9))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_1881_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(4))) OR (fsm_output(9)) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  mux_1940_nl <= MUX_s_1_2_2(or_1882_nl, or_1881_nl, fsm_output(5));
  mux_1941_nl <= MUX_s_1_2_2(or_tmp_1797, mux_1940_nl, fsm_output(8));
  or_1879_nl <= (fsm_output(4)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (fsm_output(10));
  mux_1937_nl <= MUX_s_1_2_2(or_1879_nl, or_tmp_1821, fsm_output(0));
  or_1876_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(4)) OR (fsm_output(9)) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_1938_nl <= MUX_s_1_2_2(mux_1937_nl, or_1876_nl, fsm_output(5));
  or_1875_nl <= (NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (fsm_output(4)))
      OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_1939_nl <= MUX_s_1_2_2(mux_1938_nl, or_1875_nl, fsm_output(8));
  mux_1942_nl <= MUX_s_1_2_2(mux_1941_nl, mux_1939_nl, fsm_output(7));
  mux_1947_nl <= MUX_s_1_2_2(mux_1946_nl, mux_1942_nl, fsm_output(1));
  mux_1962_nl <= MUX_s_1_2_2(mux_1961_nl, mux_1947_nl, fsm_output(2));
  or_1873_nl <= (fsm_output(8)) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(4)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(10)));
  or_1871_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(4))) OR (fsm_output(9))
      OR not_tmp_381;
  mux_1932_nl <= MUX_s_1_2_2(or_1871_nl, or_tmp_1812, fsm_output(5));
  mux_1933_nl <= MUX_s_1_2_2(mux_1932_nl, or_tmp_1811, fsm_output(8));
  mux_1934_nl <= MUX_s_1_2_2(or_1873_nl, mux_1933_nl, fsm_output(7));
  or_1867_nl <= (fsm_output(8)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(10));
  or_1866_nl <= (fsm_output(5)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (fsm_output(0))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR
      (fsm_output(4)) OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(6)) OR
      (fsm_output(10));
  mux_1930_nl <= MUX_s_1_2_2(or_1866_nl, nand_tmp_74, fsm_output(8));
  mux_1931_nl <= MUX_s_1_2_2(or_1867_nl, mux_1930_nl, fsm_output(7));
  mux_1935_nl <= MUX_s_1_2_2(mux_1934_nl, mux_1931_nl, fsm_output(1));
  or_1862_nl <= (fsm_output(7)) OR mux_tmp_1927;
  or_1850_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT (fsm_output(4))) OR (fsm_output(9))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(10)));
  mux_1923_nl <= MUX_s_1_2_2(or_tmp_1797, or_1850_nl, fsm_output(8));
  or_1848_nl <= (fsm_output(8)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (NOT (fsm_output(0))) OR (fsm_output(4))
      OR (fsm_output(9)) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(10));
  mux_1924_nl <= MUX_s_1_2_2(mux_1923_nl, or_1848_nl, fsm_output(7));
  mux_1928_nl <= MUX_s_1_2_2(or_1862_nl, mux_1924_nl, fsm_output(1));
  mux_1936_nl <= MUX_s_1_2_2(mux_1935_nl, mux_1928_nl, fsm_output(2));
  or_1847_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"));
  mux_1963_nl <= MUX_s_1_2_2(mux_1962_nl, mux_1936_nl, or_1847_nl);
  vec_rsc_0_12_i_wea_d_pff <= NOT mux_1963_nl;
  nor_850_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_1923_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_849_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_851_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1990_nl <= MUX_s_1_2_2(nor_850_cse, nor_851_nl, fsm_output(0));
  mux_1991_nl <= MUX_s_1_2_2(nor_849_nl, mux_1990_nl, fsm_output(8));
  and_612_nl <= nor_223_cse AND mux_1991_nl;
  or_1951_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1950_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_1988_nl <= MUX_s_1_2_2(or_1951_nl, or_1950_nl, fsm_output(0));
  nor_852_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1988_nl);
  nor_853_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_854_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_1987_nl <= MUX_s_1_2_2(nor_853_nl, nor_854_nl, fsm_output(7));
  mux_1989_nl <= MUX_s_1_2_2(nor_852_nl, mux_1987_nl, fsm_output(6));
  mux_1992_nl <= MUX_s_1_2_2(and_612_nl, mux_1989_nl, fsm_output(5));
  nor_855_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("110")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  or_1942_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1940_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1983_nl <= MUX_s_1_2_2(or_1942_nl, or_1940_nl, fsm_output(0));
  nor_856_nl <= NOT((fsm_output(8)) OR mux_1983_nl);
  nor_857_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1984_nl <= MUX_s_1_2_2(nor_856_nl, nor_857_nl, fsm_output(7));
  mux_1985_nl <= MUX_s_1_2_2(nor_855_nl, mux_1984_nl, fsm_output(6));
  nor_858_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  nor_859_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR
      (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_860_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1980_nl <= MUX_s_1_2_2(nor_860_nl, nor_850_cse, fsm_output(0));
  mux_1981_nl <= MUX_s_1_2_2(nor_859_nl, mux_1980_nl, fsm_output(8));
  and_613_nl <= (fsm_output(7)) AND mux_1981_nl;
  mux_1982_nl <= MUX_s_1_2_2(nor_858_nl, and_613_nl, fsm_output(6));
  mux_1986_nl <= MUX_s_1_2_2(mux_1985_nl, mux_1982_nl, fsm_output(5));
  mux_1993_nl <= MUX_s_1_2_2(mux_1992_nl, mux_1986_nl, fsm_output(2));
  or_1931_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_1930_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1976_nl <= MUX_s_1_2_2(or_1931_nl, or_1930_nl, fsm_output(0));
  or_1929_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_1927_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_1975_nl <= MUX_s_1_2_2(or_1929_nl, or_1927_nl, fsm_output(0));
  mux_1977_nl <= MUX_s_1_2_2(mux_1976_nl, mux_1975_nl, fsm_output(8));
  nor_862_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_1977_nl);
  nor_863_nl <= NOT((fsm_output(8)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_1922_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_1972_nl <= MUX_s_1_2_2(or_1923_cse, or_1922_nl, fsm_output(0));
  nor_864_nl <= NOT((fsm_output(8)) OR mux_1972_nl);
  mux_1973_nl <= MUX_s_1_2_2(nor_863_nl, nor_864_nl, fsm_output(7));
  nor_865_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR
      (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR
      (fsm_output(9)) OR not_tmp_260);
  nor_866_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_1971_nl <= MUX_s_1_2_2(nor_865_nl, nor_866_nl, fsm_output(7));
  mux_1974_nl <= MUX_s_1_2_2(mux_1973_nl, mux_1971_nl, fsm_output(6));
  mux_1978_nl <= MUX_s_1_2_2(nor_862_nl, mux_1974_nl, fsm_output(5));
  or_1916_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_1914_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_1967_nl <= MUX_s_1_2_2(or_1914_nl, or_1923_cse, fsm_output(0));
  mux_1968_nl <= MUX_s_1_2_2(or_1916_nl, mux_1967_nl, fsm_output(8));
  or_1911_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_1969_nl <= MUX_s_1_2_2(mux_1968_nl, or_1911_nl, fsm_output(7));
  nor_867_nl <= NOT((fsm_output(6)) OR mux_1969_nl);
  nor_868_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_869_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(3))) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  nor_870_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_1964_nl <= MUX_s_1_2_2(nor_869_nl, nor_870_nl, fsm_output(0));
  mux_1965_nl <= MUX_s_1_2_2(nor_868_nl, mux_1964_nl, fsm_output(8));
  and_614_nl <= (fsm_output(7)) AND mux_1965_nl;
  nor_871_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_1966_nl <= MUX_s_1_2_2(and_614_nl, nor_871_nl, fsm_output(6));
  mux_1970_nl <= MUX_s_1_2_2(nor_867_nl, mux_1966_nl, fsm_output(5));
  mux_1979_nl <= MUX_s_1_2_2(mux_1978_nl, mux_1970_nl, fsm_output(2));
  vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1993_nl, mux_1979_nl,
      fsm_output(4));
  or_2011_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_2009_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("110")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2031_nl <= MUX_s_1_2_2(or_2009_nl, mux_tmp_2017, fsm_output(4));
  mux_2032_nl <= MUX_s_1_2_2(or_2011_nl, mux_2031_nl, fsm_output(7));
  or_2008_nl <= (fsm_output(7)) OR mux_tmp_2015;
  mux_2033_nl <= MUX_s_1_2_2(mux_2032_nl, or_2008_nl, fsm_output(2));
  nand_305_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  or_2006_nl <= (fsm_output(4)) OR mux_tmp_2004;
  mux_2029_nl <= MUX_s_1_2_2(nand_305_nl, or_2006_nl, fsm_output(7));
  or_2005_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2026_nl <= MUX_s_1_2_2(or_2005_nl, or_tmp_1907, fsm_output(5));
  mux_2027_nl <= MUX_s_1_2_2(or_tmp_1911, mux_2026_nl, fsm_output(4));
  or_2004_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_2028_nl <= MUX_s_1_2_2(mux_2027_nl, or_2004_nl, fsm_output(7));
  mux_2030_nl <= MUX_s_1_2_2(mux_2029_nl, mux_2028_nl, fsm_output(2));
  mux_2034_nl <= MUX_s_1_2_2(mux_2033_nl, mux_2030_nl, fsm_output(1));
  or_2003_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_2021_nl <= MUX_s_1_2_2(or_2003_nl, or_622_cse, fsm_output(5));
  mux_2022_nl <= MUX_s_1_2_2(mux_2021_nl, or_621_cse, fsm_output(4));
  or_1994_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(3)) OR
      (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_2018_nl <= MUX_s_1_2_2(or_617_cse, or_1994_nl, fsm_output(5));
  mux_2019_nl <= MUX_s_1_2_2(mux_2018_nl, mux_tmp_2017, fsm_output(4));
  mux_2023_nl <= MUX_s_1_2_2(mux_2022_nl, mux_2019_nl, fsm_output(7));
  mux_2016_nl <= MUX_s_1_2_2(mux_tmp_2015, mux_1088_cse, fsm_output(7));
  mux_2024_nl <= MUX_s_1_2_2(mux_2023_nl, mux_2016_nl, fsm_output(2));
  nand_307_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  mux_2006_nl <= MUX_s_1_2_2(or_607_cse, nand_307_nl, fsm_output(5));
  mux_2007_nl <= MUX_s_1_2_2(or_609_cse, mux_2006_nl, fsm_output(4));
  mux_2005_nl <= MUX_s_1_2_2(mux_tmp_2004, nand_25_cse, fsm_output(4));
  mux_2008_nl <= MUX_s_1_2_2(mux_2007_nl, mux_2005_nl, fsm_output(7));
  or_1966_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_1998_nl <= MUX_s_1_2_2(or_1966_nl, or_601_cse, fsm_output(0));
  mux_1999_nl <= MUX_s_1_2_2(mux_1998_nl, or_tmp_1907, fsm_output(5));
  mux_2000_nl <= MUX_s_1_2_2(or_tmp_1911, mux_1999_nl, fsm_output(4));
  or_1959_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_1996_nl <= MUX_s_1_2_2(mux_1073_cse, or_1959_nl, fsm_output(5));
  mux_1997_nl <= MUX_s_1_2_2(mux_1996_nl, or_596_cse, fsm_output(4));
  mux_2001_nl <= MUX_s_1_2_2(mux_2000_nl, mux_1997_nl, fsm_output(7));
  mux_2009_nl <= MUX_s_1_2_2(mux_2008_nl, mux_2001_nl, fsm_output(2));
  mux_2025_nl <= MUX_s_1_2_2(mux_2024_nl, mux_2009_nl, fsm_output(1));
  and_611_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
  mux_2035_nl <= MUX_s_1_2_2(mux_2034_nl, mux_2025_nl, and_611_nl);
  vec_rsc_0_13_i_wea_d_pff <= NOT mux_2035_nl;
  nor_827_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_2029_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_826_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_828_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2062_nl <= MUX_s_1_2_2(nor_827_cse, nor_828_nl, fsm_output(0));
  mux_2063_nl <= MUX_s_1_2_2(nor_826_nl, mux_2062_nl, fsm_output(8));
  and_606_nl <= nor_223_cse AND mux_2063_nl;
  nand_302_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10))));
  or_2056_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_2060_nl <= MUX_s_1_2_2(nand_302_nl, or_2056_nl, fsm_output(0));
  nor_829_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_2060_nl);
  nor_830_nl <= NOT((NOT (fsm_output(8))) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_831_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_2059_nl <= MUX_s_1_2_2(nor_830_nl, nor_831_nl, fsm_output(7));
  mux_2061_nl <= MUX_s_1_2_2(nor_829_nl, mux_2059_nl, fsm_output(6));
  mux_2064_nl <= MUX_s_1_2_2(and_606_nl, mux_2061_nl, fsm_output(5));
  and_607_nl <= (fsm_output(7)) AND (NOT (fsm_output(8))) AND (fsm_output(0)) AND
      (VEC_LOOP_j_sva_11_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("110")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3))
      AND (fsm_output(9)) AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  or_2048_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_2046_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_2055_nl <= MUX_s_1_2_2(or_2048_nl, or_2046_nl, fsm_output(0));
  nor_832_nl <= NOT((fsm_output(8)) OR mux_2055_nl);
  nor_833_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (VEC_LOOP_j_sva_11_0(1)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2056_nl <= MUX_s_1_2_2(nor_832_nl, nor_833_nl, fsm_output(7));
  mux_2057_nl <= MUX_s_1_2_2(and_607_nl, mux_2056_nl, fsm_output(6));
  nor_834_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  and_826_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(0)) AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (NOT (VEC_LOOP_j_sva_11_0(1))) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(1))) AND (fsm_output(10));
  nor_836_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_2052_nl <= MUX_s_1_2_2(nor_836_nl, nor_827_cse, fsm_output(0));
  mux_2053_nl <= MUX_s_1_2_2(and_826_nl, mux_2052_nl, fsm_output(8));
  and_608_nl <= (fsm_output(7)) AND mux_2053_nl;
  mux_2054_nl <= MUX_s_1_2_2(nor_834_nl, and_608_nl, fsm_output(6));
  mux_2058_nl <= MUX_s_1_2_2(mux_2057_nl, mux_2054_nl, fsm_output(5));
  mux_2065_nl <= MUX_s_1_2_2(mux_2064_nl, mux_2058_nl, fsm_output(2));
  or_2037_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_2036_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_2048_nl <= MUX_s_1_2_2(or_2037_nl, or_2036_nl, fsm_output(0));
  or_2035_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_2033_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (VEC_LOOP_j_sva_11_0(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_2047_nl <= MUX_s_1_2_2(or_2035_nl, or_2033_nl, fsm_output(0));
  mux_2049_nl <= MUX_s_1_2_2(mux_2048_nl, mux_2047_nl, fsm_output(8));
  nor_838_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_2049_nl);
  nor_839_nl <= NOT((fsm_output(8)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_2028_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_2044_nl <= MUX_s_1_2_2(or_2029_cse, or_2028_nl, fsm_output(0));
  nor_840_nl <= NOT((fsm_output(8)) OR mux_2044_nl);
  mux_2045_nl <= MUX_s_1_2_2(nor_839_nl, nor_840_nl, fsm_output(7));
  nor_841_nl <= NOT((NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(8)) AND (fsm_output(0)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_260);
  nor_842_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_2043_nl <= MUX_s_1_2_2(nor_841_nl, nor_842_nl, fsm_output(7));
  mux_2046_nl <= MUX_s_1_2_2(mux_2045_nl, mux_2043_nl, fsm_output(6));
  mux_2050_nl <= MUX_s_1_2_2(nor_838_nl, mux_2046_nl, fsm_output(5));
  nand_413_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(0))) AND (fsm_output(3))
      AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (fsm_output(10)));
  or_2020_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_2039_nl <= MUX_s_1_2_2(or_2020_nl, or_2029_cse, fsm_output(0));
  mux_2040_nl <= MUX_s_1_2_2(nand_413_nl, mux_2039_nl, fsm_output(8));
  or_2017_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_2041_nl <= MUX_s_1_2_2(mux_2040_nl, or_2017_nl, fsm_output(7));
  nor_843_nl <= NOT((fsm_output(6)) OR mux_2041_nl);
  nor_844_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  and_610_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  nor_845_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_2036_nl <= MUX_s_1_2_2(and_610_nl, nor_845_nl, fsm_output(0));
  mux_2037_nl <= MUX_s_1_2_2(nor_844_nl, mux_2036_nl, fsm_output(8));
  and_609_nl <= (fsm_output(7)) AND mux_2037_nl;
  nor_846_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2038_nl <= MUX_s_1_2_2(and_609_nl, nor_846_nl, fsm_output(6));
  mux_2042_nl <= MUX_s_1_2_2(nor_843_nl, mux_2038_nl, fsm_output(5));
  mux_2051_nl <= MUX_s_1_2_2(mux_2050_nl, mux_2042_nl, fsm_output(2));
  vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2065_nl, mux_2051_nl,
      fsm_output(4));
  or_2118_nl <= (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_2102_nl <= MUX_s_1_2_2(or_2118_nl, or_622_cse, fsm_output(5));
  mux_2103_nl <= MUX_s_1_2_2(mux_2102_nl, or_621_cse, fsm_output(4));
  or_2109_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_2099_nl <= MUX_s_1_2_2(or_617_cse, or_2109_nl, fsm_output(5));
  mux_2100_nl <= MUX_s_1_2_2(mux_2099_nl, mux_tmp_2077, fsm_output(4));
  mux_2104_nl <= MUX_s_1_2_2(mux_2103_nl, mux_2100_nl, fsm_output(7));
  mux_2098_nl <= MUX_s_1_2_2(mux_tmp_2076, mux_1088_cse, fsm_output(7));
  mux_2105_nl <= MUX_s_1_2_2(mux_2104_nl, mux_2098_nl, fsm_output(2));
  nand_297_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  mux_2091_nl <= MUX_s_1_2_2(or_607_cse, nand_297_nl, fsm_output(5));
  mux_2092_nl <= MUX_s_1_2_2(or_609_cse, mux_2091_nl, fsm_output(4));
  mux_2090_nl <= MUX_s_1_2_2(mux_tmp_2071, nand_25_cse, fsm_output(4));
  mux_2093_nl <= MUX_s_1_2_2(mux_2092_nl, mux_2090_nl, fsm_output(7));
  or_2096_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2085_nl <= MUX_s_1_2_2(or_2096_nl, or_601_cse, fsm_output(0));
  mux_2086_nl <= MUX_s_1_2_2(mux_2085_nl, or_tmp_2009, fsm_output(5));
  mux_2087_nl <= MUX_s_1_2_2(or_tmp_2012, mux_2086_nl, fsm_output(4));
  or_2091_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_2083_nl <= MUX_s_1_2_2(mux_1073_cse, or_2091_nl, fsm_output(5));
  mux_2084_nl <= MUX_s_1_2_2(mux_2083_nl, or_596_cse, fsm_output(4));
  mux_2088_nl <= MUX_s_1_2_2(mux_2087_nl, mux_2084_nl, fsm_output(7));
  mux_2094_nl <= MUX_s_1_2_2(mux_2093_nl, mux_2088_nl, fsm_output(2));
  mux_2106_nl <= MUX_s_1_2_2(mux_2105_nl, mux_2094_nl, fsm_output(1));
  or_2088_nl <= (fsm_output(4)) OR (fsm_output(5)) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_2086_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(0)) OR (VEC_LOOP_j_sva_11_0(0))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2078_nl <= MUX_s_1_2_2(or_2086_nl, mux_tmp_2077, fsm_output(4));
  mux_2079_nl <= MUX_s_1_2_2(or_2088_nl, mux_2078_nl, fsm_output(7));
  or_2082_nl <= (fsm_output(7)) OR mux_tmp_2076;
  mux_2080_nl <= MUX_s_1_2_2(mux_2079_nl, or_2082_nl, fsm_output(2));
  nand_298_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  or_2074_nl <= (fsm_output(4)) OR mux_tmp_2071;
  mux_2072_nl <= MUX_s_1_2_2(nand_298_nl, or_2074_nl, fsm_output(7));
  or_2067_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2067_nl <= MUX_s_1_2_2(or_2067_nl, or_tmp_2009, fsm_output(5));
  mux_2068_nl <= MUX_s_1_2_2(or_tmp_2012, mux_2067_nl, fsm_output(4));
  or_2064_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_2069_nl <= MUX_s_1_2_2(mux_2068_nl, or_2064_nl, fsm_output(7));
  mux_2073_nl <= MUX_s_1_2_2(mux_2072_nl, mux_2069_nl, fsm_output(2));
  mux_2081_nl <= MUX_s_1_2_2(mux_2080_nl, mux_2073_nl, fsm_output(1));
  nand_299_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110")));
  mux_2107_nl <= MUX_s_1_2_2(mux_2106_nl, mux_2081_nl, nand_299_nl);
  vec_rsc_0_14_i_wea_d_pff <= NOT mux_2107_nl;
  nor_804_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  or_2136_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10));
  nor_803_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  nor_805_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2134_nl <= MUX_s_1_2_2(nor_804_cse, nor_805_nl, fsm_output(0));
  mux_2135_nl <= MUX_s_1_2_2(nor_803_nl, mux_2134_nl, fsm_output(8));
  and_601_nl <= nor_223_cse AND mux_2135_nl;
  nand_293_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10))));
  or_2163_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260;
  mux_2132_nl <= MUX_s_1_2_2(nand_293_nl, or_2163_nl, fsm_output(0));
  nor_806_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_2132_nl);
  nor_807_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_808_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_2131_nl <= MUX_s_1_2_2(nor_807_nl, nor_808_nl, fsm_output(7));
  mux_2133_nl <= MUX_s_1_2_2(nor_806_nl, mux_2131_nl, fsm_output(6));
  mux_2136_nl <= MUX_s_1_2_2(and_601_nl, mux_2133_nl, fsm_output(5));
  and_602_nl <= (fsm_output(7)) AND (NOT (fsm_output(8))) AND (fsm_output(0)) AND
      (NOT (VEC_LOOP_j_sva_11_0(0))) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3))
      AND (fsm_output(9)) AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  or_2155_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  or_2153_nl <= (fsm_output(3)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_2127_nl <= MUX_s_1_2_2(or_2155_nl, or_2153_nl, fsm_output(0));
  nor_809_nl <= NOT((fsm_output(8)) OR mux_2127_nl);
  nor_810_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2128_nl <= MUX_s_1_2_2(nor_809_nl, nor_810_nl, fsm_output(7));
  mux_2129_nl <= MUX_s_1_2_2(and_602_nl, mux_2128_nl, fsm_output(6));
  nor_811_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  and_825_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(0)) AND (NOT (VEC_LOOP_j_sva_11_0(0))) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (VEC_LOOP_j_sva_11_0(1)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(1))) AND (fsm_output(10));
  nor_813_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_2124_nl <= MUX_s_1_2_2(nor_813_nl, nor_804_cse, fsm_output(0));
  mux_2125_nl <= MUX_s_1_2_2(and_825_nl, mux_2124_nl, fsm_output(8));
  and_603_nl <= (fsm_output(7)) AND mux_2125_nl;
  mux_2126_nl <= MUX_s_1_2_2(nor_811_nl, and_603_nl, fsm_output(6));
  mux_2130_nl <= MUX_s_1_2_2(mux_2129_nl, mux_2126_nl, fsm_output(5));
  mux_2137_nl <= MUX_s_1_2_2(mux_2136_nl, mux_2130_nl, fsm_output(2));
  or_2144_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR (NOT
      (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  or_2143_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(3))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_2120_nl <= MUX_s_1_2_2(or_2144_nl, or_2143_nl, fsm_output(0));
  or_2142_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_260;
  or_2140_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR (NOT (VEC_LOOP_j_sva_11_0(2)))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (VEC_LOOP_j_sva_11_0(1))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(1)) OR (fsm_output(10));
  mux_2119_nl <= MUX_s_1_2_2(or_2142_nl, or_2140_nl, fsm_output(0));
  mux_2121_nl <= MUX_s_1_2_2(mux_2120_nl, mux_2119_nl, fsm_output(8));
  nor_815_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_2121_nl);
  nor_816_nl <= NOT((fsm_output(8)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_2135_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_2116_nl <= MUX_s_1_2_2(or_2136_cse, or_2135_nl, fsm_output(0));
  nor_817_nl <= NOT((fsm_output(8)) OR mux_2116_nl);
  mux_2117_nl <= MUX_s_1_2_2(nor_816_nl, nor_817_nl, fsm_output(7));
  nor_818_nl <= NOT((NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(8)) AND (fsm_output(0)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_260);
  nor_819_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_11_0(0))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  mux_2115_nl <= MUX_s_1_2_2(nor_818_nl, nor_819_nl, fsm_output(7));
  mux_2118_nl <= MUX_s_1_2_2(mux_2117_nl, mux_2115_nl, fsm_output(6));
  mux_2122_nl <= MUX_s_1_2_2(nor_815_nl, mux_2118_nl, fsm_output(5));
  nand_411_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(0))) AND (fsm_output(3))
      AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (fsm_output(10)));
  or_2127_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_2111_nl <= MUX_s_1_2_2(or_2127_nl, or_2136_cse, fsm_output(0));
  mux_2112_nl <= MUX_s_1_2_2(nand_411_nl, mux_2111_nl, fsm_output(8));
  or_2124_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_2113_nl <= MUX_s_1_2_2(mux_2112_nl, or_2124_nl, fsm_output(7));
  nor_820_nl <= NOT((fsm_output(6)) OR mux_2113_nl);
  nor_821_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10)));
  and_605_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  nor_822_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (VEC_LOOP_j_sva_11_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_260);
  mux_2108_nl <= MUX_s_1_2_2(and_605_nl, nor_822_nl, fsm_output(0));
  mux_2109_nl <= MUX_s_1_2_2(nor_821_nl, mux_2108_nl, fsm_output(8));
  and_604_nl <= (fsm_output(7)) AND mux_2109_nl;
  nor_823_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2110_nl <= MUX_s_1_2_2(and_604_nl, nor_823_nl, fsm_output(6));
  mux_2114_nl <= MUX_s_1_2_2(nor_820_nl, mux_2110_nl, fsm_output(5));
  mux_2123_nl <= MUX_s_1_2_2(mux_2122_nl, mux_2114_nl, fsm_output(2));
  vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2137_nl, mux_2123_nl,
      fsm_output(4));
  or_2224_nl <= (fsm_output(4)) OR (fsm_output(5)) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10)));
  or_2222_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("111")) OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2175_nl <= MUX_s_1_2_2(or_2222_nl, mux_tmp_2161, fsm_output(4));
  mux_2176_nl <= MUX_s_1_2_2(or_2224_nl, mux_2175_nl, fsm_output(7));
  or_2221_nl <= (fsm_output(7)) OR mux_tmp_2159;
  mux_2177_nl <= MUX_s_1_2_2(mux_2176_nl, or_2221_nl, fsm_output(2));
  nand_284_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  or_2219_nl <= (fsm_output(4)) OR mux_tmp_2148;
  mux_2173_nl <= MUX_s_1_2_2(nand_284_nl, or_2219_nl, fsm_output(7));
  or_2218_nl <= (fsm_output(0)) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2170_nl <= MUX_s_1_2_2(or_2218_nl, or_tmp_2120, fsm_output(5));
  mux_2171_nl <= MUX_s_1_2_2(or_tmp_2124, mux_2170_nl, fsm_output(4));
  or_2217_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_2172_nl <= MUX_s_1_2_2(mux_2171_nl, or_2217_nl, fsm_output(7));
  mux_2174_nl <= MUX_s_1_2_2(mux_2173_nl, mux_2172_nl, fsm_output(2));
  mux_2178_nl <= MUX_s_1_2_2(mux_2177_nl, mux_2174_nl, fsm_output(1));
  nand_438_nl <= NOT((NOT (fsm_output(0))) AND (VEC_LOOP_j_sva_11_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (fsm_output(3)) AND (NOT (fsm_output(6)))
      AND (fsm_output(9)) AND (NOT (fsm_output(8))) AND (fsm_output(10)));
  mux_2165_nl <= MUX_s_1_2_2(nand_438_nl, or_622_cse, fsm_output(5));
  mux_2166_nl <= MUX_s_1_2_2(mux_2165_nl, or_621_cse, fsm_output(4));
  or_2207_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(0)) OR (NOT (VEC_LOOP_j_sva_11_0(0))) OR (fsm_output(3)) OR
      (NOT (fsm_output(6))) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_2162_nl <= MUX_s_1_2_2(or_617_cse, or_2207_nl, fsm_output(5));
  mux_2163_nl <= MUX_s_1_2_2(mux_2162_nl, mux_tmp_2161, fsm_output(4));
  mux_2167_nl <= MUX_s_1_2_2(mux_2166_nl, mux_2163_nl, fsm_output(7));
  mux_2160_nl <= MUX_s_1_2_2(mux_tmp_2159, mux_1088_cse, fsm_output(7));
  mux_2168_nl <= MUX_s_1_2_2(mux_2167_nl, mux_2160_nl, fsm_output(2));
  nand_286_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (NOT (fsm_output(10))));
  mux_2150_nl <= MUX_s_1_2_2(or_607_cse, nand_286_nl, fsm_output(5));
  mux_2151_nl <= MUX_s_1_2_2(or_609_cse, mux_2150_nl, fsm_output(4));
  mux_2149_nl <= MUX_s_1_2_2(mux_tmp_2148, nand_25_cse, fsm_output(4));
  mux_2152_nl <= MUX_s_1_2_2(mux_2151_nl, mux_2149_nl, fsm_output(7));
  or_2179_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (fsm_output(10));
  mux_2142_nl <= MUX_s_1_2_2(or_2179_nl, or_601_cse, fsm_output(0));
  mux_2143_nl <= MUX_s_1_2_2(mux_2142_nl, or_tmp_2120, fsm_output(5));
  mux_2144_nl <= MUX_s_1_2_2(or_tmp_2124, mux_2143_nl, fsm_output(4));
  or_2172_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_2140_nl <= MUX_s_1_2_2(mux_1073_cse, or_2172_nl, fsm_output(5));
  mux_2141_nl <= MUX_s_1_2_2(mux_2140_nl, or_596_cse, fsm_output(4));
  mux_2145_nl <= MUX_s_1_2_2(mux_2144_nl, mux_2141_nl, fsm_output(7));
  mux_2153_nl <= MUX_s_1_2_2(mux_2152_nl, mux_2145_nl, fsm_output(2));
  mux_2169_nl <= MUX_s_1_2_2(mux_2168_nl, mux_2153_nl, fsm_output(1));
  and_600_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_12_1_1_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
  mux_2179_nl <= MUX_s_1_2_2(mux_2178_nl, mux_2169_nl, and_600_nl);
  vec_rsc_0_15_i_wea_d_pff <= NOT mux_2179_nl;
  and_591_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111")) AND (NOT
      (fsm_output(3))) AND (fsm_output(9)) AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  nand_278_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(3)) AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (NOT
      (fsm_output(10))));
  and_823_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(0))) AND (fsm_output(3))
      AND (NOT (fsm_output(9))) AND (NOT (fsm_output(1))) AND (fsm_output(10));
  nor_786_nl <= NOT((NOT (fsm_output(3))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2206_nl <= MUX_s_1_2_2(and_591_cse, nor_786_nl, fsm_output(0));
  mux_2207_nl <= MUX_s_1_2_2(and_823_nl, mux_2206_nl, fsm_output(8));
  and_590_nl <= nor_223_cse AND mux_2207_nl;
  nand_269_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10))));
  or_2269_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (NOT
      (fsm_output(3))) AND (NOT (fsm_output(9))))) OR not_tmp_260;
  mux_2204_nl <= MUX_s_1_2_2(nand_269_nl, or_2269_nl, fsm_output(0));
  nor_787_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"))
      OR mux_2204_nl);
  nor_788_nl <= NOT((NOT (fsm_output(8))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1))
      OR (fsm_output(10)));
  nor_789_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_7(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(1)) OR (NOT (fsm_output(10))));
  mux_2203_nl <= MUX_s_1_2_2(nor_788_nl, nor_789_nl, fsm_output(7));
  mux_2205_nl <= MUX_s_1_2_2(nor_787_nl, mux_2203_nl, fsm_output(6));
  mux_2208_nl <= MUX_s_1_2_2(and_590_nl, mux_2205_nl, fsm_output(5));
  and_592_nl <= (fsm_output(7)) AND (NOT (fsm_output(8))) AND (fsm_output(0)) AND
      (VEC_LOOP_j_sva_11_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3))
      AND (fsm_output(9)) AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  nand_436_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111")) AND
      (fsm_output(3)) AND (NOT (fsm_output(9))) AND (NOT (fsm_output(1))) AND (fsm_output(10)));
  nand_434_nl <= NOT((NOT (fsm_output(3))) AND CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (fsm_output(10)));
  mux_2199_nl <= MUX_s_1_2_2(nand_436_nl, nand_434_nl, fsm_output(0));
  nor_790_nl <= NOT((fsm_output(8)) OR mux_2199_nl);
  nor_791_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_11_0(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (VEC_LOOP_j_sva_11_0(1)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2200_nl <= MUX_s_1_2_2(nor_790_nl, nor_791_nl, fsm_output(7));
  mux_2201_nl <= MUX_s_1_2_2(and_592_nl, mux_2200_nl, fsm_output(6));
  nor_792_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  and_824_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(0)) AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (VEC_LOOP_j_sva_11_0(1)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (NOT (fsm_output(1))) AND (fsm_output(10));
  and_594_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(3))
      AND (NOT (fsm_output(9))) AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  mux_2196_nl <= MUX_s_1_2_2(and_594_nl, and_591_cse, fsm_output(0));
  mux_2197_nl <= MUX_s_1_2_2(and_824_nl, mux_2196_nl, fsm_output(8));
  and_593_nl <= (fsm_output(7)) AND mux_2197_nl;
  mux_2198_nl <= MUX_s_1_2_2(nor_792_nl, and_593_nl, fsm_output(6));
  mux_2202_nl <= MUX_s_1_2_2(mux_2201_nl, mux_2198_nl, fsm_output(5));
  mux_2209_nl <= MUX_s_1_2_2(mux_2208_nl, mux_2202_nl, fsm_output(2));
  nand_274_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111")) AND
      (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(1)) AND (NOT (fsm_output(10))));
  nand_275_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111")) AND
      (NOT (fsm_output(3))) AND (fsm_output(9)) AND (fsm_output(1)) AND (NOT (fsm_output(10))));
  mux_2192_nl <= MUX_s_1_2_2(nand_274_nl, nand_275_nl, fsm_output(0));
  or_2248_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (NOT (fsm_output(3))) AND (NOT
      (fsm_output(9))))) OR not_tmp_260;
  nand_277_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND (VEC_LOOP_j_sva_11_0(2)) AND
      (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (VEC_LOOP_j_sva_11_0(1))
      AND (fsm_output(3)) AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (NOT
      (fsm_output(10))));
  mux_2191_nl <= MUX_s_1_2_2(or_2248_nl, nand_277_nl, fsm_output(0));
  mux_2193_nl <= MUX_s_1_2_2(mux_2192_nl, mux_2191_nl, fsm_output(8));
  nor_794_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))
      OR mux_2193_nl);
  nor_795_nl <= NOT((fsm_output(8)) OR (NOT (VEC_LOOP_j_sva_11_0(3))) OR (NOT (fsm_output(0)))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_11_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR
      (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(10)));
  or_2241_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(10)));
  mux_2188_nl <= MUX_s_1_2_2(nand_278_cse, or_2241_nl, fsm_output(0));
  nor_796_nl <= NOT((fsm_output(8)) OR mux_2188_nl);
  mux_2189_nl <= MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output(7));
  nor_797_nl <= NOT((NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(8)) AND (fsm_output(0)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))))
      OR not_tmp_260);
  and_596_nl <= (NOT (fsm_output(8))) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_11_0(0))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  mux_2187_nl <= MUX_s_1_2_2(nor_797_nl, and_596_nl, fsm_output(7));
  mux_2190_nl <= MUX_s_1_2_2(mux_2189_nl, mux_2187_nl, fsm_output(6));
  mux_2194_nl <= MUX_s_1_2_2(nor_794_nl, mux_2190_nl, fsm_output(5));
  nand_409_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(0))) AND (fsm_output(3))
      AND (fsm_output(9)) AND (NOT (fsm_output(1))) AND (fsm_output(10)));
  or_2233_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(3))
      OR (fsm_output(9)) OR not_tmp_260;
  mux_2183_nl <= MUX_s_1_2_2(or_2233_nl, nand_278_cse, fsm_output(0));
  mux_2184_nl <= MUX_s_1_2_2(nand_409_nl, mux_2183_nl, fsm_output(8));
  or_2230_nl <= (fsm_output(8)) OR (fsm_output(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(3)) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(10));
  mux_2185_nl <= MUX_s_1_2_2(mux_2184_nl, or_2230_nl, fsm_output(7));
  nor_798_nl <= NOT((fsm_output(6)) OR mux_2185_nl);
  and_598_nl <= (fsm_output(0)) AND CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(9))) AND (fsm_output(1)) AND (NOT
      (fsm_output(10)));
  and_599_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(1)) AND (NOT (fsm_output(10)));
  nor_799_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (VEC_LOOP_j_sva_11_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (NOT
      (fsm_output(3))) AND (NOT (fsm_output(9))))) OR not_tmp_260);
  mux_2180_nl <= MUX_s_1_2_2(and_599_nl, nor_799_nl, fsm_output(0));
  mux_2181_nl <= MUX_s_1_2_2(and_598_nl, mux_2180_nl, fsm_output(8));
  and_597_nl <= (fsm_output(7)) AND mux_2181_nl;
  nor_800_nl <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(0)) OR (fsm_output(3))
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(10)));
  mux_2182_nl <= MUX_s_1_2_2(and_597_nl, nor_800_nl, fsm_output(6));
  mux_2186_nl <= MUX_s_1_2_2(nor_798_nl, mux_2182_nl, fsm_output(5));
  mux_2195_nl <= MUX_s_1_2_2(mux_2194_nl, mux_2186_nl, fsm_output(2));
  vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_2209_nl, mux_2195_nl,
      fsm_output(4));
  and_dcpl_348 <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_350 <= and_dcpl_348 AND (NOT (fsm_output(1))) AND and_dcpl_107;
  and_dcpl_351 <= NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_353 <= (fsm_output(4)) AND (NOT (fsm_output(10)));
  and_dcpl_354 <= and_dcpl_353 AND (NOT (fsm_output(9)));
  and_dcpl_356 <= and_dcpl_354 AND and_dcpl_351 AND (fsm_output(5)) AND and_dcpl_350;
  and_dcpl_358 <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_359 <= and_dcpl_358 AND (fsm_output(1));
  and_dcpl_361 <= and_dcpl_351 AND (NOT (fsm_output(5)));
  and_850_cse <= and_dcpl_354 AND and_dcpl_361 AND and_dcpl_359 AND and_dcpl_121;
  and_dcpl_365 <= and_459_cse AND (fsm_output(1));
  and_dcpl_368 <= (NOT (fsm_output(8))) AND (fsm_output(7)) AND (fsm_output(5));
  and_857_cse <= and_dcpl_354 AND and_dcpl_368 AND and_dcpl_365 AND and_dcpl_107;
  and_dcpl_373 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_374 <= and_dcpl_373 AND (NOT (fsm_output(5)));
  and_dcpl_375 <= NOT((fsm_output(4)) OR (fsm_output(10)));
  and_dcpl_376 <= and_dcpl_375 AND (NOT (fsm_output(9)));
  and_dcpl_378 <= and_dcpl_376 AND and_dcpl_374 AND and_dcpl_358 AND (NOT (fsm_output(1)))
      AND and_dcpl_107;
  and_dcpl_380 <= and_dcpl_373 AND (fsm_output(5));
  and_869_cse <= and_dcpl_376 AND and_dcpl_380 AND and_dcpl_365 AND and_dcpl_121;
  and_dcpl_384 <= and_dcpl_348 AND (fsm_output(1));
  and_dcpl_386 <= and_dcpl_353 AND (fsm_output(9));
  and_875_cse <= and_dcpl_386 AND and_dcpl_361 AND and_dcpl_384 AND nor_tmp_217;
  and_dcpl_391 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_392 <= and_dcpl_391 AND (NOT (fsm_output(5)));
  and_dcpl_394 <= and_dcpl_386 AND and_dcpl_392 AND and_459_cse AND (NOT (fsm_output(1)))
      AND and_dcpl_107;
  and_dcpl_397 <= and_dcpl_375 AND (fsm_output(9));
  and_886_cse <= and_dcpl_397 AND and_dcpl_374 AND and_dcpl_384 AND and_dcpl_99;
  and_dcpl_401 <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("011"));
  and_dcpl_404 <= and_dcpl_397 AND and_dcpl_380 AND and_dcpl_401 AND nor_tmp_217;
  and_dcpl_406 <= (fsm_output(4)) AND (fsm_output(10)) AND (NOT (fsm_output(9)));
  and_dcpl_408 <= and_dcpl_406 AND and_dcpl_368 AND and_dcpl_350;
  and_dcpl_411 <= and_dcpl_406 AND and_dcpl_392 AND and_dcpl_401 AND and_dcpl_99;
  and_dcpl_415 <= and_dcpl_406 AND and_dcpl_391 AND (fsm_output(5)) AND and_dcpl_359
      AND nor_tmp_217;
  and_dcpl_430 <= (fsm_output(8)) AND (NOT (fsm_output(7))) AND (NOT (fsm_output(5)));
  and_dcpl_433 <= and_dcpl_353 AND (fsm_output(9)) AND and_dcpl_430 AND CONV_SL_1_1(fsm_output(3
      DOWNTO 1)=STD_LOGIC_VECTOR'("110")) AND and_dcpl_107;
  and_dcpl_441 <= (fsm_output(10)) AND (fsm_output(4)) AND (NOT (fsm_output(9)))
      AND and_dcpl_430 AND (NOT (fsm_output(3))) AND (fsm_output(2)) AND (fsm_output(1))
      AND (NOT (fsm_output(6))) AND (NOT (fsm_output(0)));
  and_dcpl_480 <= CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("010"));
  and_dcpl_502 <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(5)));
  and_dcpl_503 <= (fsm_output(10)) AND (NOT (fsm_output(4)));
  and_dcpl_511 <= and_dcpl_503 AND (fsm_output(9)) AND and_dcpl_502 AND and_dcpl_480
      AND (fsm_output(6)) AND (fsm_output(0));
  and_dcpl_517 <= (fsm_output(8)) AND (fsm_output(7)) AND (fsm_output(5));
  and_dcpl_555 <= (NOT (fsm_output(10))) AND (fsm_output(4)) AND (NOT (fsm_output(9)))
      AND and_dcpl_351 AND (fsm_output(5)) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(2)))
      AND (NOT (fsm_output(1))) AND (NOT (fsm_output(6))) AND (fsm_output(0));
  not_tmp_930 <= NOT((fsm_output(6)) AND (fsm_output(2)) AND (fsm_output(7)));
  nand_450_nl <= NOT((fsm_output(9)) AND (fsm_output(3)) AND (fsm_output(6)) AND
      (fsm_output(2)) AND (fsm_output(7)));
  or_3357_nl <= (NOT (fsm_output(9))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(2))
      OR (fsm_output(7));
  mux_tmp <= MUX_s_1_2_2(nand_450_nl, or_3357_nl, fsm_output(1));
  not_tmp_933 <= NOT((fsm_output(2)) AND (fsm_output(7)));
  nand_439_nl <= NOT((fsm_output(0)) AND (NOT mux_tmp));
  or_3373_nl <= (fsm_output(0)) OR (NOT (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(3))
      OR not_tmp_930;
  mux_3721_nl <= MUX_s_1_2_2(nand_439_nl, or_3373_nl, fsm_output(10));
  or_3371_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(3))
      OR not_tmp_930;
  or_3369_nl <= (fsm_output(0)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR (fsm_output(7));
  mux_3720_nl <= MUX_s_1_2_2(or_3371_nl, or_3369_nl, fsm_output(10));
  mux_3722_nl <= MUX_s_1_2_2(mux_3721_nl, mux_3720_nl, fsm_output(4));
  or_3367_nl <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR (fsm_output(7));
  or_3366_nl <= (NOT (fsm_output(1))) OR (fsm_output(9)) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (fsm_output(7));
  mux_3718_nl <= MUX_s_1_2_2(or_3367_nl, or_3366_nl, fsm_output(0));
  or_3365_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(3))
      OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR (fsm_output(7));
  mux_3719_nl <= MUX_s_1_2_2(mux_3718_nl, or_3365_nl, fsm_output(10));
  or_3368_nl <= (fsm_output(4)) OR mux_3719_nl;
  mux_3723_nl <= MUX_s_1_2_2(mux_3722_nl, or_3368_nl, fsm_output(5));
  nor_1381_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(9)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR not_tmp_933);
  nor_1382_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (fsm_output(3))
      OR (fsm_output(6)) OR not_tmp_933);
  mux_3715_nl <= MUX_s_1_2_2(nor_1381_nl, nor_1382_nl, fsm_output(0));
  nor_1383_nl <= NOT((fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(3))
      OR (fsm_output(6)) OR (fsm_output(2)) OR (NOT (fsm_output(7))));
  mux_3716_nl <= MUX_s_1_2_2(mux_3715_nl, nor_1383_nl, fsm_output(10));
  nand_445_nl <= NOT((fsm_output(4)) AND mux_3716_nl);
  or_3358_nl <= (NOT (fsm_output(10))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(1)))
      OR (fsm_output(9)) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(2))
      OR (fsm_output(7));
  or_3356_nl <= (fsm_output(1)) OR (fsm_output(9)) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(2)) OR (fsm_output(7));
  mux_3712_nl <= MUX_s_1_2_2(mux_tmp, or_3356_nl, fsm_output(0));
  or_3355_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(3))
      OR not_tmp_930;
  mux_3713_nl <= MUX_s_1_2_2(mux_3712_nl, or_3355_nl, fsm_output(10));
  mux_3714_nl <= MUX_s_1_2_2(or_3358_nl, mux_3713_nl, fsm_output(4));
  mux_3717_nl <= MUX_s_1_2_2(nand_445_nl, mux_3714_nl, fsm_output(5));
  mux_3724_itm <= MUX_s_1_2_2(mux_3723_nl, mux_3717_nl, fsm_output(8));
  and_dcpl_564 <= NOT((fsm_output(10)) OR (fsm_output(4)) OR (fsm_output(9)) OR (NOT
      and_dcpl_351) OR (fsm_output(5)) OR (NOT (fsm_output(3))) OR (fsm_output(2))
      OR (NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(0)));
  and_dcpl_568 <= and_dcpl_348 AND (NOT (fsm_output(1))) AND (NOT (fsm_output(6)))
      AND (fsm_output(0));
  and_dcpl_574 <= (fsm_output(4)) AND (NOT (fsm_output(10))) AND (NOT (fsm_output(9)))
      AND and_dcpl_351 AND (fsm_output(5)) AND and_dcpl_568;
  or_tmp_3188 <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("01000"));
  or_tmp_3189 <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("01001"));
  mux_tmp_3724 <= MUX_s_1_2_2(or_tmp_3189, or_tmp_3188, fsm_output(2));
  or_tmp_3191 <= (fsm_output(6)) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  or_tmp_3193 <= (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_tmp_3725 <= MUX_s_1_2_2(or_tmp_3193, or_tmp_3191, fsm_output(7));
  or_tmp_3195 <= (NOT (fsm_output(6))) OR (fsm_output(9)) OR not_tmp_51;
  or_tmp_3196 <= (NOT (fsm_output(6))) OR (fsm_output(9)) OR (NOT (fsm_output(8)))
      OR (fsm_output(10));
  mux_tmp_3728 <= MUX_s_1_2_2(or_tmp_3196, or_tmp_3195, fsm_output(7));
  or_tmp_3200 <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("10000"));
  or_tmp_3202 <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("10001"));
  or_tmp_3203 <= (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(10));
  mux_tmp_3733 <= MUX_s_1_2_2(or_tmp_3195, or_tmp_3203, fsm_output(7));
  or_tmp_3204 <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("01101"));
  or_tmp_3205 <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("01110"));
  mux_tmp_3735 <= MUX_s_1_2_2(or_tmp_3205, or_tmp_3204, fsm_output(2));
  nand_455_nl <= NOT((fsm_output(6)) AND (fsm_output(9)) AND (NOT (fsm_output(8)))
      AND (fsm_output(10)));
  mux_tmp_3737 <= MUX_s_1_2_2(nand_455_nl, or_tmp_3196, fsm_output(7));
  or_tmp_3211 <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("01011"));
  or_3396_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("01010"));
  mux_tmp_3742 <= MUX_s_1_2_2(or_tmp_3211, or_3396_nl, fsm_output(2));
  or_tmp_3212 <= (fsm_output(6)) OR (fsm_output(9)) OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_tmp_3743 <= MUX_s_1_2_2(or_tmp_3212, or_tmp_3193, fsm_output(7));
  or_tmp_3213 <= NOT(CONV_SL_1_1(fsm_output(10 DOWNTO 6)=STD_LOGIC_VECTOR'("01111")));
  or_tmp_3218 <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("01100"));
  mux_tmp_3751 <= MUX_s_1_2_2(or_tmp_3200, or_tmp_3213, fsm_output(2));
  or_3406_nl <= (NOT (fsm_output(6))) OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT
      (fsm_output(10)));
  mux_tmp_3753 <= MUX_s_1_2_2(or_tmp_3203, or_3406_nl, fsm_output(7));
  or_3409_nl <= (fsm_output(6)) OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_tmp_3762 <= MUX_s_1_2_2(or_tmp_3191, or_3409_nl, fsm_output(7));
  or_3413_nl <= (fsm_output(6)) OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (NOT
      (fsm_output(10)));
  mux_3771_nl <= MUX_s_1_2_2(or_3413_nl, or_tmp_3212, fsm_output(7));
  mux_tmp_3771 <= MUX_s_1_2_2(mux_3771_nl, mux_tmp_3728, fsm_output(2));
  or_3420_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("11010"));
  mux_3783_nl <= MUX_s_1_2_2(or_3420_nl, mux_tmp_3737, fsm_output(2));
  or_3418_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("00011"));
  mux_3782_nl <= MUX_s_1_2_2(mux_tmp_3743, or_3418_nl, fsm_output(2));
  mux_3784_nl <= MUX_s_1_2_2(mux_3783_nl, mux_3782_nl, fsm_output(4));
  mux_3780_nl <= MUX_s_1_2_2(mux_tmp_3762, or_tmp_3202, fsm_output(2));
  mux_3781_nl <= MUX_s_1_2_2(mux_tmp_3742, mux_3780_nl, fsm_output(4));
  mux_3785_nl <= MUX_s_1_2_2(mux_3784_nl, mux_3781_nl, fsm_output(5));
  or_3417_nl <= (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR not_tmp_51;
  mux_3777_nl <= MUX_s_1_2_2(or_3417_nl, mux_tmp_3725, fsm_output(2));
  mux_3778_nl <= MUX_s_1_2_2(mux_tmp_3735, mux_3777_nl, fsm_output(4));
  or_3415_nl <= (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  mux_3776_nl <= MUX_s_1_2_2(or_3415_nl, mux_tmp_3771, fsm_output(4));
  mux_3779_nl <= MUX_s_1_2_2(mux_3778_nl, mux_3776_nl, fsm_output(5));
  mux_3786_nl <= MUX_s_1_2_2(mux_3785_nl, mux_3779_nl, fsm_output(0));
  mux_3770_nl <= MUX_s_1_2_2(or_tmp_3204, or_tmp_3218, fsm_output(2));
  mux_3773_nl <= MUX_s_1_2_2(mux_tmp_3771, mux_3770_nl, fsm_output(4));
  or_3411_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("10011"));
  mux_3768_nl <= MUX_s_1_2_2(or_tmp_3189, or_3411_nl, fsm_output(2));
  mux_3769_nl <= MUX_s_1_2_2(mux_3768_nl, mux_tmp_3751, fsm_output(4));
  mux_3774_nl <= MUX_s_1_2_2(mux_3773_nl, mux_3769_nl, fsm_output(5));
  mux_3765_nl <= MUX_s_1_2_2(or_tmp_3218, or_tmp_3211, fsm_output(2));
  mux_3764_nl <= MUX_s_1_2_2(mux_tmp_3753, mux_tmp_3762, fsm_output(2));
  mux_3766_nl <= MUX_s_1_2_2(mux_3765_nl, mux_3764_nl, fsm_output(4));
  mux_3761_nl <= MUX_s_1_2_2(or_tmp_3188, mux_tmp_3737, fsm_output(2));
  or_3407_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("00100"));
  mux_3760_nl <= MUX_s_1_2_2(or_3407_nl, or_tmp_3205, fsm_output(2));
  mux_3762_nl <= MUX_s_1_2_2(mux_3761_nl, mux_3760_nl, fsm_output(4));
  mux_3767_nl <= MUX_s_1_2_2(mux_3766_nl, mux_3762_nl, fsm_output(5));
  mux_3775_nl <= MUX_s_1_2_2(mux_3774_nl, mux_3767_nl, fsm_output(0));
  mux_3787_nl <= MUX_s_1_2_2(mux_3786_nl, mux_3775_nl, fsm_output(3));
  mux_3755_nl <= MUX_s_1_2_2(mux_tmp_3725, mux_tmp_3753, fsm_output(2));
  mux_3756_nl <= MUX_s_1_2_2(mux_3755_nl, mux_tmp_3724, fsm_output(4));
  or_3403_nl <= (NOT (fsm_output(7))) OR (fsm_output(6)) OR (fsm_output(9)) OR not_tmp_51;
  mux_3751_nl <= MUX_s_1_2_2(or_tmp_3218, or_3403_nl, fsm_output(2));
  mux_3753_nl <= MUX_s_1_2_2(mux_tmp_3751, mux_3751_nl, fsm_output(4));
  mux_3757_nl <= MUX_s_1_2_2(mux_3756_nl, mux_3753_nl, fsm_output(5));
  or_3401_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("10010"));
  mux_3748_nl <= MUX_s_1_2_2(or_tmp_3188, or_3401_nl, fsm_output(2));
  mux_3747_nl <= MUX_s_1_2_2(or_tmp_3213, or_tmp_3205, fsm_output(2));
  mux_3749_nl <= MUX_s_1_2_2(mux_3748_nl, mux_3747_nl, fsm_output(4));
  mux_3745_nl <= MUX_s_1_2_2(mux_tmp_3743, mux_tmp_3733, fsm_output(2));
  mux_3746_nl <= MUX_s_1_2_2(mux_3745_nl, mux_tmp_3742, fsm_output(4));
  mux_3750_nl <= MUX_s_1_2_2(mux_3749_nl, mux_3746_nl, fsm_output(5));
  mux_3758_nl <= MUX_s_1_2_2(mux_3757_nl, mux_3750_nl, fsm_output(0));
  or_3395_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(6))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_3392_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("00110"));
  mux_3739_nl <= MUX_s_1_2_2(mux_tmp_3737, or_3392_nl, fsm_output(2));
  mux_3740_nl <= MUX_s_1_2_2(or_3395_nl, mux_3739_nl, fsm_output(4));
  mux_3735_nl <= MUX_s_1_2_2(mux_tmp_3733, mux_tmp_3725, fsm_output(2));
  mux_3737_nl <= MUX_s_1_2_2(mux_tmp_3735, mux_3735_nl, fsm_output(4));
  mux_3741_nl <= MUX_s_1_2_2(mux_3740_nl, mux_3737_nl, fsm_output(5));
  mux_3731_nl <= MUX_s_1_2_2(or_tmp_3202, or_tmp_3200, fsm_output(2));
  or_3384_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("11000"));
  mux_3730_nl <= MUX_s_1_2_2(or_3384_nl, mux_tmp_3728, fsm_output(2));
  mux_3732_nl <= MUX_s_1_2_2(mux_3731_nl, mux_3730_nl, fsm_output(4));
  or_3376_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 6)/=STD_LOGIC_VECTOR'("00001"));
  mux_3727_nl <= MUX_s_1_2_2(mux_tmp_3725, or_3376_nl, fsm_output(2));
  mux_3728_nl <= MUX_s_1_2_2(mux_3727_nl, mux_tmp_3724, fsm_output(4));
  mux_3733_nl <= MUX_s_1_2_2(mux_3732_nl, mux_3728_nl, fsm_output(5));
  mux_3742_nl <= MUX_s_1_2_2(mux_3741_nl, mux_3733_nl, fsm_output(0));
  mux_3759_nl <= MUX_s_1_2_2(mux_3758_nl, mux_3742_nl, fsm_output(3));
  mux_3788_itm <= MUX_s_1_2_2(mux_3787_nl, mux_3759_nl, fsm_output(1));
  and_dcpl_579 <= (NOT (fsm_output(4))) AND (NOT (fsm_output(10))) AND (NOT (fsm_output(9)))
      AND and_dcpl_351 AND (NOT (fsm_output(5))) AND and_dcpl_568;
  and_dcpl_588 <= (NOT (fsm_output(4))) AND (fsm_output(10)) AND (fsm_output(9))
      AND (NOT (fsm_output(8))) AND (fsm_output(7)) AND (NOT (fsm_output(5))) AND
      and_dcpl_348 AND (fsm_output(1)) AND (NOT (fsm_output(6))) AND (NOT (fsm_output(0)));
  and_dcpl_591 <= and_dcpl_348 AND (NOT (fsm_output(1)));
  and_dcpl_592 <= and_dcpl_591 AND and_dcpl_107;
  and_dcpl_598 <= and_dcpl_354 AND and_dcpl_351 AND (fsm_output(5)) AND and_dcpl_592;
  and_dcpl_614 <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_615 <= and_dcpl_614 AND (NOT (fsm_output(1)));
  and_dcpl_618 <= and_dcpl_391 AND (fsm_output(5));
  and_dcpl_622 <= and_dcpl_376 AND and_dcpl_618 AND and_dcpl_615 AND and_dcpl_99;
  and_dcpl_623 <= and_dcpl_358 AND (NOT (fsm_output(1)));
  and_dcpl_624 <= and_dcpl_623 AND and_dcpl_107;
  and_dcpl_628 <= and_dcpl_376 AND and_dcpl_374 AND and_dcpl_624;
  and_dcpl_641 <= and_dcpl_386 AND and_dcpl_368 AND and_dcpl_623 AND and_dcpl_99;
  and_dcpl_642 <= and_459_cse AND (NOT (fsm_output(1)));
  and_dcpl_646 <= and_dcpl_386 AND and_dcpl_392 AND and_dcpl_642 AND and_dcpl_107;
  and_dcpl_651 <= and_dcpl_614 AND (fsm_output(1));
  and_dcpl_654 <= and_dcpl_397 AND and_dcpl_380 AND and_dcpl_651 AND nor_tmp_217;
  and_dcpl_657 <= and_dcpl_503 AND (NOT (fsm_output(9)));
  and_dcpl_659 <= and_dcpl_657 AND and_dcpl_361 AND and_dcpl_642 AND and_dcpl_121;
  and_dcpl_663 <= and_dcpl_406 AND and_dcpl_368 AND and_dcpl_592;
  and_dcpl_666 <= and_dcpl_406 AND and_dcpl_392 AND and_dcpl_651 AND and_dcpl_99;
  and_dcpl_669 <= and_dcpl_406 AND and_dcpl_618 AND and_dcpl_359 AND nor_tmp_217;
  and_dcpl_672 <= and_dcpl_657 AND and_dcpl_380 AND and_dcpl_591 AND and_dcpl_121;
  and_dcpl_676 <= and_dcpl_503 AND (fsm_output(9)) AND and_dcpl_361 AND and_dcpl_615
      AND nor_tmp_217;
  and_dcpl_678 <= and_dcpl_376 AND and_dcpl_361 AND and_dcpl_624;
  and_dcpl_688 <= NOT(CONV_SL_1_1(fsm_output/=STD_LOGIC_VECTOR'("00100100100")));
  and_dcpl_698 <= (NOT (fsm_output(4))) AND (fsm_output(10)) AND (NOT (fsm_output(9)))
      AND and_dcpl_351 AND (NOT (fsm_output(5))) AND (fsm_output(3)) AND (fsm_output(2))
      AND (NOT (fsm_output(1))) AND (fsm_output(6)) AND (NOT (fsm_output(0)));
  nor_1369_nl <= NOT((fsm_output(10)) OR (NOT((fsm_output(9)) AND (fsm_output(1))
      AND (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6)))));
  nor_1370_nl <= NOT((fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(3)) OR nand_257_cse);
  nor_1371_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(8)) OR (fsm_output(6)));
  mux_3799_nl <= MUX_s_1_2_2(nor_1370_nl, nor_1371_nl, fsm_output(9));
  and_1249_nl <= (fsm_output(10)) AND mux_3799_nl;
  mux_3800_nl <= MUX_s_1_2_2(nor_1369_nl, and_1249_nl, fsm_output(2));
  and_1248_nl <= (fsm_output(4)) AND mux_3800_nl;
  or_3441_nl <= (fsm_output(10)) OR (fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(0))
      OR (fsm_output(3)) OR nand_257_cse;
  or_3439_nl <= (NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(0)) OR (NOT
      (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(6));
  or_3438_nl <= (fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (fsm_output(8)) OR (fsm_output(6));
  mux_3797_nl <= MUX_s_1_2_2(or_3439_nl, or_3438_nl, fsm_output(10));
  mux_3798_nl <= MUX_s_1_2_2(or_3441_nl, mux_3797_nl, fsm_output(2));
  nor_1372_nl <= NOT((fsm_output(4)) OR mux_3798_nl);
  mux_3801_nl <= MUX_s_1_2_2(and_1248_nl, nor_1372_nl, fsm_output(5));
  nor_1373_nl <= NOT((NOT (fsm_output(9))) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(3)) OR nand_257_cse);
  nor_1374_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(1))) OR (fsm_output(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(6)));
  mux_3793_nl <= MUX_s_1_2_2(nor_1373_nl, nor_1374_nl, fsm_output(10));
  nor_1375_nl <= NOT((fsm_output(10)) OR (fsm_output(9)) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR nand_257_cse);
  mux_3794_nl <= MUX_s_1_2_2(mux_3793_nl, nor_1375_nl, fsm_output(2));
  or_3431_nl <= (fsm_output(1)) OR (fsm_output(0)) OR (NOT (fsm_output(3))) OR (fsm_output(8))
      OR (fsm_output(6));
  or_3430_nl <= (fsm_output(1)) OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(8))
      OR (fsm_output(6));
  mux_3792_nl <= MUX_s_1_2_2(or_3431_nl, or_3430_nl, fsm_output(9));
  nor_1376_nl <= NOT((fsm_output(2)) OR (fsm_output(10)) OR mux_3792_nl);
  mux_3795_nl <= MUX_s_1_2_2(mux_3794_nl, nor_1376_nl, fsm_output(4));
  and_1250_nl <= (fsm_output(2)) AND (fsm_output(10)) AND (NOT (fsm_output(9))) AND
      (fsm_output(1)) AND (fsm_output(0)) AND (fsm_output(3)) AND (NOT (fsm_output(8)))
      AND (fsm_output(6));
  nor_1378_nl <= NOT((NOT (fsm_output(10))) OR (fsm_output(9)) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(8)))
      OR (fsm_output(6)));
  or_3424_nl <= (fsm_output(1)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(8)) OR (NOT (fsm_output(6)));
  or_3422_nl <= (NOT (fsm_output(1))) OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(8))
      OR (NOT (fsm_output(6)));
  mux_3789_nl <= MUX_s_1_2_2(or_3424_nl, or_3422_nl, fsm_output(9));
  nor_1379_nl <= NOT((fsm_output(10)) OR mux_3789_nl);
  mux_3790_nl <= MUX_s_1_2_2(nor_1378_nl, nor_1379_nl, fsm_output(2));
  mux_3791_nl <= MUX_s_1_2_2(and_1250_nl, mux_3790_nl, fsm_output(4));
  mux_3796_nl <= MUX_s_1_2_2(mux_3795_nl, mux_3791_nl, fsm_output(5));
  not_tmp_980 <= MUX_s_1_2_2(mux_3801_nl, mux_3796_nl, fsm_output(7));
  and_dcpl_707 <= (fsm_output(4)) AND (NOT (fsm_output(10))) AND (NOT (fsm_output(9)))
      AND and_dcpl_351 AND (fsm_output(5)) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(2)))
      AND (fsm_output(1)) AND (NOT (fsm_output(6))) AND (fsm_output(0));
  and_dcpl_717 <= and_dcpl_353 AND (fsm_output(9)) AND (NOT (fsm_output(8))) AND
      (fsm_output(7)) AND (fsm_output(5)) AND and_dcpl_358 AND (NOT (fsm_output(1)))
      AND and_dcpl_99;
  and_dcpl_727 <= (fsm_output(10)) AND (NOT (fsm_output(4))) AND (NOT (fsm_output(9)))
      AND and_dcpl_373 AND (fsm_output(5)) AND and_dcpl_348 AND (NOT (fsm_output(1)))
      AND and_dcpl_121;
  and_dcpl_734 <= and_dcpl_353 AND (NOT (fsm_output(9))) AND (NOT (fsm_output(8)))
      AND (NOT (fsm_output(7))) AND (NOT (fsm_output(5))) AND and_dcpl_358 AND (fsm_output(1))
      AND and_dcpl_121;
  and_dcpl_741 <= (NOT (fsm_output(10))) AND (NOT (fsm_output(4))) AND (fsm_output(9))
      AND and_dcpl_373 AND (NOT (fsm_output(5))) AND and_dcpl_348 AND (fsm_output(1))
      AND and_dcpl_99;
  COMP_LOOP_or_55_ssc <= and_857_cse OR and_dcpl_628 OR and_875_cse OR and_dcpl_672;
  COMP_LOOP_or_56_ssc <= and_dcpl_622 OR and_dcpl_641 OR and_dcpl_659 OR and_dcpl_676;
  COMP_LOOP_or_57_ssc <= and_869_cse OR and_dcpl_654 OR and_dcpl_663 OR and_dcpl_669;
  COMP_LOOP_or_58_ssc <= and_dcpl_646 OR and_dcpl_666;
  or_tmp <= (fsm_output(9)) OR (NOT (fsm_output(4)));
  nor_tmp <= (fsm_output(2)) AND (fsm_output(4));
  mux_tmp_3818 <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), fsm_output(2));
  not_tmp_1007 <= NOT((fsm_output(2)) OR (fsm_output(4)));
  mux_tmp_3819 <= MUX_s_1_2_2(not_tmp_1007, mux_tmp_3818, fsm_output(0));
  mux_tmp_3822 <= MUX_s_1_2_2(mux_tmp_3818, nor_tmp, or_2348_cse);
  or_tmp_3291 <= and_563_cse OR (fsm_output(4));
  or_tmp_3293 <= (fsm_output(9)) OR (NOT or_tmp_3291);
  nor_tmp_535 <= ((fsm_output(9)) OR (fsm_output(2))) AND (fsm_output(4));
  nor_tmp_536 <= or_2348_cse AND (fsm_output(2)) AND (fsm_output(4));
  mux_tmp_3828 <= MUX_s_1_2_2((NOT or_tmp_3291), nor_tmp_536, fsm_output(9));
  mux_tmp_3834 <= MUX_s_1_2_2(mux_tmp_3822, (fsm_output(4)), fsm_output(9));
  nor_tmp_539 <= or_3280_cse AND (fsm_output(4));
  nor_tmp_540 <= or_2385_cse AND (fsm_output(4));
  or_tmp_3303 <= and_573_cse OR (fsm_output(2)) OR (fsm_output(4));
  or_tmp_3304 <= ((fsm_output(9)) AND (fsm_output(2))) OR (fsm_output(4));
  mux_tmp_3846 <= MUX_s_1_2_2(mux_tmp_3818, nor_tmp, fsm_output(0));
  mux_tmp_3853 <= MUX_s_1_2_2((NOT or_tmp_3291), nor_tmp_540, fsm_output(9));
  not_tmp_1021 <= NOT(((fsm_output(9)) AND (fsm_output(1)) AND (fsm_output(0)) AND
      (fsm_output(2))) OR (fsm_output(4)));
  nor_1460_nl <= NOT((fsm_output(0)) OR (fsm_output(2)) OR (fsm_output(4)));
  and_1267_nl <= (fsm_output(0)) AND (fsm_output(2)) AND (fsm_output(4));
  mux_tmp_3861 <= MUX_s_1_2_2(nor_1460_nl, and_1267_nl, fsm_output(1));
  mux_tmp_3878 <= MUX_s_1_2_2(mux_tmp_3819, mux_tmp_3846, fsm_output(1));
  or_tmp_3320 <= (fsm_output(1)) OR (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(8)))
      OR (fsm_output(10)) OR (fsm_output(9)) OR (fsm_output(4));
  not_tmp_1034 <= NOT((fsm_output(9)) AND (fsm_output(4)));
  or_tmp_3327 <= (fsm_output(10)) OR not_tmp_1034;
  mux_3898_nl <= MUX_s_1_2_2(or_tmp_3327, or_tmp_2652, fsm_output(8));
  or_3516_nl <= (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8)) OR (fsm_output(10))
      OR not_tmp_1034;
  mux_tmp_3898 <= MUX_s_1_2_2(mux_3898_nl, or_3516_nl, fsm_output(1));
  or_tmp_3332 <= (fsm_output(8)) OR (fsm_output(10)) OR (NOT (fsm_output(9))) OR
      (fsm_output(4));
  nand_470_nl <= NOT(COMP_LOOP_nor_11_itm AND (fsm_output(8)) AND (fsm_output(10))
      AND (NOT (fsm_output(9))) AND (fsm_output(4)));
  mux_3902_nl <= MUX_s_1_2_2(or_tmp_3332, nand_470_nl, fsm_output(1));
  nand_tmp <= NOT((fsm_output(6)) AND (NOT mux_3902_nl));
  mux_tmp_3902 <= MUX_s_1_2_2(or_tmp_195, or_tmp_3327, fsm_output(8));
  or_3531_nl <= (fsm_output(8)) OR (NOT (fsm_output(10))) OR (fsm_output(9)) OR (fsm_output(4));
  mux_3906_nl <= MUX_s_1_2_2(or_tmp, or_2747_cse, fsm_output(10));
  or_3530_nl <= (fsm_output(8)) OR mux_3906_nl;
  mux_tmp_3906 <= MUX_s_1_2_2(or_3531_nl, or_3530_nl, COMP_LOOP_nor_11_itm);
  or_tmp_3343 <= (NOT (fsm_output(1))) OR (fsm_output(8)) OR (fsm_output(10)) OR
      (fsm_output(9)) OR (fsm_output(4));
  mux_tmp_3915 <= MUX_s_1_2_2(or_2415_cse, or_tmp_182, fsm_output(8));
  or_tmp_3369 <= (fsm_output(8)) OR (fsm_output(10)) OR (fsm_output(9)) OR (NOT (fsm_output(4)));
  COMP_LOOP_or_60_itm <= and_850_cse OR and_857_cse OR and_dcpl_378 OR and_869_cse
      OR and_875_cse OR and_dcpl_394 OR and_886_cse OR and_dcpl_404 OR and_dcpl_408
      OR and_dcpl_411 OR and_dcpl_415;
  COMP_LOOP_or_24_itm <= and_dcpl_433 OR and_dcpl_441;
  COMP_LOOP_COMP_LOOP_or_6_cse <= (NOT and_dcpl_441) OR (and_dcpl_353 AND (NOT (fsm_output(9)))
      AND and_dcpl_351 AND (fsm_output(5)) AND nor_738_cse AND and_dcpl_107) OR and_dcpl_433;
  COMP_LOOP_or_67_itm <= and_dcpl_688 OR and_dcpl_698;
  COMP_LOOP_COMP_LOOP_or_9_cse <= (NOT(and_dcpl_688 OR and_dcpl_698)) OR not_tmp_980
      OR and_dcpl_707;
  COMP_LOOP_nor_680_itm <= NOT(not_tmp_980 OR and_dcpl_707);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_219 = '0' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((and_dcpl_103 AND and_dcpl_98) OR STAGE_LOOP_i_3_0_sva_mx0c1) = '1' )
          THEN
        STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "0001"), STAGE_LOOP_i_3_0_sva_2,
            STAGE_LOOP_i_3_0_sva_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_219 = '0' ) THEN
        r_sva <= r_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= '0';
        COMP_LOOP_nor_11_itm <= '0';
        modExp_exp_1_7_1_sva <= '0';
        COMP_LOOP_nor_12_itm <= '0';
        COMP_LOOP_nor_134_itm <= '0';
        COMP_LOOP_nor_137_itm <= '0';
        COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= '0';
        COMP_LOOP_COMP_LOOP_nor_1_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_139_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_140_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_141_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_143_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_144_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_145_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_146_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_147_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_148_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_149_itm <= '0';
      ELSE
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_111 AND and_dcpl_97 AND and_dcpl_50
            AND (NOT STAGE_LOOP_acc_itm_2_1);
        COMP_LOOP_nor_11_itm <= (COMP_LOOP_mux1h_428_nl AND (mux_2888_nl OR (fsm_output(0))))
            OR (mux_2983_nl AND (fsm_output(0)));
        modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_464_nl AND (NOT mux_3396_nl);
        COMP_LOOP_nor_12_itm <= (COMP_LOOP_mux1h_474_nl AND (NOT(mux_3417_nl AND
            (fsm_output(1))))) OR (NOT(mux_3513_nl OR (fsm_output(1))));
        COMP_LOOP_nor_134_itm <= (COMP_LOOP_mux1h_477_nl AND mux_3584_nl) OR mux_3591_nl;
        COMP_LOOP_nor_137_itm <= (COMP_LOOP_mux1h_479_nl AND (mux_3598_nl OR (fsm_output(10))))
            OR mux_3605_nl;
        COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= COMP_LOOP_mux1h_480_nl AND (NOT and_dcpl_283);
        COMP_LOOP_COMP_LOOP_nor_1_itm <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_COMP_LOOP_and_139_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_140_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_141_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_COMP_LOOP_and_143_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_144_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_145_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_146_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_147_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_148_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_149_itm <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      modulo_result_rem_cmp_a <= MUX1HOT_v_64_6_2(z_out_10, operator_64_false_acc_mut_63_0,
          COMP_LOOP_10_acc_8_itm, COMP_LOOP_1_modExp_1_while_if_mul_mut_1, COMP_LOOP_10_mul_mut,
          z_out_5, STD_LOGIC_VECTOR'( modulo_result_or_nl & (NOT mux_2303_nl) & (NOT
          mux_2378_nl) & mux_2394_nl & (NOT mux_2461_nl) & (NOT mux_2475_itm)));
      modulo_result_rem_cmp_b <= p_sva;
      operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_6, (operator_64_false_acc_mut_64
          & operator_64_false_acc_mut_63_0), and_dcpl_266);
      operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
          STAGE_LOOP_lshift_psp_sva, and_dcpl_266);
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_2495_nl = '0' ) THEN
        STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_3896_nl = '0' ) THEN
        operator_64_false_acc_mut_64 <= operator_64_false_mux1h_2_rgt(64);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_3949_nl = '0' ) THEN
        operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_2_rgt(63 DOWNTO
            0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_j_sva_11_0 <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (and_dcpl_273 OR VEC_LOOP_j_sva_11_0_mx0c1) = '1' ) THEN
        VEC_LOOP_j_sva_11_0 <= MUX_v_12_2_2(STD_LOGIC_VECTOR'("000000000000"), (z_out_6(11
            DOWNTO 0)), VEC_LOOP_j_sva_11_0_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_k_9_4_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( (NOT(mux_3952_nl OR (fsm_output(8)))) = '1' ) THEN
        COMP_LOOP_k_9_4_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (COMP_LOOP_k_9_4_sva_2(4
            DOWNTO 0)), or_3477_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((modExp_while_and_3 OR modExp_while_and_5 OR modExp_result_sva_mx0c0
          OR (NOT mux_2675_nl)) AND (modExp_result_sva_mx0c0 OR modExp_result_and_rgt
          OR modExp_result_and_1_rgt)) = '1' ) THEN
        modExp_result_sva <= MUX1HOT_v_64_3_2(STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
            modulo_result_rem_cmp_z, (z_out_6(63 DOWNTO 0)), STD_LOGIC_VECTOR'( modExp_result_sva_mx0c0
            & modExp_result_and_rgt & modExp_result_and_1_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        tmp_10_lpi_4_dfm <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
      ELSIF ( (MUX_s_1_2_2((NOT mux_2740_nl), mux_2705_nl, fsm_output(9))) = '1'
          ) THEN
        tmp_10_lpi_4_dfm <= MUX1HOT_v_64_17_2(('0' & operator_64_false_slc_modExp_exp_63_1_3),
            vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
            vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d,
            vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d,
            vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d,
            STD_LOGIC_VECTOR'( and_dcpl_273 & COMP_LOOP_or_8_nl & COMP_LOOP_or_9_nl
            & COMP_LOOP_or_10_nl & COMP_LOOP_or_11_nl & COMP_LOOP_or_12_nl & COMP_LOOP_or_13_nl
            & COMP_LOOP_or_14_nl & COMP_LOOP_or_15_nl & COMP_LOOP_or_16_nl & COMP_LOOP_or_17_nl
            & COMP_LOOP_or_18_nl & COMP_LOOP_or_19_nl & COMP_LOOP_or_20_nl & COMP_LOOP_or_21_nl
            & COMP_LOOP_or_22_nl & COMP_LOOP_or_23_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2867_nl, mux_2822_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_10_mul_mut <= MUX1HOT_v_64_21_2(r_sva, modulo_result_rem_cmp_z,
            (z_out_6(63 DOWNTO 0)), modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
            vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d,
            vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d,
            vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d,
            vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d, COMP_LOOP_1_modExp_1_while_if_mul_mut_1,
            STD_LOGIC_VECTOR'( and_340_nl & COMP_LOOP_or_30_nl & COMP_LOOP_or_31_nl
            & not_tmp_596 & COMP_LOOP_and_277_nl & COMP_LOOP_COMP_LOOP_and_932_nl
            & COMP_LOOP_COMP_LOOP_and_934_nl & COMP_LOOP_and_1_nl & COMP_LOOP_COMP_LOOP_and_936_nl
            & COMP_LOOP_and_2_nl & COMP_LOOP_and_3_nl & COMP_LOOP_and_4_nl & COMP_LOOP_COMP_LOOP_and_930_nl
            & COMP_LOOP_and_5_nl & COMP_LOOP_and_6_nl & COMP_LOOP_and_7_nl & COMP_LOOP_and_8_nl
            & COMP_LOOP_and_9_nl & COMP_LOOP_and_10_nl & COMP_LOOP_and_11_nl & mux_114_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= '0';
      ELSIF ( (and_dcpl_260 OR and_dcpl_332 OR and_dcpl_126 OR and_dcpl_141 OR and_dcpl_147
          OR and_dcpl_158 OR and_dcpl_164 OR and_dcpl_175 OR and_dcpl_182 OR and_dcpl_192
          OR and_dcpl_198 OR and_dcpl_206 OR and_dcpl_217 OR and_dcpl_225 OR and_dcpl_232
          OR and_dcpl_242 OR and_dcpl_247 OR and_dcpl_255) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= MUX1HOT_s_1_3_2((NOT (z_out_5(63))), (NOT
            (z_out_8_8_7(1))), COMP_LOOP_COMP_LOOP_and_17_nl, STD_LOGIC_VECTOR'(
            and_dcpl_260 & and_dcpl_332 & COMP_LOOP_or_32_cse));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_3181_nl OR (NOT mux_2475_itm)) = '1' ) THEN
        COMP_LOOP_10_acc_8_itm <= MUX_v_64_2_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(COMP_LOOP_1_acc_8_nl),
            64)), z_out_10, mux_2475_itm);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(or_tmp_9 OR (NOT (fsm_output(0))) OR (fsm_output(6)) OR (fsm_output(7))
          OR (NOT (fsm_output(5))) OR (fsm_output(2)) OR (fsm_output(8)) OR (NOT
          (fsm_output(4))) OR (fsm_output(9)))) = '1' ) THEN
        COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= NOT(CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_305_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_305_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_62_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_62_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_2_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_2_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_64_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_64_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_4_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_4_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_5_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_5_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_6_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_6_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_68_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_68_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_8_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_8_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_9_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_9_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_10_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(nor_nl, and_1253_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_10_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_10_nl,
            (NOT (COMP_LOOP_1_acc_nl(9))), and_dcpl_255);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_11_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_11_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_12_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_12_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_13_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_13_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_14_itm <= '0';
      ELSIF ( not_tmp_708 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_14_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (mux_3224_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_6_sva <= COMP_LOOP_acc_1_cse_6_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_2_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (mux_3234_nl OR CONV_SL_1_1(fsm_output(10 DOWNTO 8)/=STD_LOGIC_VECTOR'("000")))
          = '1' ) THEN
        COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (NOT((NOT mux_3242_nl) AND nor_601_cse)) = '1' ) THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "001")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_4_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (NOT(mux_3243_nl AND nor_601_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_4_sva <= z_out_5(11 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_3249_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_13_psp_sva <= z_out;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (mux_3251_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "011")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_8_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (mux_3255_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_8_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "0111")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_16_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (mux_3263_nl OR (fsm_output(10))) = '1' ) THEN
        COMP_LOOP_acc_16_psp_sva <= z_out_7(8 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_10_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3267_nl, mux_3264_nl, fsm_output(4))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_10_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1001")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_17_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3276_nl, (fsm_output(10)), fsm_output(9))) = '1' )
          THEN
        COMP_LOOP_acc_17_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "101")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_12_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3288_nl, mux_3287_nl, fsm_output(4))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_12_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1011")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_19_psp_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3292_nl, (fsm_output(10)), fsm_output(9))) = '1' )
          THEN
        COMP_LOOP_acc_19_psp_sva <= z_out_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_14_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3297_nl, (fsm_output(10)), fsm_output(9))) = '1' )
          THEN
        COMP_LOOP_acc_1_cse_14_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1101")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_20_psp_sva <= STD_LOGIC_VECTOR'( "00000000000");
      ELSIF ( (MUX_s_1_2_2(nor_1420_nl, and_1254_nl, fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_20_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0(11
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "111")), 8), 11), 11));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3304_nl, and_816_cse, or_2935_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_11_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1111")), 9), 12), 12));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        modExp_exp_1_6_1_sva <= '0';
        modExp_exp_1_5_1_sva <= '0';
        modExp_exp_1_4_1_sva <= '0';
      ELSIF ( mux_3369_itm = '1' ) THEN
        modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0(2)), modExp_exp_1_7_1_sva,
            (COMP_LOOP_k_9_4_sva_4_0(3)), STD_LOGIC_VECTOR'( and_dcpl_283 & not_tmp_776
            & not_tmp_762));
        modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0(1)), modExp_exp_1_6_1_sva,
            (COMP_LOOP_k_9_4_sva_4_0(2)), STD_LOGIC_VECTOR'( and_dcpl_283 & not_tmp_776
            & not_tmp_762));
        modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0(0)), modExp_exp_1_5_1_sva,
            (COMP_LOOP_k_9_4_sva_4_0(1)), STD_LOGIC_VECTOR'( and_dcpl_283 & not_tmp_776
            & not_tmp_762));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_12_1_1_sva <= STD_LOGIC_VECTOR'( "000000000000");
      ELSIF ( COMP_LOOP_or_32_cse = '1' ) THEN
        COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_7(12 DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_126 OR not_tmp_519 OR and_dcpl_141 OR and_dcpl_158 OR and_dcpl_164
          OR and_dcpl_175 OR and_dcpl_192 OR and_dcpl_198 OR and_dcpl_206 OR and_dcpl_225
          OR and_dcpl_232 OR and_dcpl_242) = '1' ) THEN
        COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((z_out(9)), (z_out_8_8_7(1)),
            not_tmp_519);
      END IF;
    END IF;
  END PROCESS;
  modulo_result_or_nl <= and_dcpl_260 OR not_tmp_519;
  mux_2296_nl <= MUX_s_1_2_2(and_dcpl_123, (fsm_output(3)), and_573_cse);
  mux_2297_nl <= MUX_s_1_2_2(or_tmp_2233, (NOT mux_2296_nl), fsm_output(6));
  mux_2298_nl <= MUX_s_1_2_2(mux_2297_nl, mux_tmp_2220, fsm_output(7));
  mux_2295_nl <= MUX_s_1_2_2((NOT and_tmp_10), mux_tmp_2218, fsm_output(7));
  mux_2299_nl <= MUX_s_1_2_2((NOT mux_2298_nl), mux_2295_nl, fsm_output(5));
  mux_2291_nl <= MUX_s_1_2_2((fsm_output(3)), or_tmp_2260, fsm_output(1));
  mux_2292_nl <= MUX_s_1_2_2(mux_tmp_2254, mux_2291_nl, fsm_output(6));
  nand_264_nl <= NOT((fsm_output(6)) AND nor_tmp_295);
  mux_2293_nl <= MUX_s_1_2_2(mux_2292_nl, nand_264_nl, fsm_output(7));
  mux_2294_nl <= MUX_s_1_2_2(mux_2293_nl, mux_tmp_2290, fsm_output(5));
  mux_2300_nl <= MUX_s_1_2_2(mux_2299_nl, mux_2294_nl, fsm_output(2));
  mux_2286_nl <= MUX_s_1_2_2(mux_tmp_2285, or_tmp_2223, fsm_output(7));
  mux_2283_nl <= MUX_s_1_2_2(or_tmp_2230, (NOT nor_tmp_6), fsm_output(6));
  mux_2282_nl <= MUX_s_1_2_2(nor_tmp_295, (fsm_output(10)), fsm_output(6));
  mux_2284_nl <= MUX_s_1_2_2(mux_2283_nl, mux_2282_nl, fsm_output(7));
  mux_2287_nl <= MUX_s_1_2_2(mux_2286_nl, mux_2284_nl, fsm_output(5));
  mux_2278_nl <= MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, fsm_output(6));
  mux_2280_nl <= MUX_s_1_2_2(mux_28_cse, (NOT mux_2278_nl), fsm_output(7));
  nand_265_nl <= NOT((and_574_cse OR (fsm_output(3))) AND (fsm_output(10)));
  mux_2276_nl <= MUX_s_1_2_2((fsm_output(10)), or_tmp_2248, fsm_output(6));
  mux_2277_nl <= MUX_s_1_2_2(nand_265_nl, mux_2276_nl, fsm_output(7));
  mux_2281_nl <= MUX_s_1_2_2(mux_2280_nl, mux_2277_nl, fsm_output(5));
  mux_2288_nl <= MUX_s_1_2_2(mux_2287_nl, mux_2281_nl, fsm_output(2));
  mux_2301_nl <= MUX_s_1_2_2(mux_2300_nl, mux_2288_nl, fsm_output(8));
  mux_2272_nl <= MUX_s_1_2_2(or_tmp_14, nand_tmp_92, fsm_output(7));
  mux_2270_nl <= MUX_s_1_2_2((NOT (fsm_output(3))), nor_tmp_6, fsm_output(6));
  mux_2271_nl <= MUX_s_1_2_2(mux_2270_nl, or_tmp_14, fsm_output(7));
  mux_2273_nl <= MUX_s_1_2_2(mux_2272_nl, mux_2271_nl, fsm_output(5));
  mux_2267_nl <= MUX_s_1_2_2((NOT nor_tmp_291), mux_tmp_2250, fsm_output(6));
  mux_2268_nl <= MUX_s_1_2_2(or_tmp_2257, mux_2267_nl, fsm_output(7));
  mux_2266_nl <= MUX_s_1_2_2(mux_tmp_2265, or_tmp_2255, fsm_output(7));
  mux_2269_nl <= MUX_s_1_2_2(mux_2268_nl, mux_2266_nl, fsm_output(5));
  mux_2274_nl <= MUX_s_1_2_2(mux_2273_nl, mux_2269_nl, fsm_output(2));
  nor_778_nl <= NOT((fsm_output(6)) OR nor_tmp_6);
  mux_2261_nl <= MUX_s_1_2_2(nor_tmp_9, or_tmp_2253, fsm_output(6));
  mux_2262_nl <= MUX_s_1_2_2(nor_778_nl, mux_2261_nl, fsm_output(7));
  mux_2259_nl <= MUX_s_1_2_2(or_tmp_2253, (NOT mux_tmp_2251), fsm_output(6));
  mux_2258_nl <= MUX_s_1_2_2((NOT or_tmp_2238), nor_tmp_6, fsm_output(6));
  mux_2260_nl <= MUX_s_1_2_2(mux_2259_nl, mux_2258_nl, fsm_output(7));
  mux_2263_nl <= MUX_s_1_2_2(mux_2262_nl, mux_2260_nl, fsm_output(5));
  nor_779_nl <= NOT((fsm_output(6)) OR nor_tmp_9);
  mux_2255_nl <= MUX_s_1_2_2(or_tmp_2233, (NOT mux_tmp_2254), fsm_output(6));
  mux_2256_nl <= MUX_s_1_2_2(nor_779_nl, mux_2255_nl, fsm_output(7));
  mux_2252_nl <= MUX_s_1_2_2(mux_tmp_2251, mux_tmp_2250, fsm_output(6));
  mux_2253_nl <= MUX_s_1_2_2((NOT mux_2252_nl), and_tmp_10, fsm_output(7));
  mux_2257_nl <= MUX_s_1_2_2(mux_2256_nl, mux_2253_nl, fsm_output(5));
  mux_2264_nl <= MUX_s_1_2_2(mux_2263_nl, mux_2257_nl, fsm_output(2));
  mux_2275_nl <= MUX_s_1_2_2(mux_2274_nl, (NOT mux_2264_nl), fsm_output(8));
  mux_2302_nl <= MUX_s_1_2_2(mux_2301_nl, mux_2275_nl, fsm_output(4));
  mux_2245_nl <= MUX_s_1_2_2(mux_tmp_2239, nor_tmp_6, fsm_output(6));
  or_2306_nl <= (fsm_output(7)) OR mux_2245_nl;
  mux_2244_nl <= MUX_s_1_2_2(not_tmp_426, or_tmp_2246, fsm_output(7));
  mux_2246_nl <= MUX_s_1_2_2(or_2306_nl, mux_2244_nl, fsm_output(5));
  mux_2242_nl <= MUX_s_1_2_2(nor_tmp_286, or_tmp_2237, fsm_output(7));
  mux_2241_nl <= MUX_s_1_2_2(nand_tmp_92, or_tmp_14, fsm_output(7));
  mux_2243_nl <= MUX_s_1_2_2(mux_2242_nl, mux_2241_nl, fsm_output(5));
  mux_2247_nl <= MUX_s_1_2_2(mux_2246_nl, mux_2243_nl, fsm_output(2));
  mux_2235_nl <= MUX_s_1_2_2(or_tmp_2220, or_tmp_21, fsm_output(6));
  or_2300_nl <= (fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(10));
  mux_2236_nl <= MUX_s_1_2_2(mux_2235_nl, or_2300_nl, fsm_output(7));
  nand_91_nl <= NOT((fsm_output(7)) AND (NOT((((fsm_output(6)) OR (fsm_output(1)))
      AND (fsm_output(3))) OR (fsm_output(10)))));
  mux_2237_nl <= MUX_s_1_2_2(mux_2236_nl, nand_91_nl, fsm_output(5));
  mux_2233_nl <= MUX_s_1_2_2(or_tmp_237, or_tmp_2238, fsm_output(6));
  or_2297_nl <= (fsm_output(7)) OR mux_2233_nl;
  or_2293_nl <= ((fsm_output(6)) AND (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(10));
  mux_2232_nl <= MUX_s_1_2_2(or_tmp_2237, or_2293_nl, fsm_output(7));
  mux_2234_nl <= MUX_s_1_2_2(or_2297_nl, mux_2232_nl, fsm_output(5));
  mux_2238_nl <= MUX_s_1_2_2(mux_2237_nl, mux_2234_nl, fsm_output(2));
  mux_2248_nl <= MUX_s_1_2_2(mux_2247_nl, mux_2238_nl, fsm_output(8));
  mux_2225_nl <= MUX_s_1_2_2(and_dcpl_101, nor_tmp_6, fsm_output(1));
  mux_2226_nl <= MUX_s_1_2_2(and_dcpl_102, mux_2225_nl, fsm_output(0));
  mux_2227_nl <= MUX_s_1_2_2(and_dcpl_101, mux_2226_nl, fsm_output(6));
  mux_2228_nl <= MUX_s_1_2_2((NOT mux_2227_nl), or_tmp_4, fsm_output(7));
  mux_2224_nl <= MUX_s_1_2_2(mux_tmp_2223, or_tmp_2223, fsm_output(7));
  mux_2229_nl <= MUX_s_1_2_2(mux_2228_nl, mux_2224_nl, fsm_output(5));
  mux_2221_nl <= MUX_s_1_2_2((NOT mux_tmp_2220), or_tmp_4, fsm_output(7));
  or_2288_nl <= (fsm_output(6)) OR or_tmp_2230;
  mux_2219_nl <= MUX_s_1_2_2(mux_tmp_2218, or_2288_nl, fsm_output(7));
  mux_2222_nl <= MUX_s_1_2_2(mux_2221_nl, mux_2219_nl, fsm_output(5));
  mux_2230_nl <= MUX_s_1_2_2(mux_2229_nl, mux_2222_nl, fsm_output(2));
  or_2285_nl <= (NOT(and_574_cse OR (fsm_output(3)))) OR (fsm_output(10));
  mux_2215_nl <= MUX_s_1_2_2(or_tmp_14, or_2285_nl, fsm_output(7));
  mux_2214_nl <= MUX_s_1_2_2(or_tmp_2225, (fsm_output(10)), fsm_output(6));
  or_2283_nl <= (fsm_output(7)) OR mux_2214_nl;
  mux_2216_nl <= MUX_s_1_2_2(mux_2215_nl, or_2283_nl, fsm_output(5));
  or_2279_nl <= (NOT((fsm_output(3)) OR (fsm_output(6)))) OR (fsm_output(10));
  mux_2212_nl <= MUX_s_1_2_2(or_tmp_2223, or_2279_nl, fsm_output(7));
  nand_90_nl <= NOT((fsm_output(6)) AND (NOT or_tmp_2220));
  mux_2211_nl <= MUX_s_1_2_2((fsm_output(10)), nand_90_nl, fsm_output(7));
  mux_2213_nl <= MUX_s_1_2_2(mux_2212_nl, mux_2211_nl, fsm_output(5));
  mux_2217_nl <= MUX_s_1_2_2(mux_2216_nl, mux_2213_nl, fsm_output(2));
  mux_2231_nl <= MUX_s_1_2_2(mux_2230_nl, mux_2217_nl, fsm_output(8));
  mux_2249_nl <= MUX_s_1_2_2(mux_2248_nl, mux_2231_nl, fsm_output(4));
  mux_2303_nl <= MUX_s_1_2_2(mux_2302_nl, mux_2249_nl, fsm_output(9));
  or_2355_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(10));
  mux_2373_nl <= MUX_s_1_2_2(or_2355_nl, or_tmp_2267, fsm_output(7));
  mux_2372_nl <= MUX_s_1_2_2(or_tmp_2281, (NOT mux_tmp_2218), fsm_output(7));
  mux_2374_nl <= MUX_s_1_2_2(mux_2373_nl, mux_2372_nl, fsm_output(5));
  mux_2369_nl <= MUX_s_1_2_2((NOT nor_tmp_300), or_tmp_2271, fsm_output(6));
  or_2354_nl <= (fsm_output(6)) OR ((fsm_output(0)) AND (fsm_output(1)) AND (NOT
      (fsm_output(3))) AND (fsm_output(10)));
  mux_2370_nl <= MUX_s_1_2_2(mux_2369_nl, or_2354_nl, fsm_output(7));
  or_2351_nl <= (fsm_output(6)) OR and_dcpl_223;
  mux_2367_nl <= MUX_s_1_2_2(or_tmp_21, mux_tmp_2362, fsm_output(6));
  mux_2368_nl <= MUX_s_1_2_2(or_2351_nl, mux_2367_nl, fsm_output(7));
  mux_2371_nl <= MUX_s_1_2_2(mux_2370_nl, mux_2368_nl, fsm_output(5));
  mux_2375_nl <= MUX_s_1_2_2(mux_2374_nl, mux_2371_nl, fsm_output(2));
  mux_2364_nl <= MUX_s_1_2_2(mux_tmp_2285, (fsm_output(6)), fsm_output(7));
  nand_100_nl <= NOT((fsm_output(6)) AND (NOT mux_tmp_2362));
  mux_2363_nl <= MUX_s_1_2_2(nand_100_nl, or_tmp_2293, fsm_output(7));
  mux_2365_nl <= MUX_s_1_2_2((NOT mux_2364_nl), mux_2363_nl, fsm_output(5));
  nand_99_nl <= NOT((fsm_output(6)) AND (NOT mux_tmp_2239));
  mux_2360_nl <= MUX_s_1_2_2((NOT mux_28_cse), nand_99_nl, fsm_output(7));
  nand_98_nl <= NOT((fsm_output(6)) AND (NOT nor_tmp_295));
  mux_2359_nl <= MUX_s_1_2_2(nand_98_nl, or_tmp_434, fsm_output(7));
  mux_2361_nl <= MUX_s_1_2_2(mux_2360_nl, mux_2359_nl, fsm_output(5));
  mux_2366_nl <= MUX_s_1_2_2(mux_2365_nl, mux_2361_nl, fsm_output(2));
  mux_2376_nl <= MUX_s_1_2_2(mux_2375_nl, mux_2366_nl, fsm_output(8));
  mux_2354_nl <= MUX_s_1_2_2((fsm_output(10)), (NOT or_tmp_2248), fsm_output(6));
  mux_2355_nl <= MUX_s_1_2_2(mux_2354_nl, mux_tmp_2327, fsm_output(7));
  mux_2352_nl <= MUX_s_1_2_2(and_dcpl_109, nor_tmp_6, fsm_output(6));
  mux_2353_nl <= MUX_s_1_2_2(mux_2352_nl, and_tmp_16, fsm_output(7));
  mux_2356_nl <= MUX_s_1_2_2(mux_2355_nl, mux_2353_nl, fsm_output(5));
  nand_261_nl <= NOT(or_2348_cse AND mux_tmp_2239);
  mux_2348_nl <= MUX_s_1_2_2(nand_261_nl, nor_tmp_6, fsm_output(6));
  mux_2350_nl <= MUX_s_1_2_2((NOT mux_tmp_2349), mux_2348_nl, fsm_output(7));
  and_275_nl <= (fsm_output(6)) AND ((fsm_output(1)) OR (NOT (fsm_output(3))) OR
      (fsm_output(10)));
  mux_2347_nl <= MUX_s_1_2_2(mux_tmp_2265, and_275_nl, fsm_output(7));
  mux_2351_nl <= MUX_s_1_2_2(mux_2350_nl, mux_2347_nl, fsm_output(5));
  mux_2357_nl <= MUX_s_1_2_2(mux_2356_nl, mux_2351_nl, fsm_output(2));
  mux_2344_nl <= MUX_s_1_2_2(not_tmp_463, nand_tmp_96, fsm_output(7));
  or_2342_nl <= (fsm_output(1)) OR (NOT nor_tmp_6);
  mux_2342_nl <= MUX_s_1_2_2(or_tmp_2266, or_2342_nl, fsm_output(0));
  or_2343_nl <= (fsm_output(6)) OR (NOT mux_2342_nl);
  mux_2343_nl <= MUX_s_1_2_2(or_tmp_3, or_2343_nl, fsm_output(7));
  mux_2345_nl <= MUX_s_1_2_2(mux_2344_nl, mux_2343_nl, fsm_output(5));
  or_2341_nl <= (fsm_output(1)) OR (fsm_output(3)) OR (NOT (fsm_output(10)));
  mux_2339_nl <= MUX_s_1_2_2(or_2341_nl, or_tmp_2282, fsm_output(0));
  nand_262_nl <= NOT((fsm_output(6)) AND mux_2339_nl);
  mux_2340_nl <= MUX_s_1_2_2(nand_262_nl, or_tmp_3, fsm_output(7));
  mux_2337_nl <= MUX_s_1_2_2((NOT and_dcpl_240), or_tmp_2238, fsm_output(6));
  mux_2338_nl <= MUX_s_1_2_2(mux_2337_nl, or_tmp_2281, fsm_output(7));
  mux_2341_nl <= MUX_s_1_2_2(mux_2340_nl, mux_2338_nl, fsm_output(5));
  mux_2346_nl <= MUX_s_1_2_2(mux_2345_nl, mux_2341_nl, fsm_output(2));
  mux_2358_nl <= MUX_s_1_2_2((NOT mux_2357_nl), mux_2346_nl, fsm_output(8));
  mux_2377_nl <= MUX_s_1_2_2(mux_2376_nl, mux_2358_nl, fsm_output(4));
  mux_2332_nl <= MUX_s_1_2_2(or_36_cse, or_tmp_14, fsm_output(7));
  mux_2331_nl <= MUX_s_1_2_2(or_tmp_2280, or_15_cse, fsm_output(7));
  mux_2333_nl <= MUX_s_1_2_2(mux_2332_nl, mux_2331_nl, fsm_output(5));
  mux_2329_nl <= MUX_s_1_2_2(or_36_cse, or_tmp_2255, fsm_output(7));
  mux_2328_nl <= MUX_s_1_2_2((NOT mux_tmp_2327), or_tmp_4, fsm_output(7));
  mux_2330_nl <= MUX_s_1_2_2(mux_2329_nl, mux_2328_nl, fsm_output(5));
  mux_2334_nl <= MUX_s_1_2_2(mux_2333_nl, mux_2330_nl, fsm_output(2));
  mux_2323_nl <= MUX_s_1_2_2(or_tmp_2248, or_tmp_237, fsm_output(6));
  nand_97_nl <= NOT((fsm_output(6)) AND (NOT or_tmp_2275));
  mux_2324_nl <= MUX_s_1_2_2(mux_2323_nl, nand_97_nl, fsm_output(7));
  mux_2322_nl <= MUX_s_1_2_2(or_tmp_4, or_tmp_2276, fsm_output(7));
  mux_2325_nl <= MUX_s_1_2_2(mux_2324_nl, mux_2322_nl, fsm_output(5));
  mux_2319_nl <= MUX_s_1_2_2(or_tmp_21, or_tmp_2275, fsm_output(6));
  mux_2320_nl <= MUX_s_1_2_2(mux_2319_nl, or_tmp_4, fsm_output(7));
  mux_2318_nl <= MUX_s_1_2_2(nand_tmp_96, or_tmp_2246, fsm_output(7));
  mux_2321_nl <= MUX_s_1_2_2(mux_2320_nl, mux_2318_nl, fsm_output(5));
  mux_2326_nl <= MUX_s_1_2_2(mux_2325_nl, mux_2321_nl, fsm_output(2));
  mux_2335_nl <= MUX_s_1_2_2(mux_2334_nl, mux_2326_nl, fsm_output(8));
  or_2330_nl <= (fsm_output(6)) OR mux_tmp_2254;
  or_2329_nl <= (fsm_output(6)) OR or_tmp_2271;
  mux_2314_nl <= MUX_s_1_2_2(or_2330_nl, or_2329_nl, fsm_output(7));
  mux_2313_nl <= MUX_s_1_2_2((NOT mux_tmp_2223), nand_tmp_95, fsm_output(7));
  mux_2315_nl <= MUX_s_1_2_2(mux_2314_nl, mux_2313_nl, fsm_output(5));
  mux_2311_nl <= MUX_s_1_2_2(or_tmp_2267, or_tmp_14, fsm_output(7));
  nand_94_nl <= NOT((fsm_output(6)) AND (NOT or_tmp_2225));
  mux_2308_nl <= MUX_s_1_2_2((NOT mux_tmp_2218), nand_94_nl, fsm_output(7));
  mux_2312_nl <= MUX_s_1_2_2(mux_2311_nl, mux_2308_nl, fsm_output(5));
  mux_2316_nl <= MUX_s_1_2_2(mux_2315_nl, mux_2312_nl, fsm_output(2));
  mux_2305_nl <= MUX_s_1_2_2(or_tmp_3, nand_tmp_93, fsm_output(7));
  or_2321_nl <= (NOT (fsm_output(7))) OR (fsm_output(6)) OR (fsm_output(10));
  mux_2306_nl <= MUX_s_1_2_2(mux_2305_nl, or_2321_nl, fsm_output(5));
  or_2319_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")) OR or_tmp_2248;
  mux_2304_nl <= MUX_s_1_2_2(or_tmp_2263, or_2319_nl, fsm_output(5));
  mux_2307_nl <= MUX_s_1_2_2(mux_2306_nl, mux_2304_nl, fsm_output(2));
  mux_2317_nl <= MUX_s_1_2_2(mux_2316_nl, mux_2307_nl, fsm_output(8));
  mux_2336_nl <= MUX_s_1_2_2(mux_2335_nl, mux_2317_nl, fsm_output(4));
  mux_2378_nl <= MUX_s_1_2_2(mux_2377_nl, mux_2336_nl, fsm_output(9));
  nor_758_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(2)))
      OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(5)) OR (fsm_output(10)));
  nor_759_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(8))) OR (fsm_output(2)) OR
      (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10))));
  mux_2391_nl <= MUX_s_1_2_2(nor_758_nl, nor_759_nl, fsm_output(4));
  nor_760_nl <= NOT((fsm_output(8)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10)));
  nor_761_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(2)) OR (fsm_output(3)) OR
      (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_2390_nl <= MUX_s_1_2_2(nor_760_nl, nor_761_nl, fsm_output(7));
  and_568_nl <= (fsm_output(4)) AND mux_2390_nl;
  mux_2392_nl <= MUX_s_1_2_2(mux_2391_nl, and_568_nl, fsm_output(6));
  nor_762_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(2)))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  nor_763_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(8)) OR (fsm_output(2)) OR
      (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(5))) OR
      (fsm_output(10)));
  mux_2388_nl <= MUX_s_1_2_2(nor_762_nl, nor_763_nl, fsm_output(4));
  or_2372_nl <= (fsm_output(8)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT (fsm_output(10)));
  or_2370_nl <= (NOT (fsm_output(8))) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_45;
  mux_2387_nl <= MUX_s_1_2_2(or_2372_nl, or_2370_nl, fsm_output(7));
  nor_764_nl <= NOT((fsm_output(4)) OR mux_2387_nl);
  mux_2389_nl <= MUX_s_1_2_2(mux_2388_nl, nor_764_nl, fsm_output(6));
  mux_2393_nl <= MUX_s_1_2_2(mux_2392_nl, mux_2389_nl, fsm_output(1));
  nor_765_nl <= NOT((fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(5))
      OR (fsm_output(10)));
  nor_766_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_2384_nl <= MUX_s_1_2_2(nor_765_nl, nor_766_nl, fsm_output(8));
  and_570_nl <= (fsm_output(7)) AND mux_2384_nl;
  or_2365_nl <= (NOT (fsm_output(2))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (fsm_output(10));
  or_2364_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (fsm_output(9))
      OR not_tmp_45;
  mux_2383_nl <= MUX_s_1_2_2(or_2365_nl, or_2364_nl, fsm_output(8));
  nor_767_nl <= NOT((fsm_output(7)) OR mux_2383_nl);
  mux_2385_nl <= MUX_s_1_2_2(and_570_nl, nor_767_nl, fsm_output(4));
  and_569_nl <= (fsm_output(6)) AND mux_2385_nl;
  nor_768_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(8))) OR (fsm_output(2))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10)));
  nor_769_nl <= NOT((fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT
      (fsm_output(5))) OR (fsm_output(10)));
  nor_770_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (fsm_output(10)));
  mux_2379_nl <= MUX_s_1_2_2(nor_769_nl, nor_770_nl, fsm_output(8));
  nor_771_nl <= NOT((fsm_output(8)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(9))
      OR not_tmp_45);
  mux_2380_nl <= MUX_s_1_2_2(mux_2379_nl, nor_771_nl, fsm_output(7));
  mux_2381_nl <= MUX_s_1_2_2(nor_768_nl, mux_2380_nl, fsm_output(4));
  nor_772_nl <= NOT((fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(8)) OR (NOT
      (fsm_output(2))) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (NOT (fsm_output(10))));
  mux_2382_nl <= MUX_s_1_2_2(mux_2381_nl, nor_772_nl, fsm_output(6));
  mux_2386_nl <= MUX_s_1_2_2(and_569_nl, mux_2382_nl, fsm_output(1));
  mux_2394_nl <= MUX_s_1_2_2(mux_2393_nl, mux_2386_nl, fsm_output(0));
  nand_109_nl <= NOT((fsm_output(5)) AND (NOT mux_tmp_2425));
  mux_2456_nl <= MUX_s_1_2_2(nand_109_nl, nand_tmp_108, or_2348_cse);
  mux_2455_nl <= MUX_s_1_2_2(nand_tmp_108, nand_tmp_107, and_573_cse);
  mux_2457_nl <= MUX_s_1_2_2(mux_2456_nl, mux_2455_nl, fsm_output(2));
  mux_2452_nl <= MUX_s_1_2_2((NOT or_tmp_2342), mux_tmp_2426, fsm_output(0));
  mux_2453_nl <= MUX_s_1_2_2((NOT or_tmp_2343), mux_2452_nl, fsm_output(1));
  mux_2451_nl <= MUX_s_1_2_2(mux_tmp_2426, mux_tmp_2436, fsm_output(1));
  mux_2454_nl <= MUX_s_1_2_2(mux_2453_nl, mux_2451_nl, fsm_output(2));
  mux_2458_nl <= MUX_s_1_2_2(mux_2457_nl, (NOT mux_2454_nl), fsm_output(7));
  mux_2447_nl <= MUX_s_1_2_2(mux_tmp_2401, (NOT nor_tmp_307), fsm_output(5));
  mux_2446_nl <= MUX_s_1_2_2(mux_tmp_2401, nand_257_cse, fsm_output(5));
  mux_2448_nl <= MUX_s_1_2_2(mux_2447_nl, mux_2446_nl, or_2348_cse);
  mux_2443_nl <= MUX_s_1_2_2(or_tmp_434, (NOT (fsm_output(6))), fsm_output(8));
  mux_2444_nl <= MUX_s_1_2_2(or_tmp_2334, mux_2443_nl, fsm_output(5));
  mux_2445_nl <= MUX_s_1_2_2(mux_2444_nl, mux_tmp_2423, or_2348_cse);
  mux_2449_nl <= MUX_s_1_2_2(mux_2448_nl, mux_2445_nl, fsm_output(2));
  mux_2450_nl <= MUX_s_1_2_2(mux_tmp_2406, mux_2449_nl, fsm_output(7));
  mux_2459_nl <= MUX_s_1_2_2(mux_2458_nl, mux_2450_nl, fsm_output(4));
  mux_2439_nl <= MUX_s_1_2_2(nand_tmp_107, nand_tmp_105, and_573_cse);
  mux_2438_nl <= MUX_s_1_2_2(nand_tmp_105, mux_tmp_2406, and_573_cse);
  mux_2440_nl <= MUX_s_1_2_2(mux_2439_nl, mux_2438_nl, fsm_output(2));
  mux_2434_nl <= MUX_s_1_2_2((NOT mux_2433_itm), nor_tmp_307, fsm_output(5));
  mux_2437_nl <= MUX_s_1_2_2(mux_tmp_2436, mux_2434_nl, fsm_output(2));
  mux_2441_nl <= MUX_s_1_2_2(mux_2440_nl, (NOT mux_2437_nl), fsm_output(7));
  mux_2430_nl <= MUX_s_1_2_2(mux_tmp_2406, or_tmp_2343, or_2348_cse);
  mux_2428_nl <= MUX_s_1_2_2(or_tmp_2343, or_tmp_2342, fsm_output(0));
  mux_2429_nl <= MUX_s_1_2_2(mux_2428_nl, (NOT mux_tmp_2426), fsm_output(1));
  mux_2431_nl <= MUX_s_1_2_2(mux_2430_nl, mux_2429_nl, fsm_output(2));
  nand_106_nl <= NOT((fsm_output(5)) AND (NOT mux_tmp_917));
  mux_2424_nl <= MUX_s_1_2_2(mux_tmp_2423, nand_106_nl, and_563_cse);
  mux_2432_nl <= MUX_s_1_2_2(mux_2431_nl, mux_2424_nl, fsm_output(7));
  mux_2442_nl <= MUX_s_1_2_2(mux_2441_nl, mux_2432_nl, fsm_output(4));
  mux_2460_nl <= MUX_s_1_2_2(mux_2459_nl, mux_2442_nl, fsm_output(3));
  or_2397_nl <= (fsm_output(8)) OR (fsm_output(6)) OR (fsm_output(10));
  mux_2416_nl <= MUX_s_1_2_2(or_2397_nl, mux_tmp_2401, fsm_output(5));
  mux_2417_nl <= MUX_s_1_2_2(mux_2416_nl, nand_tmp_105, and_573_cse);
  mux_2418_nl <= MUX_s_1_2_2(mux_2417_nl, nand_tmp_105, fsm_output(2));
  mux_2414_nl <= MUX_s_1_2_2(or_tmp_2329, or_tmp_2335, or_2348_cse);
  mux_2415_nl <= MUX_s_1_2_2(or_tmp_2329, mux_2414_nl, fsm_output(2));
  mux_2419_nl <= MUX_s_1_2_2(mux_2418_nl, mux_2415_nl, fsm_output(7));
  mux_2411_nl <= MUX_s_1_2_2(mux_tmp_2406, or_tmp_2338, fsm_output(1));
  mux_2410_nl <= MUX_s_1_2_2(or_tmp_2338, or_tmp_2331, fsm_output(1));
  mux_2412_nl <= MUX_s_1_2_2(mux_2411_nl, mux_2410_nl, fsm_output(2));
  mux_2409_nl <= MUX_s_1_2_2(mux_tmp_2400, or_tmp_2327, and_565_cse);
  mux_2413_nl <= MUX_s_1_2_2(mux_2412_nl, mux_2409_nl, fsm_output(7));
  mux_2420_nl <= MUX_s_1_2_2(mux_2419_nl, mux_2413_nl, fsm_output(4));
  mux_2404_nl <= MUX_s_1_2_2(or_tmp_2335, mux_tmp_2402, fsm_output(1));
  mux_2403_nl <= MUX_s_1_2_2(mux_tmp_2402, mux_tmp_2400, or_2348_cse);
  mux_2405_nl <= MUX_s_1_2_2(mux_2404_nl, mux_2403_nl, fsm_output(2));
  mux_2407_nl <= MUX_s_1_2_2(mux_tmp_2406, mux_2405_nl, fsm_output(7));
  mux_2398_nl <= MUX_s_1_2_2(or_tmp_2331, or_tmp_2329, or_2385_cse);
  mux_2395_nl <= MUX_s_1_2_2(or_tmp_14, or_tmp_4, fsm_output(8));
  nand_104_nl <= NOT((fsm_output(5)) AND (NOT mux_2395_nl));
  mux_2396_nl <= MUX_s_1_2_2(or_tmp_2327, nand_104_nl, and_573_cse);
  or_2381_nl <= (NOT (fsm_output(5))) OR (fsm_output(8)) OR (fsm_output(6)) OR (fsm_output(10));
  mux_2397_nl <= MUX_s_1_2_2(mux_2396_nl, or_2381_nl, fsm_output(2));
  mux_2399_nl <= MUX_s_1_2_2(mux_2398_nl, mux_2397_nl, fsm_output(7));
  mux_2408_nl <= MUX_s_1_2_2(mux_2407_nl, mux_2399_nl, fsm_output(4));
  mux_2421_nl <= MUX_s_1_2_2(mux_2420_nl, mux_2408_nl, fsm_output(3));
  mux_2461_nl <= MUX_s_1_2_2(mux_2460_nl, mux_2421_nl, fsm_output(9));
  COMP_LOOP_nor_11_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_and_274_nl <= (NOT and_dcpl_281) AND and_dcpl_273;
  or_2728_nl <= (fsm_output(8)) OR ((fsm_output(4)) AND or_tmp_187);
  mux_2971_nl <= MUX_s_1_2_2(or_2729_cse, or_2728_nl, fsm_output(1));
  mux_2972_nl <= MUX_s_1_2_2(mux_tmp_413, mux_2971_nl, fsm_output(6));
  mux_2969_nl <= MUX_s_1_2_2(mux_tmp_2930, mux_tmp_2907, or_2348_cse);
  mux_2970_nl <= MUX_s_1_2_2(mux_2969_nl, nand_tmp_140, fsm_output(6));
  mux_2973_nl <= MUX_s_1_2_2(mux_2972_nl, mux_2970_nl, fsm_output(7));
  mux_2965_nl <= MUX_s_1_2_2((NOT mux_tmp_2911), or_tmp_182, fsm_output(8));
  mux_2966_nl <= MUX_s_1_2_2(mux_2965_nl, or_tmp_2663, and_573_cse);
  mux_2964_nl <= MUX_s_1_2_2(nand_tmp_140, nand_tmp_13, fsm_output(1));
  mux_2967_nl <= MUX_s_1_2_2(mux_2966_nl, mux_2964_nl, fsm_output(6));
  mux_2963_nl <= MUX_s_1_2_2(or_tmp_189, mux_tmp_2930, fsm_output(6));
  mux_2968_nl <= MUX_s_1_2_2(mux_2967_nl, mux_2963_nl, fsm_output(7));
  mux_2974_nl <= MUX_s_1_2_2(mux_2973_nl, mux_2968_nl, fsm_output(5));
  mux_426_nl <= MUX_s_1_2_2(or_tmp_187, nor_tmp_46, fsm_output(8));
  mux_427_nl <= MUX_s_1_2_2(mux_tmp_412, mux_426_nl, fsm_output(1));
  mux_2956_nl <= MUX_s_1_2_2(mux_tmp_2912, mux_tmp_2919, fsm_output(1));
  mux_2957_nl <= MUX_s_1_2_2(mux_tmp_2913, mux_2956_nl, fsm_output(0));
  mux_2960_nl <= MUX_s_1_2_2(mux_427_nl, mux_2957_nl, fsm_output(6));
  mux_2955_nl <= MUX_s_1_2_2(mux_tmp_2905, nand_tmp_13, fsm_output(6));
  mux_2961_nl <= MUX_s_1_2_2(mux_2960_nl, mux_2955_nl, fsm_output(7));
  mux_421_nl <= MUX_s_1_2_2(nand_tmp_13, nand_tmp_12, fsm_output(1));
  mux_422_nl <= MUX_s_1_2_2(or_tmp_191, mux_421_nl, fsm_output(6));
  mux_2950_nl <= MUX_s_1_2_2(or_tmp_2659, mux_tmp_2912, or_2348_cse);
  mux_2951_nl <= MUX_s_1_2_2(mux_2950_nl, mux_tmp_2907, fsm_output(6));
  mux_2954_nl <= MUX_s_1_2_2(mux_422_nl, mux_2951_nl, fsm_output(7));
  mux_2962_nl <= MUX_s_1_2_2(mux_2961_nl, mux_2954_nl, fsm_output(5));
  mux_2975_nl <= MUX_s_1_2_2(mux_2974_nl, mux_2962_nl, fsm_output(3));
  mux_414_nl <= MUX_s_1_2_2(mux_tmp_413, mux_tmp_412, or_2348_cse);
  mux_2940_nl <= MUX_s_1_2_2(mux_726_cse, or_tmp_187, fsm_output(4));
  mux_2941_nl <= MUX_s_1_2_2(mux_2940_nl, or_tmp_2652, fsm_output(8));
  mux_2942_nl <= MUX_s_1_2_2(mux_tmp_2912, mux_2941_nl, nor_412_cse);
  mux_2946_nl <= MUX_s_1_2_2(mux_414_nl, mux_2942_nl, fsm_output(6));
  mux_2938_nl <= MUX_s_1_2_2(nand_tmp_140, nand_tmp_13, and_573_cse);
  mux_2939_nl <= MUX_s_1_2_2(mux_tmp_2907, mux_2938_nl, fsm_output(6));
  mux_2947_nl <= MUX_s_1_2_2(mux_2946_nl, mux_2939_nl, fsm_output(7));
  mux_2934_nl <= MUX_s_1_2_2(or_tmp_2663, or_tmp_191, or_2348_cse);
  mux_2935_nl <= MUX_s_1_2_2(mux_2934_nl, nand_tmp_13, fsm_output(6));
  mux_2932_nl <= MUX_s_1_2_2(or_tmp_189, or_tmp_2659, and_573_cse);
  mux_2931_nl <= MUX_s_1_2_2(mux_tmp_2930, mux_tmp_2907, fsm_output(1));
  mux_2933_nl <= MUX_s_1_2_2(mux_2932_nl, mux_2931_nl, fsm_output(6));
  mux_2936_nl <= MUX_s_1_2_2(mux_2935_nl, mux_2933_nl, fsm_output(7));
  mux_2948_nl <= MUX_s_1_2_2(mux_2947_nl, mux_2936_nl, fsm_output(5));
  or_2718_nl <= (NOT (fsm_output(8))) OR (fsm_output(4));
  mux_2924_nl <= MUX_s_1_2_2(and_816_cse, or_tmp_187, or_2718_nl);
  mux_2925_nl <= MUX_s_1_2_2(mux_2924_nl, mux_tmp_2921, fsm_output(1));
  mux_2922_nl <= MUX_s_1_2_2(or_tmp_182, mux_tmp_2911, fsm_output(8));
  mux_2923_nl <= MUX_s_1_2_2(mux_2922_nl, mux_tmp_2921, fsm_output(1));
  mux_2926_nl <= MUX_s_1_2_2(mux_2925_nl, mux_2923_nl, fsm_output(0));
  mux_2927_nl <= MUX_s_1_2_2(mux_2926_nl, mux_tmp_2919, fsm_output(6));
  mux_386_nl <= MUX_s_1_2_2(nand_tmp_13, nand_tmp_12, and_573_cse);
  mux_2918_nl <= MUX_s_1_2_2(or_tmp_2649, mux_386_nl, fsm_output(6));
  mux_2928_nl <= MUX_s_1_2_2(mux_2927_nl, mux_2918_nl, fsm_output(7));
  mux_2908_nl <= MUX_s_1_2_2(mux_tmp_2907, nand_tmp_136, fsm_output(1));
  mux_2909_nl <= MUX_s_1_2_2(mux_2908_nl, mux_tmp_2905, fsm_output(0));
  mux_2914_nl <= MUX_s_1_2_2(mux_tmp_2913, mux_2909_nl, fsm_output(6));
  mux_2916_nl <= MUX_s_1_2_2(mux_384_cse, mux_2914_nl, fsm_output(7));
  mux_2929_nl <= MUX_s_1_2_2(mux_2928_nl, mux_2916_nl, fsm_output(5));
  mux_2949_nl <= MUX_s_1_2_2(mux_2948_nl, mux_2929_nl, fsm_output(3));
  mux_2976_nl <= MUX_s_1_2_2(mux_2975_nl, mux_2949_nl, fsm_output(2));
  COMP_LOOP_mux1h_428_nl <= MUX1HOT_s_1_6_2((operator_66_true_div_cmp_z(0)), (tmp_10_lpi_4_dfm(0)),
      (z_out_6(5)), COMP_LOOP_nor_12_itm, COMP_LOOP_nor_11_itm, COMP_LOOP_nor_11_nl,
      STD_LOGIC_VECTOR'( COMP_LOOP_and_274_nl & and_dcpl_281 & and_dcpl_119 & not_tmp_646
      & (NOT mux_2976_nl) & COMP_LOOP_or_32_cse));
  or_3351_nl <= (fsm_output(4)) OR (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(3))
      OR (fsm_output(8)) OR (fsm_output(9)) OR not_tmp_45;
  or_2678_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_45;
  mux_2885_nl <= MUX_s_1_2_2(or_2679_cse, or_2678_nl, fsm_output(3));
  nor_667_nl <= NOT((fsm_output(6)) OR mux_2885_nl);
  nor_668_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(8))
      OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_2886_nl <= MUX_s_1_2_2(nor_667_nl, nor_668_nl, fsm_output(2));
  nand_421_nl <= NOT((fsm_output(4)) AND mux_2886_nl);
  mux_2887_nl <= MUX_s_1_2_2(or_3351_nl, nand_421_nl, fsm_output(7));
  or_2674_nl <= (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(9)) OR (NOT (fsm_output(5)))
      OR (fsm_output(10));
  or_2673_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(9)))
      OR (fsm_output(5)) OR (fsm_output(10));
  mux_2883_nl <= MUX_s_1_2_2(or_2674_nl, or_2673_nl, fsm_output(6));
  or_3352_nl <= (NOT (fsm_output(4))) OR (fsm_output(2)) OR mux_2883_nl;
  nor_671_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_45);
  mux_2882_nl <= MUX_s_1_2_2(nor_670_cse, nor_671_nl, fsm_output(3));
  nand_422_nl <= NOT(nor_381_cse AND mux_2882_nl);
  mux_2884_nl <= MUX_s_1_2_2(or_3352_nl, nand_422_nl, fsm_output(7));
  mux_2888_nl <= MUX_s_1_2_2(mux_2887_nl, mux_2884_nl, fsm_output(1));
  nor_646_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (fsm_output(5)) OR (NOT (fsm_output(10))));
  nor_647_nl <= NOT((fsm_output(7)) OR (fsm_output(1)) OR (fsm_output(3)) OR (NOT
      (fsm_output(6))) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_2980_nl <= MUX_s_1_2_2(nor_646_nl, nor_647_nl, fsm_output(8));
  nor_648_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(7)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(5)) OR (NOT (fsm_output(10))));
  mux_2981_nl <= MUX_s_1_2_2(mux_2980_nl, nor_648_nl, fsm_output(4));
  nor_649_nl <= NOT((fsm_output(4)) OR (fsm_output(8)) OR (fsm_output(7)) OR (NOT
      (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(5)))
      OR (fsm_output(10)));
  mux_2982_nl <= MUX_s_1_2_2(mux_2981_nl, nor_649_nl, fsm_output(9));
  nor_650_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(8)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(5))
      OR (fsm_output(10)));
  nor_651_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR
      (fsm_output(5)) OR (NOT (fsm_output(10))));
  nor_652_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (NOT (fsm_output(6))) OR
      (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_2977_nl <= MUX_s_1_2_2(nor_651_nl, nor_652_nl, fsm_output(7));
  nor_653_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_2978_nl <= MUX_s_1_2_2(mux_2977_nl, nor_653_nl, fsm_output(8));
  and_490_nl <= (fsm_output(4)) AND mux_2978_nl;
  mux_2979_nl <= MUX_s_1_2_2(nor_650_nl, and_490_nl, fsm_output(9));
  mux_2983_nl <= MUX_s_1_2_2(mux_2982_nl, mux_2979_nl, fsm_output(2));
  COMP_LOOP_mux1h_464_nl <= MUX1HOT_s_1_4_2((COMP_LOOP_k_9_4_sva_4_0(3)), COMP_LOOP_nor_134_itm,
      modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_4_sva_4_0(4)), STD_LOGIC_VECTOR'( and_dcpl_283
      & and_dcpl_332 & (NOT mux_3369_itm) & not_tmp_762));
  nor_580_nl <= NOT((fsm_output(6)) OR mux_3394_cse);
  mux_3395_nl <= MUX_s_1_2_2(nor_580_nl, mux_3392_cse, fsm_output(3));
  mux_3396_nl <= MUX_s_1_2_2(mux_3395_nl, mux_3388_cse, fsm_output(9));
  COMP_LOOP_nor_12_nl <= NOT((z_out_7(4)) OR (z_out_7(3)) OR (z_out_7(1)));
  mux_3487_nl <= MUX_s_1_2_2(mux_tmp_3452, mux_tmp_3450, and_573_cse);
  mux_3486_nl <= MUX_s_1_2_2(mux_tmp_3450, mux_tmp_3449, or_2348_cse);
  mux_3488_nl <= MUX_s_1_2_2(mux_3487_nl, mux_3486_nl, fsm_output(2));
  mux_3483_nl <= MUX_s_1_2_2((NOT or_212_cse), and_tmp_36, fsm_output(5));
  mux_3482_nl <= MUX_s_1_2_2((NOT or_212_cse), (fsm_output(8)), fsm_output(5));
  mux_3484_nl <= MUX_s_1_2_2(mux_3483_nl, mux_3482_nl, fsm_output(1));
  mux_3480_nl <= MUX_s_1_2_2(mux_tmp_3456, (fsm_output(8)), fsm_output(5));
  mux_3481_nl <= MUX_s_1_2_2(mux_3480_nl, mux_tmp_3471, fsm_output(1));
  mux_3485_nl <= MUX_s_1_2_2(mux_3484_nl, mux_3481_nl, fsm_output(2));
  mux_3489_nl <= MUX_s_1_2_2(mux_3488_nl, (NOT mux_3485_nl), fsm_output(6));
  mux_3478_nl <= MUX_s_1_2_2(mux_tmp_3426, or_2729_cse, fsm_output(5));
  mux_3476_nl <= MUX_s_1_2_2((NOT and_tmp_36), mux_tmp_3426, fsm_output(5));
  mux_3477_nl <= MUX_s_1_2_2(mux_3476_nl, mux_tmp_3452, and_565_cse);
  mux_3479_nl <= MUX_s_1_2_2(mux_3478_nl, mux_3477_nl, fsm_output(6));
  mux_3490_nl <= MUX_s_1_2_2(mux_3489_nl, mux_3479_nl, fsm_output(7));
  mux_3469_nl <= MUX_s_1_2_2((NOT mux_tmp_3468), nand_tmp_167, fsm_output(5));
  mux_3470_nl <= MUX_s_1_2_2(mux_3469_nl, mux_tmp_3467, fsm_output(0));
  mux_3472_nl <= MUX_s_1_2_2((NOT mux_tmp_3471), mux_3470_nl, fsm_output(1));
  mux_3473_nl <= MUX_s_1_2_2(mux_3472_nl, mux_tmp_3467, fsm_output(2));
  mux_3474_nl <= MUX_s_1_2_2(mux_tmp_3449, mux_3473_nl, fsm_output(6));
  mux_3462_nl <= MUX_s_1_2_2(or_tmp_150, or_2729_cse, fsm_output(5));
  mux_3461_nl <= MUX_s_1_2_2((NOT or_tmp_150), mux_tmp_3458, fsm_output(5));
  mux_3463_nl <= MUX_s_1_2_2((NOT mux_3462_nl), mux_3461_nl, fsm_output(0));
  mux_3464_nl <= MUX_s_1_2_2(mux_3463_nl, mux_tmp_3459, fsm_output(1));
  mux_3457_nl <= MUX_s_1_2_2((NOT or_tmp_191), mux_tmp_3456, fsm_output(5));
  mux_3460_nl <= MUX_s_1_2_2(mux_tmp_3459, mux_3457_nl, fsm_output(1));
  mux_3465_nl <= MUX_s_1_2_2(mux_3464_nl, mux_3460_nl, fsm_output(2));
  mux_3453_nl <= MUX_s_1_2_2(mux_tmp_3452, mux_tmp_3450, fsm_output(0));
  mux_3451_nl <= MUX_s_1_2_2(mux_tmp_3450, mux_tmp_3449, fsm_output(0));
  mux_3454_nl <= MUX_s_1_2_2(mux_3453_nl, mux_3451_nl, fsm_output(1));
  mux_3455_nl <= MUX_s_1_2_2(mux_tmp_3452, mux_3454_nl, fsm_output(2));
  mux_3466_nl <= MUX_s_1_2_2((NOT mux_3465_nl), mux_3455_nl, fsm_output(6));
  mux_3475_nl <= MUX_s_1_2_2(mux_3474_nl, mux_3466_nl, fsm_output(7));
  mux_3491_nl <= MUX_s_1_2_2(mux_3490_nl, mux_3475_nl, fsm_output(3));
  mux_3443_nl <= MUX_s_1_2_2(or_2729_cse, or_tmp_118, fsm_output(5));
  mux_3442_nl <= MUX_s_1_2_2(or_212_cse, or_tmp_118, fsm_output(5));
  mux_3444_nl <= MUX_s_1_2_2(mux_3443_nl, mux_3442_nl, fsm_output(1));
  mux_3445_nl <= MUX_s_1_2_2(mux_3444_nl, mux_tmp_226, fsm_output(2));
  mux_3446_nl <= MUX_s_1_2_2(mux_tmp_3430, mux_3445_nl, fsm_output(6));
  mux_3438_nl <= MUX_s_1_2_2(or_163_cse, or_tmp_110, fsm_output(5));
  mux_3439_nl <= MUX_s_1_2_2(mux_3438_nl, mux_tmp_3436, or_2348_cse);
  mux_3437_nl <= MUX_s_1_2_2(mux_tmp_3436, mux_tmp_207, and_573_cse);
  mux_3440_nl <= MUX_s_1_2_2(mux_3439_nl, mux_3437_nl, fsm_output(2));
  mux_3434_nl <= MUX_s_1_2_2(or_tmp_118, or_163_cse, fsm_output(5));
  mux_3435_nl <= MUX_s_1_2_2(mux_3434_nl, mux_tmp_3418, and_563_cse);
  mux_3441_nl <= MUX_s_1_2_2(mux_3440_nl, mux_3435_nl, fsm_output(6));
  mux_3447_nl <= MUX_s_1_2_2(mux_3446_nl, mux_3441_nl, fsm_output(7));
  mux_3428_nl <= MUX_s_1_2_2(or_163_cse, (fsm_output(8)), fsm_output(5));
  mux_3427_nl <= MUX_s_1_2_2(mux_tmp_3426, (fsm_output(8)), fsm_output(5));
  mux_3429_nl <= MUX_s_1_2_2(mux_3428_nl, mux_3427_nl, fsm_output(1));
  mux_3431_nl <= MUX_s_1_2_2(mux_tmp_3430, mux_3429_nl, fsm_output(2));
  mux_3424_nl <= MUX_s_1_2_2(mux_tmp_226, mux_tmp_3422, and_573_cse);
  mux_3425_nl <= MUX_s_1_2_2(mux_3424_nl, mux_tmp_3422, fsm_output(2));
  mux_3432_nl <= MUX_s_1_2_2(mux_3431_nl, mux_3425_nl, fsm_output(6));
  mux_3420_nl <= MUX_s_1_2_2(mux_tmp_207, mux_tmp_3418, fsm_output(6));
  mux_3433_nl <= MUX_s_1_2_2(mux_3432_nl, mux_3420_nl, fsm_output(7));
  mux_3448_nl <= MUX_s_1_2_2(mux_3447_nl, mux_3433_nl, fsm_output(3));
  mux_3492_nl <= MUX_s_1_2_2(mux_3491_nl, mux_3448_nl, fsm_output(9));
  or_3090_nl <= (fsm_output(6)) OR mux_3394_cse;
  or_3084_nl <= (fsm_output(0)) OR mux_tmp_3386;
  or_3083_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR (fsm_output(2))
      OR (fsm_output(7)) OR not_tmp_34;
  mux_3499_nl <= MUX_s_1_2_2(or_3002_cse, mux_3498_cse, fsm_output(1));
  or_3079_nl <= (fsm_output(1)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  mux_3500_nl <= MUX_s_1_2_2(mux_3499_nl, or_3079_nl, fsm_output(5));
  mux_3501_nl <= MUX_s_1_2_2(or_3083_nl, mux_3500_nl, fsm_output(0));
  mux_3502_nl <= MUX_s_1_2_2(or_3084_nl, mux_3501_nl, fsm_output(6));
  mux_3505_nl <= MUX_s_1_2_2(or_3090_nl, mux_3502_nl, fsm_output(3));
  nand_168_nl <= NOT((fsm_output(0)) AND (NOT mux_tmp_3386));
  or_3076_nl <= (fsm_output(0)) OR mux_3385_cse;
  mux_3496_nl <= MUX_s_1_2_2(nand_168_nl, or_3076_nl, fsm_output(6));
  or_3071_nl <= (fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR (NOT (fsm_output(2))) OR (fsm_output(7)) OR (NOT (fsm_output(8))) OR (NOT
      (fsm_output(4))) OR (fsm_output(10));
  mux_3497_nl <= MUX_s_1_2_2(mux_3496_nl, or_3071_nl, fsm_output(3));
  mux_3506_nl <= MUX_s_1_2_2(mux_3505_nl, mux_3497_nl, fsm_output(9));
  COMP_LOOP_mux1h_474_nl <= MUX1HOT_s_1_3_2(COMP_LOOP_nor_12_itm, COMP_LOOP_nor_134_itm,
      COMP_LOOP_nor_12_nl, STD_LOGIC_VECTOR'( (NOT mux_3492_nl) & (NOT mux_3506_nl)
      & COMP_LOOP_or_32_cse));
  or_3055_nl <= (fsm_output(6)) OR (fsm_output(8)) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(0))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(10));
  or_3054_nl <= (fsm_output(8)) OR (NOT (fsm_output(5))) OR (fsm_output(0)) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(10));
  or_3052_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(10));
  or_3051_nl <= (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(10)));
  mux_3414_nl <= MUX_s_1_2_2(or_3052_nl, or_3051_nl, fsm_output(0));
  or_3053_nl <= (NOT (fsm_output(8))) OR (fsm_output(5)) OR mux_3414_nl;
  mux_3415_nl <= MUX_s_1_2_2(or_3054_nl, or_3053_nl, fsm_output(6));
  mux_3416_nl <= MUX_s_1_2_2(or_3055_nl, mux_3415_nl, fsm_output(4));
  nor_569_nl <= NOT((fsm_output(7)) OR mux_3416_nl);
  nor_570_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (NOT (fsm_output(10))));
  nor_571_nl <= NOT((fsm_output(5)) OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(10)));
  mux_3412_nl <= MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output(8));
  and_410_nl <= (fsm_output(6)) AND mux_3412_nl;
  or_3044_nl <= (fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(3)) OR (fsm_output(9))
      OR (fsm_output(10));
  nand_208_nl <= NOT((fsm_output(5)) AND (fsm_output(0)) AND (fsm_output(3)) AND
      (fsm_output(9)) AND (NOT (fsm_output(10))));
  mux_3411_nl <= MUX_s_1_2_2(or_3044_nl, nand_208_nl, fsm_output(8));
  nor_572_nl <= NOT((fsm_output(6)) OR mux_3411_nl);
  mux_3413_nl <= MUX_s_1_2_2(and_410_nl, nor_572_nl, fsm_output(4));
  and_409_nl <= (fsm_output(7)) AND mux_3413_nl;
  mux_3417_nl <= MUX_s_1_2_2(nor_569_nl, and_409_nl, fsm_output(2));
  or_3348_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(5))) OR (fsm_output(3)) OR (fsm_output(8)) OR (NOT (fsm_output(10)));
  or_3099_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (fsm_output(3))
      OR (NOT (fsm_output(8))) OR (fsm_output(10));
  mux_3510_nl <= MUX_s_1_2_2(or_3099_nl, or_tmp_3025, fsm_output(7));
  or_3349_nl <= (fsm_output(2)) OR mux_3510_nl;
  mux_3511_nl <= MUX_s_1_2_2(or_3348_nl, or_3349_nl, fsm_output(0));
  or_3097_nl <= (NOT (fsm_output(7))) OR (fsm_output(6)) OR (NOT((fsm_output(5))
      AND (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(10))));
  or_3095_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(10));
  mux_3509_nl <= MUX_s_1_2_2(or_3097_nl, or_3095_nl, fsm_output(2));
  or_3350_nl <= (fsm_output(0)) OR mux_3509_nl;
  mux_3512_nl <= MUX_s_1_2_2(mux_3511_nl, or_3350_nl, fsm_output(4));
  nor_567_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(6)) OR
      (fsm_output(5)) OR (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(10)));
  or_3091_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (fsm_output(3))
      OR (fsm_output(8)) OR (fsm_output(10));
  mux_3507_nl <= MUX_s_1_2_2(or_tmp_3025, or_3091_nl, fsm_output(7));
  and_402_nl <= (fsm_output(2)) AND (NOT mux_3507_nl);
  mux_3508_nl <= MUX_s_1_2_2(nor_567_nl, and_402_nl, fsm_output(0));
  nand_420_nl <= NOT((fsm_output(4)) AND mux_3508_nl);
  mux_3513_nl <= MUX_s_1_2_2(mux_3512_nl, nand_420_nl, fsm_output(9));
  COMP_LOOP_nor_14_nl <= NOT((z_out_7(4)) OR (z_out_7(2)) OR (z_out_7(1)));
  mux_3558_nl <= MUX_s_1_2_2(mux_tmp_379, mux_tmp_3323, fsm_output(1));
  mux_3559_nl <= MUX_s_1_2_2(mux_382_cse, mux_3558_nl, fsm_output(0));
  mux_3560_nl <= MUX_s_1_2_2(nand_tmp_12, mux_3559_nl, fsm_output(6));
  mux_3561_nl <= MUX_s_1_2_2(mux_3560_nl, mux_3557_cse, fsm_output(5));
  mux_3562_nl <= MUX_s_1_2_2(mux_3561_nl, mux_3555_cse, fsm_output(7));
  mux_3576_nl <= MUX_s_1_2_2(mux_3575_cse, mux_3562_nl, fsm_output(3));
  mux_3577_nl <= MUX_s_1_2_2(mux_3576_nl, mux_3551_cse, fsm_output(2));
  COMP_LOOP_mux1h_477_nl <= MUX1HOT_s_1_4_2((COMP_LOOP_k_9_4_sva_4_0(4)), COMP_LOOP_nor_137_itm,
      COMP_LOOP_nor_134_itm, COMP_LOOP_nor_14_nl, STD_LOGIC_VECTOR'( and_dcpl_283
      & not_tmp_776 & (NOT mux_3577_nl) & COMP_LOOP_or_32_cse));
  nor_558_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(3)) OR (fsm_output(6)) OR
      (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(4)) OR (NOT (fsm_output(10))));
  nor_559_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  mux_3582_nl <= MUX_s_1_2_2(nor_558_nl, nor_559_nl, fsm_output(7));
  nand_452_nl <= NOT((fsm_output(2)) AND mux_3582_nl);
  or_3474_nl <= CONV_SL_1_1(fsm_output(10 DOWNTO 2)/=STD_LOGIC_VECTOR'("011010110"));
  mux_3583_nl <= MUX_s_1_2_2(nand_452_nl, or_3474_nl, fsm_output(1));
  or_3127_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(6))) OR (fsm_output(9))
      OR (fsm_output(8)) OR (NOT (fsm_output(4))) OR (fsm_output(10));
  or_3126_nl <= (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(9)) OR (NOT
      (fsm_output(8))) OR (fsm_output(4)) OR (fsm_output(10));
  mux_3579_nl <= MUX_s_1_2_2(or_3127_nl, or_3126_nl, fsm_output(5));
  or_3125_nl <= (fsm_output(5)) OR (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(9))
      OR (fsm_output(8)) OR (fsm_output(4)) OR (NOT (fsm_output(10)));
  mux_3580_nl <= MUX_s_1_2_2(mux_3579_nl, or_3125_nl, fsm_output(7));
  or_3475_nl <= (fsm_output(2)) OR mux_3580_nl;
  nor_562_nl <= NOT((fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(9)) OR (fsm_output(8))
      OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  nor_563_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(9)))
      OR (NOT (fsm_output(8))) OR (NOT (fsm_output(4))) OR (fsm_output(10)));
  mux_3578_nl <= MUX_s_1_2_2(nor_562_nl, nor_563_nl, fsm_output(5));
  nand_453_nl <= NOT((fsm_output(2)) AND (fsm_output(7)) AND mux_3578_nl);
  mux_3581_nl <= MUX_s_1_2_2(or_3475_nl, nand_453_nl, fsm_output(1));
  mux_3584_nl <= MUX_s_1_2_2(mux_3583_nl, mux_3581_nl, fsm_output(0));
  or_3145_nl <= (NOT (fsm_output(5))) OR (fsm_output(9)) OR not_tmp_51;
  mux_3589_nl <= MUX_s_1_2_2(or_2679_cse, or_3145_nl, fsm_output(3));
  nor_552_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(4))) OR (fsm_output(6)) OR
      mux_3589_nl);
  nor_554_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(8)) OR
      (NOT (fsm_output(10))));
  mux_3588_nl <= MUX_s_1_2_2(nor_670_cse, nor_554_nl, fsm_output(3));
  and_392_nl <= nor_381_cse AND mux_3588_nl;
  mux_3590_nl <= MUX_s_1_2_2(nor_552_nl, and_392_nl, fsm_output(1));
  and_391_nl <= (fsm_output(7)) AND mux_3590_nl;
  nor_555_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(4))) OR (fsm_output(6))
      OR (NOT (fsm_output(3))) OR (fsm_output(5)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(10))));
  or_3136_nl <= (fsm_output(6)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10));
  or_3135_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(5)) OR (fsm_output(9))
      OR not_tmp_51;
  mux_3585_nl <= MUX_s_1_2_2(or_3136_nl, or_3135_nl, fsm_output(4));
  nor_556_nl <= NOT((fsm_output(2)) OR mux_3585_nl);
  mux_3586_nl <= MUX_s_1_2_2(nor_555_nl, nor_556_nl, fsm_output(1));
  nor_557_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT (fsm_output(5))) OR (NOT
      (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(10)));
  mux_3587_nl <= MUX_s_1_2_2(mux_3586_nl, nor_557_nl, fsm_output(7));
  mux_3591_nl <= MUX_s_1_2_2(and_391_nl, mux_3587_nl, fsm_output(0));
  COMP_LOOP_nor_17_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_mux1h_479_nl <= MUX1HOT_s_1_3_2(COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      COMP_LOOP_nor_137_itm, COMP_LOOP_nor_17_nl, STD_LOGIC_VECTOR'( not_tmp_776
      & (NOT mux_3369_itm) & COMP_LOOP_or_32_cse));
  or_3158_nl <= (fsm_output(6)) OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT
      (fsm_output(4))) OR (fsm_output(8)) OR (NOT (fsm_output(9)));
  or_3156_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (fsm_output(4)) OR (NOT (fsm_output(8))) OR (fsm_output(9));
  mux_3596_nl <= MUX_s_1_2_2(or_3158_nl, or_3156_nl, fsm_output(1));
  or_3155_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(9));
  mux_3597_nl <= MUX_s_1_2_2(mux_3596_nl, or_3155_nl, fsm_output(0));
  or_3342_nl <= (fsm_output(3)) OR mux_3597_nl;
  or_3343_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(9));
  nor_548_nl <= NOT((fsm_output(7)) OR (fsm_output(4)) OR (NOT (fsm_output(8))) OR
      (fsm_output(9)));
  and_820_nl <= (fsm_output(7)) AND (fsm_output(4)) AND (NOT (fsm_output(8))) AND
      (fsm_output(9));
  mux_3593_nl <= MUX_s_1_2_2(nor_548_nl, and_820_nl, fsm_output(2));
  nand_419_nl <= NOT((NOT((fsm_output(1)) OR (NOT (fsm_output(6))))) AND mux_3593_nl);
  mux_3594_nl <= MUX_s_1_2_2(or_3343_nl, nand_419_nl, fsm_output(0));
  or_3344_nl <= (fsm_output(1)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(4))) OR (fsm_output(8)) OR (fsm_output(9));
  or_3345_nl <= (NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(7))
      OR (fsm_output(4)) OR (fsm_output(8)) OR (NOT (fsm_output(9)));
  mux_3592_nl <= MUX_s_1_2_2(or_3344_nl, or_3345_nl, fsm_output(0));
  mux_3595_nl <= MUX_s_1_2_2(mux_3594_nl, mux_3592_nl, fsm_output(3));
  mux_3598_nl <= MUX_s_1_2_2(or_3342_nl, mux_3595_nl, fsm_output(5));
  nand_181_nl <= NOT((fsm_output(5)) AND mux_3603_cse);
  nor_541_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR nand_398_cse);
  nor_542_nl <= NOT((fsm_output(2)) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(4))
      OR (NOT (fsm_output(10))));
  mux_3602_nl <= MUX_s_1_2_2(nor_541_nl, nor_542_nl, fsm_output(7));
  nand_180_nl <= NOT(nor_515_cse AND mux_3602_nl);
  mux_3604_nl <= MUX_s_1_2_2(nand_181_nl, nand_180_nl, fsm_output(0));
  nor_538_nl <= NOT((fsm_output(6)) OR mux_3604_nl);
  and_389_nl <= (fsm_output(0)) AND (fsm_output(5)) AND (fsm_output(3)) AND (fsm_output(7))
      AND (fsm_output(2)) AND (fsm_output(9)) AND (fsm_output(8)) AND (fsm_output(4))
      AND (NOT (fsm_output(10)));
  nor_543_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(7)) OR (fsm_output(2)) OR
      (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(4))) OR
      (fsm_output(10)));
  mux_3599_nl <= MUX_s_1_2_2(nor_543_nl, nor_544_cse, fsm_output(5));
  mux_3600_nl <= MUX_s_1_2_2(mux_3599_nl, nor_545_cse, fsm_output(0));
  mux_3601_nl <= MUX_s_1_2_2(and_389_nl, mux_3600_nl, fsm_output(6));
  mux_3605_nl <= MUX_s_1_2_2(nor_538_nl, mux_3601_nl, fsm_output(1));
  mux_3668_nl <= MUX_s_1_2_2(nand_tmp_119, or_tmp_3107, fsm_output(7));
  mux_3667_nl <= MUX_s_1_2_2((NOT nor_tmp_286), (fsm_output(6)), fsm_output(7));
  mux_3669_nl <= MUX_s_1_2_2(mux_3668_nl, mux_3667_nl, fsm_output(5));
  nand_195_nl <= NOT((fsm_output(6)) AND (CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT nor_tmp_6)));
  mux_3665_nl <= MUX_s_1_2_2(nand_195_nl, or_tmp_434, fsm_output(7));
  and_388_nl <= ((fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3)))
      AND (fsm_output(10));
  mux_3664_nl <= MUX_s_1_2_2(and_388_nl, nand_tmp_119, fsm_output(7));
  mux_3666_nl <= MUX_s_1_2_2((NOT mux_3665_nl), mux_3664_nl, fsm_output(5));
  mux_3670_nl <= MUX_s_1_2_2((NOT mux_3669_nl), mux_3666_nl, fsm_output(2));
  mux_3661_nl <= MUX_s_1_2_2(not_tmp_378, mux_tmp_2696, fsm_output(7));
  mux_3659_nl <= MUX_s_1_2_2((NOT or_tmp_2269), or_tmp_9, fsm_output(6));
  and_386_nl <= (fsm_output(6)) AND or_tmp_2483;
  mux_3660_nl <= MUX_s_1_2_2(mux_3659_nl, and_386_nl, fsm_output(7));
  mux_3662_nl <= MUX_s_1_2_2(mux_3661_nl, mux_3660_nl, fsm_output(5));
  or_3182_nl <= (fsm_output(6)) OR (NOT or_tmp_2275);
  and_385_nl <= (fsm_output(6)) AND or_tmp_2220;
  mux_3657_nl <= MUX_s_1_2_2(or_3182_nl, and_385_nl, fsm_output(7));
  mux_3658_nl <= MUX_s_1_2_2(mux_tmp_2290, mux_3657_nl, fsm_output(5));
  mux_3663_nl <= MUX_s_1_2_2(mux_3662_nl, mux_3658_nl, fsm_output(2));
  mux_3671_nl <= MUX_s_1_2_2(mux_3670_nl, mux_3663_nl, fsm_output(8));
  mux_3653_nl <= MUX_s_1_2_2(and_tmp_16, (NOT or_tmp_2479), fsm_output(7));
  mux_3652_nl <= MUX_s_1_2_2(or_15_cse, mux_tmp_893, fsm_output(7));
  mux_3654_nl <= MUX_s_1_2_2(mux_3653_nl, mux_3652_nl, fsm_output(5));
  nand_196_nl <= NOT((fsm_output(6)) AND or_tmp_237);
  mux_3650_nl <= MUX_s_1_2_2(nand_196_nl, or_tmp_2479, fsm_output(7));
  mux_3648_nl <= MUX_s_1_2_2((NOT or_tmp_2253), or_tmp_2248, fsm_output(6));
  mux_3649_nl <= MUX_s_1_2_2(or_tmp_4, mux_3648_nl, fsm_output(7));
  mux_3651_nl <= MUX_s_1_2_2((NOT mux_3650_nl), mux_3649_nl, fsm_output(5));
  mux_3655_nl <= MUX_s_1_2_2(mux_3654_nl, mux_3651_nl, fsm_output(2));
  mux_3644_nl <= MUX_s_1_2_2((NOT nor_tmp_6), or_tmp_2260, fsm_output(6));
  mux_3645_nl <= MUX_s_1_2_2(mux_3644_nl, (fsm_output(6)), fsm_output(7));
  mux_3642_nl <= MUX_s_1_2_2((fsm_output(10)), and_dcpl_240, fsm_output(6));
  mux_3641_nl <= MUX_s_1_2_2(nor_tmp_291, (fsm_output(10)), fsm_output(6));
  mux_3643_nl <= MUX_s_1_2_2((NOT mux_3642_nl), mux_3641_nl, fsm_output(7));
  mux_3646_nl <= MUX_s_1_2_2(mux_3645_nl, mux_3643_nl, fsm_output(5));
  nor_536_nl <= NOT((fsm_output(6)) OR (NOT nor_tmp_9));
  mux_3639_nl <= MUX_s_1_2_2(nor_536_nl, nand_tmp_119, fsm_output(7));
  nand_197_nl <= NOT(((NOT (fsm_output(6))) OR (fsm_output(3))) AND (fsm_output(10)));
  mux_3638_nl <= MUX_s_1_2_2(nand_197_nl, nor_tmp_286, fsm_output(7));
  mux_3640_nl <= MUX_s_1_2_2((NOT mux_3639_nl), mux_3638_nl, fsm_output(5));
  mux_3647_nl <= MUX_s_1_2_2(mux_3646_nl, mux_3640_nl, fsm_output(2));
  mux_3656_nl <= MUX_s_1_2_2(mux_3655_nl, mux_3647_nl, fsm_output(8));
  mux_3672_nl <= MUX_s_1_2_2(mux_3671_nl, mux_3656_nl, fsm_output(4));
  mux_3632_nl <= MUX_s_1_2_2((NOT (fsm_output(10))), nor_tmp_6, fsm_output(6));
  mux_3633_nl <= MUX_s_1_2_2(mux_3632_nl, or_tmp_4, fsm_output(7));
  mux_3631_nl <= MUX_s_1_2_2(or_tmp_434, (fsm_output(10)), fsm_output(7));
  mux_3634_nl <= MUX_s_1_2_2(mux_3633_nl, mux_3631_nl, fsm_output(5));
  mux_3629_nl <= MUX_s_1_2_2(mux_tmp_893, or_tmp_4, fsm_output(7));
  mux_3627_nl <= MUX_s_1_2_2(or_tmp_2479, (fsm_output(10)), fsm_output(7));
  mux_3630_nl <= MUX_s_1_2_2(mux_3629_nl, mux_3627_nl, fsm_output(5));
  mux_3635_nl <= MUX_s_1_2_2(mux_3634_nl, mux_3630_nl, fsm_output(2));
  mux_3624_nl <= MUX_s_1_2_2(or_tmp_14, mux_tmp_2788, fsm_output(7));
  mux_3625_nl <= MUX_s_1_2_2(mux_3624_nl, mux_3_cse, fsm_output(5));
  mux_2589_nl <= MUX_s_1_2_2(or_tmp_14, or_tmp_4, fsm_output(7));
  or_3179_nl <= (NOT (fsm_output(6))) OR (fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(10));
  mux_3622_nl <= MUX_s_1_2_2(or_tmp_4, or_3179_nl, fsm_output(7));
  mux_3623_nl <= MUX_s_1_2_2(mux_2589_nl, mux_3622_nl, fsm_output(5));
  mux_3626_nl <= MUX_s_1_2_2(mux_3625_nl, mux_3623_nl, fsm_output(2));
  mux_3636_nl <= MUX_s_1_2_2(mux_3635_nl, mux_3626_nl, fsm_output(8));
  mux_3617_nl <= MUX_s_1_2_2((NOT (fsm_output(10))), or_tmp_9, fsm_output(6));
  or_3178_nl <= (NOT((fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(3))))
      OR (fsm_output(10));
  mux_3618_nl <= MUX_s_1_2_2(mux_3617_nl, or_3178_nl, fsm_output(7));
  or_3176_nl <= (NOT((fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT
      (fsm_output(3))))) OR (fsm_output(10));
  mux_3616_nl <= MUX_s_1_2_2((fsm_output(6)), or_3176_nl, fsm_output(7));
  mux_3619_nl <= MUX_s_1_2_2(mux_3618_nl, mux_3616_nl, fsm_output(5));
  mux_3614_nl <= MUX_s_1_2_2(or_tmp_3107, (fsm_output(10)), fsm_output(7));
  mux_3611_nl <= MUX_s_1_2_2(or_tmp_2269, or_tmp_2271, fsm_output(6));
  mux_3612_nl <= MUX_s_1_2_2((fsm_output(6)), mux_3611_nl, fsm_output(7));
  mux_3615_nl <= MUX_s_1_2_2(mux_3614_nl, mux_3612_nl, fsm_output(5));
  mux_3620_nl <= MUX_s_1_2_2(mux_3619_nl, mux_3615_nl, fsm_output(2));
  mux_3608_nl <= MUX_s_1_2_2(mux_9_cse, or_tmp_4, fsm_output(7));
  mux_3609_nl <= MUX_s_1_2_2(mux_3608_nl, or_tmp_2263, fsm_output(5));
  mux_3606_nl <= MUX_s_1_2_2(mux_tmp_2790, or_tmp_4, fsm_output(7));
  mux_3607_nl <= MUX_s_1_2_2(mux_3606_nl, or_tmp_2263, fsm_output(5));
  mux_3610_nl <= MUX_s_1_2_2(mux_3609_nl, mux_3607_nl, fsm_output(2));
  mux_3621_nl <= MUX_s_1_2_2(mux_3620_nl, mux_3610_nl, fsm_output(8));
  mux_3637_nl <= MUX_s_1_2_2(mux_3636_nl, mux_3621_nl, fsm_output(4));
  mux_3673_nl <= MUX_s_1_2_2(mux_3672_nl, (NOT mux_3637_nl), fsm_output(9));
  COMP_LOOP_or_28_nl <= and_dcpl_147 OR and_dcpl_217;
  COMP_LOOP_mux1h_480_nl <= MUX1HOT_s_1_6_2(modExp_exp_1_4_1_sva, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      (COMP_LOOP_k_9_4_sva_4_0(0)), (z_out_8_8_7(0)), (z_out_9(6)), (z_out_9(5)),
      STD_LOGIC_VECTOR'( not_tmp_776 & mux_3673_nl & not_tmp_762 & COMP_LOOP_or_28_nl
      & and_dcpl_182 & and_dcpl_247));
  or_3297_nl <= (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(10));
  nand_250_nl <= NOT((fsm_output(0)) AND (fsm_output(7)) AND (fsm_output(9)) AND
      (fsm_output(10)));
  mux_2493_nl <= MUX_s_1_2_2(or_3297_nl, nand_250_nl, fsm_output(1));
  mux_2494_nl <= MUX_s_1_2_2(mux_2493_nl, nand_375_cse, or_495_cse);
  mux_2495_nl <= MUX_s_1_2_2(mux_2494_nl, nand_376_cse, fsm_output(8));
  nor_1453_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))))
      OR (fsm_output(4)));
  mux_3890_nl <= MUX_s_1_2_2(nor_1453_nl, mux_tmp_3878, fsm_output(9));
  mux_3891_nl <= MUX_s_1_2_2(mux_3890_nl, mux_tmp_3834, fsm_output(3));
  mux_3889_nl <= MUX_s_1_2_2(not_tmp_1021, mux_tmp_3828, fsm_output(3));
  mux_3892_nl <= MUX_s_1_2_2((NOT mux_3891_nl), mux_3889_nl, fsm_output(10));
  and_1258_nl <= ((fsm_output(9)) OR (fsm_output(1)) OR (NOT (fsm_output(0))) OR
      (fsm_output(2))) AND (fsm_output(4));
  mux_3886_nl <= MUX_s_1_2_2((fsm_output(4)), or_tmp_3303, fsm_output(9));
  mux_3887_nl <= MUX_s_1_2_2(and_1258_nl, mux_3886_nl, fsm_output(3));
  or_3508_nl <= (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(2)) OR (fsm_output(4));
  mux_3888_nl <= MUX_s_1_2_2(mux_3887_nl, or_3508_nl, fsm_output(10));
  mux_3893_nl <= MUX_s_1_2_2(mux_3892_nl, mux_3888_nl, fsm_output(5));
  and_1259_nl <= (fsm_output(3)) AND (fsm_output(9)) AND (fsm_output(1)) AND (fsm_output(0))
      AND (fsm_output(2)) AND (fsm_output(4));
  mux_3883_nl <= MUX_s_1_2_2((fsm_output(9)), or_2747_cse, fsm_output(3));
  mux_3884_nl <= MUX_s_1_2_2(and_1259_nl, mux_3883_nl, fsm_output(10));
  and_1260_nl <= ((fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(2)))
      AND (fsm_output(4));
  mux_3881_nl <= MUX_s_1_2_2(mux_tmp_3853, and_1260_nl, fsm_output(3));
  or_3506_nl <= (fsm_output(9)) OR mux_tmp_3878;
  mux_3880_nl <= MUX_s_1_2_2(or_tmp, or_3506_nl, fsm_output(3));
  mux_3882_nl <= MUX_s_1_2_2((NOT mux_3881_nl), mux_3880_nl, fsm_output(10));
  mux_3885_nl <= MUX_s_1_2_2(mux_3884_nl, mux_3882_nl, fsm_output(5));
  mux_3894_nl <= MUX_s_1_2_2((NOT mux_3893_nl), mux_3885_nl, fsm_output(8));
  or_3505_nl <= (fsm_output(3)) OR (fsm_output(9));
  mux_3875_nl <= MUX_s_1_2_2(mux_tmp_3861, (fsm_output(4)), or_3505_nl);
  or_3504_nl <= (fsm_output(9)) OR (NOT((fsm_output(1)) OR (fsm_output(0)) OR (fsm_output(2))
      OR (fsm_output(4))));
  mux_3874_nl <= MUX_s_1_2_2(or_tmp, or_3504_nl, fsm_output(3));
  mux_3876_nl <= MUX_s_1_2_2((NOT mux_3875_nl), mux_3874_nl, fsm_output(10));
  and_1256_nl <= (fsm_output(3)) AND (fsm_output(9)) AND nor_tmp_540;
  or_3502_nl <= (fsm_output(9)) OR nor_tmp_539;
  mux_3872_nl <= MUX_s_1_2_2(or_3502_nl, or_2747_cse, fsm_output(3));
  mux_3873_nl <= MUX_s_1_2_2(and_1256_nl, mux_3872_nl, fsm_output(10));
  mux_3877_nl <= MUX_s_1_2_2(mux_3876_nl, mux_3873_nl, fsm_output(5));
  mux_3867_nl <= MUX_s_1_2_2(not_tmp_1007, mux_tmp_3818, and_573_cse);
  mux_3868_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), mux_3867_nl, fsm_output(9));
  mux_3865_nl <= MUX_s_1_2_2(not_tmp_1007, mux_tmp_3846, fsm_output(1));
  mux_3866_nl <= MUX_s_1_2_2(mux_3865_nl, (fsm_output(4)), fsm_output(9));
  mux_3869_nl <= MUX_s_1_2_2(mux_3868_nl, mux_3866_nl, fsm_output(3));
  mux_3870_nl <= MUX_s_1_2_2((NOT mux_3869_nl), or_tmp, fsm_output(10));
  mux_3863_nl <= MUX_s_1_2_2((fsm_output(4)), (NOT mux_tmp_3861), and_1262_cse);
  or_3500_nl <= (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(4));
  mux_3861_nl <= MUX_s_1_2_2(or_3500_nl, or_tmp, fsm_output(3));
  mux_3864_nl <= MUX_s_1_2_2(mux_3863_nl, mux_3861_nl, fsm_output(10));
  mux_3871_nl <= MUX_s_1_2_2(mux_3870_nl, mux_3864_nl, fsm_output(5));
  mux_3878_nl <= MUX_s_1_2_2(mux_3877_nl, mux_3871_nl, fsm_output(8));
  mux_3895_nl <= MUX_s_1_2_2(mux_3894_nl, mux_3878_nl, fsm_output(7));
  and_1255_nl <= (fsm_output(9)) AND nor_tmp_536;
  mux_3856_nl <= MUX_s_1_2_2(and_1255_nl, nor_tmp_535, fsm_output(3));
  mux_3855_nl <= MUX_s_1_2_2(not_tmp_1021, mux_tmp_3853, fsm_output(3));
  mux_3857_nl <= MUX_s_1_2_2(mux_3856_nl, (NOT mux_3855_nl), fsm_output(10));
  nor_1456_nl <= NOT(and_565_cse OR (fsm_output(4)));
  mux_3851_nl <= MUX_s_1_2_2(nor_1456_nl, nor_tmp_540, fsm_output(9));
  mux_3852_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), mux_3851_nl, fsm_output(3));
  and_1264_nl <= ((fsm_output(0)) OR (fsm_output(2))) AND (fsm_output(4));
  mux_3848_nl <= MUX_s_1_2_2(mux_tmp_3846, and_1264_nl, fsm_output(1));
  mux_3849_nl <= MUX_s_1_2_2(mux_3848_nl, (fsm_output(4)), fsm_output(9));
  mux_3850_nl <= MUX_s_1_2_2(mux_3849_nl, or_tmp_3304, fsm_output(3));
  mux_3853_nl <= MUX_s_1_2_2(mux_3852_nl, mux_3850_nl, fsm_output(10));
  mux_3858_nl <= MUX_s_1_2_2(mux_3857_nl, mux_3853_nl, fsm_output(5));
  mux_3843_nl <= MUX_s_1_2_2(or_tmp_3303, (NOT nor_tmp_540), fsm_output(9));
  mux_3844_nl <= MUX_s_1_2_2(or_tmp_3304, mux_3843_nl, fsm_output(3));
  or_3493_nl <= (fsm_output(9)) OR (NOT nor_tmp_539);
  mux_3842_nl <= MUX_s_1_2_2(or_3493_nl, or_tmp, fsm_output(3));
  mux_3845_nl <= MUX_s_1_2_2(mux_3844_nl, mux_3842_nl, fsm_output(10));
  nor_1457_nl <= NOT((fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR (fsm_output(4)));
  or_3490_nl <= (fsm_output(9)) OR nor_tmp_536;
  mux_3840_nl <= MUX_s_1_2_2((fsm_output(9)), or_3490_nl, fsm_output(3));
  mux_3841_nl <= MUX_s_1_2_2(nor_1457_nl, mux_3840_nl, fsm_output(10));
  mux_3846_nl <= MUX_s_1_2_2(mux_3845_nl, mux_3841_nl, fsm_output(5));
  mux_3859_nl <= MUX_s_1_2_2(mux_3858_nl, mux_3846_nl, fsm_output(8));
  nor_1458_nl <= NOT(((fsm_output(0)) AND (fsm_output(2))) OR (fsm_output(4)));
  mux_3833_nl <= MUX_s_1_2_2(nor_1458_nl, mux_tmp_3819, fsm_output(1));
  mux_3834_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), mux_3833_nl, fsm_output(9));
  mux_3836_nl <= MUX_s_1_2_2((NOT mux_tmp_3834), mux_3834_nl, fsm_output(3));
  mux_3832_nl <= MUX_s_1_2_2(or_tmp_3293, or_2747_cse, fsm_output(3));
  mux_3837_nl <= MUX_s_1_2_2(mux_3836_nl, mux_3832_nl, fsm_output(10));
  mux_3830_nl <= MUX_s_1_2_2(mux_tmp_3828, nor_tmp_535, fsm_output(3));
  mux_3828_nl <= MUX_s_1_2_2(or_tmp, or_tmp_3293, fsm_output(3));
  mux_3831_nl <= MUX_s_1_2_2((NOT mux_3830_nl), mux_3828_nl, fsm_output(10));
  mux_3838_nl <= MUX_s_1_2_2(mux_3837_nl, mux_3831_nl, fsm_output(5));
  nor_1459_nl <= NOT((fsm_output(3)) OR (fsm_output(9)) OR or_tmp_3291);
  mux_3826_nl <= MUX_s_1_2_2(nor_1459_nl, (fsm_output(9)), fsm_output(10));
  mux_3824_nl <= MUX_s_1_2_2((fsm_output(4)), (NOT mux_tmp_3822), and_1262_cse);
  mux_3821_nl <= MUX_s_1_2_2(mux_tmp_3819, nor_tmp, fsm_output(1));
  or_3480_nl <= (fsm_output(9)) OR (NOT mux_3821_nl);
  mux_3822_nl <= MUX_s_1_2_2(or_3480_nl, or_tmp, fsm_output(3));
  mux_3825_nl <= MUX_s_1_2_2(mux_3824_nl, mux_3822_nl, fsm_output(10));
  mux_3827_nl <= MUX_s_1_2_2(mux_3826_nl, mux_3825_nl, fsm_output(5));
  mux_3839_nl <= MUX_s_1_2_2(mux_3838_nl, mux_3827_nl, fsm_output(8));
  mux_3860_nl <= MUX_s_1_2_2(mux_3859_nl, mux_3839_nl, fsm_output(7));
  mux_3896_nl <= MUX_s_1_2_2(mux_3895_nl, mux_3860_nl, fsm_output(6));
  or_3579_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(1))) OR (NOT COMP_LOOP_nor_11_itm)
      OR (fsm_output(8)) OR (fsm_output(10)) OR not_tmp_1034;
  mux_3943_nl <= MUX_s_1_2_2(nand_201_cse, or_tmp_3327, fsm_output(8));
  nand_463_nl <= NOT((fsm_output(1)) AND (NOT mux_3943_nl));
  mux_3944_nl <= MUX_s_1_2_2(or_tmp_3343, nand_463_nl, fsm_output(6));
  mux_3945_nl <= MUX_s_1_2_2(or_3579_nl, mux_3944_nl, fsm_output(3));
  mux_3941_nl <= MUX_s_1_2_2(or_tmp_3369, mux_tmp_3902, fsm_output(1));
  or_3577_nl <= (fsm_output(6)) OR mux_3941_nl;
  mux_3942_nl <= MUX_s_1_2_2(or_3577_nl, nand_tmp, fsm_output(3));
  mux_3946_nl <= MUX_s_1_2_2(mux_3945_nl, mux_3942_nl, fsm_output(5));
  nor_1448_nl <= NOT((NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8)) OR (NOT (fsm_output(10)))
      OR (NOT (fsm_output(9))) OR (fsm_output(4)));
  nor_1449_nl <= NOT((NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8)) OR (fsm_output(10))
      OR (fsm_output(9)) OR (fsm_output(4)));
  mux_3938_nl <= MUX_s_1_2_2(nor_1448_nl, nor_1449_nl, fsm_output(1));
  nand_462_nl <= NOT((fsm_output(6)) AND mux_3938_nl);
  or_3574_nl <= (fsm_output(1)) OR (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(8)))
      OR (fsm_output(10)) OR not_tmp_1034;
  mux_3939_nl <= MUX_s_1_2_2(nand_462_nl, or_3574_nl, fsm_output(3));
  or_3572_nl <= (fsm_output(3)) OR (fsm_output(6)) OR nor_1450_cse OR (fsm_output(8))
      OR (NOT (fsm_output(10))) OR (fsm_output(9)) OR (fsm_output(4));
  mux_3940_nl <= MUX_s_1_2_2(mux_3939_nl, or_3572_nl, fsm_output(5));
  mux_3947_nl <= MUX_s_1_2_2(mux_3946_nl, mux_3940_nl, fsm_output(2));
  or_3568_nl <= (fsm_output(6)) OR mux_tmp_3898;
  mux_3935_nl <= MUX_s_1_2_2(or_3568_nl, or_tmp_3320, fsm_output(3));
  or_3567_nl <= (fsm_output(1)) OR (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8))
      OR (NOT (fsm_output(10))) OR (fsm_output(9)) OR (NOT (fsm_output(4)));
  or_3565_nl <= (fsm_output(6)) OR nor_1450_cse OR (NOT (fsm_output(8))) OR (NOT
      (fsm_output(10))) OR (fsm_output(9)) OR (NOT (fsm_output(4)));
  mux_3934_nl <= MUX_s_1_2_2(or_3567_nl, or_3565_nl, fsm_output(3));
  mux_3936_nl <= MUX_s_1_2_2(mux_3935_nl, mux_3934_nl, fsm_output(5));
  mux_3931_nl <= MUX_s_1_2_2(or_tmp_3369, mux_tmp_3915, fsm_output(1));
  nand_461_nl <= NOT((fsm_output(6)) AND (NOT mux_3931_nl));
  or_3559_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(8)))
      OR (fsm_output(10)) OR (fsm_output(9)) OR (NOT (fsm_output(4)));
  mux_3932_nl <= MUX_s_1_2_2(nand_461_nl, or_3559_nl, fsm_output(3));
  nand_465_nl <= NOT((fsm_output(6)) AND (fsm_output(1)) AND COMP_LOOP_nor_11_itm
      AND (fsm_output(8)) AND (NOT (fsm_output(10))) AND (fsm_output(9)) AND (NOT
      (fsm_output(4))));
  or_3556_nl <= (NOT (fsm_output(1))) OR (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8))
      OR (fsm_output(10)) OR (fsm_output(9)) OR (NOT (fsm_output(4)));
  mux_3928_nl <= MUX_s_1_2_2(mux_tmp_3902, mux_tmp_3906, fsm_output(1));
  mux_3929_nl <= MUX_s_1_2_2(or_3556_nl, mux_3928_nl, fsm_output(6));
  mux_3930_nl <= MUX_s_1_2_2(nand_465_nl, mux_3929_nl, fsm_output(3));
  mux_3933_nl <= MUX_s_1_2_2(mux_3932_nl, mux_3930_nl, fsm_output(5));
  mux_3937_nl <= MUX_s_1_2_2(mux_3936_nl, mux_3933_nl, fsm_output(2));
  mux_3948_nl <= MUX_s_1_2_2(mux_3947_nl, mux_3937_nl, fsm_output(7));
  or_3554_nl <= (fsm_output(8)) OR (fsm_output(10)) OR (fsm_output(9)) OR (fsm_output(4));
  mux_3922_nl <= MUX_s_1_2_2(or_3554_nl, or_tmp_3332, fsm_output(1));
  nand_471_nl <= NOT((fsm_output(1)) AND (fsm_output(8)) AND (fsm_output(10)) AND
      (NOT (fsm_output(9))) AND (fsm_output(4)));
  mux_3923_nl <= MUX_s_1_2_2(mux_3922_nl, nand_471_nl, fsm_output(6));
  or_3551_nl <= (fsm_output(1)) OR (fsm_output(8)) OR (fsm_output(10)) OR (fsm_output(9))
      OR (fsm_output(4));
  or_3550_nl <= (NOT (fsm_output(1))) OR (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8))
      OR (NOT (fsm_output(10))) OR (fsm_output(9)) OR (fsm_output(4));
  mux_3921_nl <= MUX_s_1_2_2(or_3551_nl, or_3550_nl, fsm_output(6));
  mux_3924_nl <= MUX_s_1_2_2(mux_3923_nl, mux_3921_nl, fsm_output(3));
  mux_3918_nl <= MUX_s_1_2_2(or_tmp_195, or_tmp_182, fsm_output(8));
  nand_460_nl <= NOT((fsm_output(1)) AND COMP_LOOP_nor_11_itm AND (NOT mux_3918_nl));
  or_3548_nl <= (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(8))) OR (fsm_output(10))
      OR (fsm_output(9)) OR (fsm_output(4));
  mux_3917_nl <= MUX_s_1_2_2(mux_tmp_3915, or_3548_nl, fsm_output(1));
  mux_3919_nl <= MUX_s_1_2_2(nand_460_nl, mux_3917_nl, fsm_output(6));
  or_3546_nl <= (NOT (fsm_output(8))) OR (fsm_output(10)) OR (fsm_output(9)) OR (NOT
      (fsm_output(4)));
  or_3544_nl <= (fsm_output(10)) OR (NOT (fsm_output(9))) OR (fsm_output(4));
  mux_3914_nl <= MUX_s_1_2_2(or_3544_nl, or_2415_cse, fsm_output(8));
  mux_3915_nl <= MUX_s_1_2_2(or_3546_nl, mux_3914_nl, fsm_output(1));
  or_3547_nl <= (fsm_output(6)) OR mux_3915_nl;
  mux_3920_nl <= MUX_s_1_2_2(mux_3919_nl, or_3547_nl, fsm_output(3));
  mux_3925_nl <= MUX_s_1_2_2(mux_3924_nl, mux_3920_nl, fsm_output(5));
  or_3542_nl <= (fsm_output(1)) OR (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(8)))
      OR (NOT (fsm_output(10))) OR (fsm_output(9)) OR (NOT (fsm_output(4)));
  or_3540_nl <= (fsm_output(6)) OR nor_1450_cse OR (fsm_output(8)) OR nand_201_cse;
  mux_3912_nl <= MUX_s_1_2_2(or_3542_nl, or_3540_nl, fsm_output(3));
  or_3536_nl <= (fsm_output(1)) OR (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8))
      OR (fsm_output(10)) OR (NOT (fsm_output(9))) OR (fsm_output(4));
  mux_3911_nl <= MUX_s_1_2_2(or_3536_nl, or_tmp_3343, fsm_output(6));
  nand_459_nl <= NOT((fsm_output(3)) AND (NOT mux_3911_nl));
  mux_3913_nl <= MUX_s_1_2_2(mux_3912_nl, nand_459_nl, fsm_output(5));
  mux_3926_nl <= MUX_s_1_2_2(mux_3925_nl, mux_3913_nl, fsm_output(2));
  or_3533_nl <= (fsm_output(1)) OR (NOT COMP_LOOP_nor_11_itm) OR (NOT (fsm_output(8)))
      OR (fsm_output(10)) OR (NOT (fsm_output(9))) OR (fsm_output(4));
  or_3527_nl <= (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8)) OR (NOT (fsm_output(10)))
      OR (fsm_output(9)) OR (fsm_output(4));
  mux_3908_nl <= MUX_s_1_2_2(mux_tmp_3906, or_3527_nl, fsm_output(1));
  or_3532_nl <= (fsm_output(6)) OR mux_3908_nl;
  mux_3909_nl <= MUX_s_1_2_2(or_3533_nl, or_3532_nl, fsm_output(3));
  or_3534_nl <= (fsm_output(5)) OR mux_3909_nl;
  or_3589_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR mux_tmp_3902;
  mux_3904_nl <= MUX_s_1_2_2(or_3589_nl, nand_tmp, fsm_output(3));
  or_3521_nl <= (NOT (fsm_output(1))) OR (NOT COMP_LOOP_nor_11_itm) OR (fsm_output(8))
      OR (fsm_output(10)) OR not_tmp_1034;
  mux_3900_nl <= MUX_s_1_2_2(or_3521_nl, mux_tmp_3898, fsm_output(6));
  or_3514_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(8))) OR (fsm_output(10))
      OR not_tmp_1034;
  mux_3897_nl <= MUX_s_1_2_2(or_3514_nl, or_tmp_3320, fsm_output(6));
  mux_3901_nl <= MUX_s_1_2_2(mux_3900_nl, mux_3897_nl, fsm_output(3));
  mux_3905_nl <= MUX_s_1_2_2(mux_3904_nl, mux_3901_nl, fsm_output(5));
  mux_3910_nl <= MUX_s_1_2_2(or_3534_nl, mux_3905_nl, fsm_output(2));
  mux_3927_nl <= MUX_s_1_2_2(mux_3926_nl, mux_3910_nl, fsm_output(7));
  mux_3949_nl <= MUX_s_1_2_2(mux_3948_nl, mux_3927_nl, fsm_output(0));
  or_2515_nl <= (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(0))) OR (fsm_output(1))
      OR (NOT (fsm_output(3))) OR (fsm_output(10));
  or_2514_nl <= (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(10));
  mux_2648_nl <= MUX_s_1_2_2(or_2515_nl, or_2514_nl, fsm_output(4));
  or_2513_nl <= (fsm_output(4)) OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(0))
      OR (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(10)));
  mux_2649_nl <= MUX_s_1_2_2(mux_2648_nl, or_2513_nl, fsm_output(9));
  or_3477_nl <= mux_2649_nl OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(8));
  or_3584_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("110"));
  or_3583_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("001"));
  mux_3950_nl <= MUX_s_1_2_2(or_3584_nl, or_3583_nl, fsm_output(0));
  or_3585_nl <= (fsm_output(1)) OR (fsm_output(9)) OR (fsm_output(10)) OR mux_3950_nl;
  or_3581_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(10)))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(5));
  mux_3951_nl <= MUX_s_1_2_2(or_3585_nl, or_3581_nl, fsm_output(7));
  or_3587_nl <= (fsm_output(6)) OR mux_3951_nl;
  or_3588_nl <= (NOT (fsm_output(6))) OR (fsm_output(7)) OR (fsm_output(1)) OR (NOT
      (fsm_output(9))) OR (NOT (fsm_output(10))) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (fsm_output(4)) OR (fsm_output(5));
  mux_3952_nl <= MUX_s_1_2_2(or_3587_nl, or_3588_nl, fsm_output(2));
  nor_725_nl <= NOT((fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(10)));
  mux_2670_nl <= MUX_s_1_2_2(nor_725_nl, mux_tmp_2650, and_573_cse);
  mux_2669_nl <= MUX_s_1_2_2(mux_tmp_2650, and_815_cse, fsm_output(1));
  mux_2671_nl <= MUX_s_1_2_2(mux_2670_nl, mux_2669_nl, fsm_output(3));
  mux_2668_nl <= MUX_s_1_2_2(mux_tmp_2650, and_815_cse, fsm_output(3));
  mux_2672_nl <= MUX_s_1_2_2(mux_2671_nl, mux_2668_nl, fsm_output(2));
  nand_244_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101")));
  mux_2667_nl <= MUX_s_1_2_2(mux_tmp_2650, and_815_cse, nand_244_nl);
  mux_2673_nl <= MUX_s_1_2_2(mux_2672_nl, mux_2667_nl, fsm_output(4));
  or_4_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"));
  mux_2674_nl <= MUX_s_1_2_2(mux_2673_nl, and_815_cse, or_4_nl);
  mux_2675_nl <= MUX_s_1_2_2(mux_2674_nl, and_816_cse, fsm_output(8));
  COMP_LOOP_or_8_nl <= (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_339_m1c);
  COMP_LOOP_or_9_nl <= (COMP_LOOP_COMP_LOOP_and_305_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_339_m1c);
  COMP_LOOP_or_10_nl <= (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_339_m1c);
  COMP_LOOP_or_11_nl <= (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_339_m1c);
  COMP_LOOP_or_12_nl <= (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_339_m1c);
  COMP_LOOP_or_13_nl <= (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_339_m1c);
  COMP_LOOP_or_14_nl <= (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_339_m1c);
  COMP_LOOP_or_15_nl <= (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_339_m1c);
  COMP_LOOP_or_16_nl <= (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_339_m1c);
  COMP_LOOP_or_17_nl <= (COMP_LOOP_COMP_LOOP_and_8_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_339_m1c);
  COMP_LOOP_or_18_nl <= (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_339_m1c);
  COMP_LOOP_or_19_nl <= (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_339_m1c);
  COMP_LOOP_or_20_nl <= (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_339_m1c);
  COMP_LOOP_or_21_nl <= (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_339_m1c);
  COMP_LOOP_or_22_nl <= (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_339_m1c);
  COMP_LOOP_or_23_nl <= (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_283) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_305_m1c) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_307_m1c) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_309_m1c) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_312_m1c) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_315_m1c) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_317_m1c) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_320_m1c) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_322_m1c) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_324_m1c) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_327_m1c) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_329_m1c) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_331_m1c) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_334_m1c) OR (COMP_LOOP_COMP_LOOP_and_305_itm AND and_336_m1c) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_339_m1c);
  nor_716_nl <= NOT((fsm_output(6)) OR and_dcpl_124);
  mux_2736_nl <= MUX_s_1_2_2(nor_716_nl, mux_tmp_2687, fsm_output(7));
  mux_2734_nl <= MUX_s_1_2_2(and_dcpl_109, nor_tmp_9, fsm_output(6));
  mux_2735_nl <= MUX_s_1_2_2(mux_2734_nl, (fsm_output(6)), fsm_output(7));
  mux_2737_nl <= MUX_s_1_2_2(mux_2736_nl, mux_2735_nl, fsm_output(5));
  or_3268_nl <= (fsm_output(6)) OR and_dcpl_123;
  mux_2731_nl <= MUX_s_1_2_2(nor_tmp_6, (NOT nor_tmp_288), fsm_output(6));
  mux_2732_nl <= MUX_s_1_2_2(or_3268_nl, mux_2731_nl, fsm_output(7));
  mux_2729_nl <= MUX_s_1_2_2(or_tmp_2483, (NOT or_tmp_2233), fsm_output(6));
  mux_2730_nl <= MUX_s_1_2_2(mux_2729_nl, nand_tmp_119, fsm_output(7));
  mux_2733_nl <= MUX_s_1_2_2(mux_2732_nl, mux_2730_nl, fsm_output(5));
  mux_2738_nl <= MUX_s_1_2_2((NOT mux_2737_nl), mux_2733_nl, fsm_output(2));
  mux_55_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), or_tmp_3, fsm_output(7));
  mux_2724_nl <= MUX_s_1_2_2((NOT nor_tmp_300), or_tmp_9, fsm_output(6));
  mux_2725_nl <= MUX_s_1_2_2(mux_2724_nl, (fsm_output(6)), fsm_output(7));
  mux_2727_nl <= MUX_s_1_2_2(mux_55_nl, mux_2725_nl, fsm_output(5));
  mux_2722_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), nand_tmp_93, fsm_output(7));
  mux_50_nl <= MUX_s_1_2_2(or_36_cse, (fsm_output(6)), fsm_output(7));
  mux_2723_nl <= MUX_s_1_2_2(mux_2722_nl, mux_50_nl, fsm_output(5));
  mux_2728_nl <= MUX_s_1_2_2(mux_2727_nl, mux_2723_nl, fsm_output(2));
  mux_2739_nl <= MUX_s_1_2_2(mux_2738_nl, mux_2728_nl, fsm_output(8));
  mux_2717_nl <= MUX_s_1_2_2(and_dcpl_243, mux_tmp_2696, fsm_output(7));
  mux_2718_nl <= MUX_s_1_2_2((NOT mux_2717_nl), mux_tmp_2701, fsm_output(5));
  mux_2715_nl <= MUX_s_1_2_2(and_dcpl_243, or_tmp_2479, fsm_output(7));
  mux_2716_nl <= MUX_s_1_2_2((NOT mux_2715_nl), mux_tmp_2698, fsm_output(5));
  mux_2719_nl <= MUX_s_1_2_2(mux_2718_nl, mux_2716_nl, fsm_output(2));
  nand_118_nl <= NOT((fsm_output(6)) AND (NOT nor_tmp_6));
  mux_2712_nl <= MUX_s_1_2_2(nand_118_nl, or_tmp_434, fsm_output(7));
  or_3269_nl <= (fsm_output(6)) OR (NOT or_tmp_2248);
  mux_2710_nl <= MUX_s_1_2_2(nor_tmp_291, (NOT nor_tmp_6), fsm_output(6));
  mux_2711_nl <= MUX_s_1_2_2(or_3269_nl, mux_2710_nl, fsm_output(7));
  mux_2713_nl <= MUX_s_1_2_2(mux_2712_nl, mux_2711_nl, fsm_output(5));
  or_2540_nl <= (fsm_output(6)) OR (NOT or_tmp_2253);
  mux_2708_nl <= MUX_s_1_2_2(or_tmp_4, or_2540_nl, fsm_output(7));
  mux_2706_nl <= MUX_s_1_2_2(nor_tmp_6, (NOT nor_tmp_9), fsm_output(6));
  mux_2707_nl <= MUX_s_1_2_2(or_tmp_2479, mux_2706_nl, fsm_output(7));
  mux_2709_nl <= MUX_s_1_2_2(mux_2708_nl, mux_2707_nl, fsm_output(5));
  mux_2714_nl <= MUX_s_1_2_2(mux_2713_nl, mux_2709_nl, fsm_output(2));
  mux_2720_nl <= MUX_s_1_2_2(mux_2719_nl, mux_2714_nl, fsm_output(8));
  mux_2740_nl <= MUX_s_1_2_2(mux_2739_nl, mux_2720_nl, fsm_output(4));
  mux_29_nl <= MUX_s_1_2_2(mux_28_cse, or_tmp_14, fsm_output(7));
  mux_2702_nl <= MUX_s_1_2_2(mux_tmp_2701, mux_29_nl, fsm_output(5));
  mux_2697_nl <= MUX_s_1_2_2(mux_tmp_2696, or_tmp_14, fsm_output(7));
  mux_2699_nl <= MUX_s_1_2_2(mux_tmp_2698, mux_2697_nl, fsm_output(5));
  mux_2703_nl <= MUX_s_1_2_2(mux_2702_nl, mux_2699_nl, fsm_output(2));
  or_25_nl <= (NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"))))
      OR (fsm_output(10));
  or_24_nl <= nor_223_cse OR (fsm_output(10));
  mux_22_nl <= MUX_s_1_2_2(or_25_nl, or_24_nl, fsm_output(5));
  mux_2704_nl <= MUX_s_1_2_2(mux_2703_nl, mux_22_nl, fsm_output(8));
  nand_116_nl <= NOT((fsm_output(6)) AND (NOT and_dcpl_240));
  mux_2691_nl <= MUX_s_1_2_2(nand_116_nl, or_tmp_2474, fsm_output(7));
  mux_17_nl <= MUX_s_1_2_2((fsm_output(6)), or_tmp_8, fsm_output(7));
  mux_2692_nl <= MUX_s_1_2_2(mux_2691_nl, mux_17_nl, fsm_output(5));
  mux_2688_nl <= MUX_s_1_2_2(mux_tmp_2687, or_tmp_14, fsm_output(7));
  or_18_nl <= (NOT((NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1))))
      OR (fsm_output(10));
  mux_13_nl <= MUX_s_1_2_2((fsm_output(6)), or_18_nl, fsm_output(7));
  mux_2689_nl <= MUX_s_1_2_2(mux_2688_nl, mux_13_nl, fsm_output(5));
  mux_2693_nl <= MUX_s_1_2_2(mux_2692_nl, mux_2689_nl, fsm_output(2));
  mux_10_nl <= MUX_s_1_2_2(mux_9_cse, or_15_cse, fsm_output(7));
  mux_8_nl <= MUX_s_1_2_2(mux_7_cse, or_tmp_4, fsm_output(7));
  mux_11_nl <= MUX_s_1_2_2(mux_10_nl, mux_8_nl, fsm_output(5));
  mux_2677_nl <= MUX_s_1_2_2(or_tmp_2230, (fsm_output(10)), fsm_output(6));
  mux_2678_nl <= MUX_s_1_2_2(or_tmp_8, mux_2677_nl, fsm_output(7));
  mux_2679_nl <= MUX_s_1_2_2(mux_2678_nl, mux_3_cse, fsm_output(5));
  mux_2685_nl <= MUX_s_1_2_2(mux_11_nl, mux_2679_nl, fsm_output(2));
  mux_2694_nl <= MUX_s_1_2_2(mux_2693_nl, mux_2685_nl, fsm_output(8));
  mux_2705_nl <= MUX_s_1_2_2(mux_2704_nl, mux_2694_nl, fsm_output(4));
  and_340_nl <= and_dcpl_191 AND and_dcpl_98;
  COMP_LOOP_or_30_nl <= ((NOT (modulo_result_rem_cmp_z(63))) AND and_345_m1c) OR
      (not_tmp_634 AND (NOT (modulo_result_rem_cmp_z(63))));
  COMP_LOOP_or_31_nl <= ((modulo_result_rem_cmp_z(63)) AND and_345_m1c) OR (not_tmp_634
      AND (modulo_result_rem_cmp_z(63)));
  COMP_LOOP_and_277_nl <= COMP_LOOP_COMP_LOOP_nor_1_itm AND mux_2770_m1c;
  COMP_LOOP_COMP_LOOP_and_932_nl <= (COMP_LOOP_acc_10_cse_12_1_1_sva(0)) AND COMP_LOOP_nor_11_itm
      AND mux_2770_m1c;
  COMP_LOOP_COMP_LOOP_and_934_nl <= (COMP_LOOP_acc_10_cse_12_1_1_sva(1)) AND COMP_LOOP_nor_12_itm
      AND mux_2770_m1c;
  COMP_LOOP_and_1_nl <= COMP_LOOP_COMP_LOOP_and_137_itm AND mux_2770_m1c;
  COMP_LOOP_COMP_LOOP_and_936_nl <= (COMP_LOOP_acc_10_cse_12_1_1_sva(2)) AND COMP_LOOP_nor_134_itm
      AND mux_2770_m1c;
  COMP_LOOP_and_2_nl <= COMP_LOOP_COMP_LOOP_and_139_itm AND mux_2770_m1c;
  COMP_LOOP_and_3_nl <= COMP_LOOP_COMP_LOOP_and_140_itm AND mux_2770_m1c;
  COMP_LOOP_and_4_nl <= COMP_LOOP_COMP_LOOP_and_141_itm AND mux_2770_m1c;
  COMP_LOOP_COMP_LOOP_and_930_nl <= (COMP_LOOP_acc_10_cse_12_1_1_sva(3)) AND COMP_LOOP_nor_137_itm
      AND mux_2770_m1c;
  COMP_LOOP_and_5_nl <= COMP_LOOP_COMP_LOOP_and_143_itm AND mux_2770_m1c;
  COMP_LOOP_and_6_nl <= COMP_LOOP_COMP_LOOP_and_144_itm AND mux_2770_m1c;
  COMP_LOOP_and_7_nl <= COMP_LOOP_COMP_LOOP_and_145_itm AND mux_2770_m1c;
  COMP_LOOP_and_8_nl <= COMP_LOOP_COMP_LOOP_and_146_itm AND mux_2770_m1c;
  COMP_LOOP_and_9_nl <= COMP_LOOP_COMP_LOOP_and_147_itm AND mux_2770_m1c;
  COMP_LOOP_and_10_nl <= COMP_LOOP_COMP_LOOP_and_148_itm AND mux_2770_m1c;
  COMP_LOOP_and_11_nl <= COMP_LOOP_COMP_LOOP_and_149_itm AND mux_2770_m1c;
  nor_1265_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(7)))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(5))
      OR (fsm_output(10)));
  nor_1266_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(8))) OR (fsm_output(7))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(5))
      OR (NOT (fsm_output(10))));
  mux_112_nl <= MUX_s_1_2_2(nor_1265_nl, nor_1266_nl, fsm_output(4));
  or_113_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(0))) OR (fsm_output(3))
      OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  nand_395_nl <= NOT((fsm_output(7)) AND (fsm_output(0)) AND (fsm_output(3)) AND
      (fsm_output(9)) AND (fsm_output(5)) AND (NOT (fsm_output(10))));
  mux_110_nl <= MUX_s_1_2_2(or_113_nl, nand_395_nl, fsm_output(8));
  nor_1267_nl <= NOT((fsm_output(2)) OR mux_110_nl);
  nor_1268_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(7))) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  or_109_nl <= (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10));
  or_108_nl <= (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(5)) OR (fsm_output(10));
  mux_107_nl <= MUX_s_1_2_2(or_109_nl, or_108_nl, fsm_output(0));
  nor_1269_nl <= NOT((fsm_output(7)) OR mux_107_nl);
  nor_1270_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR not_tmp_45);
  mux_108_nl <= MUX_s_1_2_2(nor_1269_nl, nor_1270_nl, fsm_output(8));
  mux_109_nl <= MUX_s_1_2_2(nor_1268_nl, mux_108_nl, fsm_output(2));
  mux_111_nl <= MUX_s_1_2_2(nor_1267_nl, mux_109_nl, fsm_output(4));
  mux_113_nl <= MUX_s_1_2_2(mux_112_nl, mux_111_nl, fsm_output(6));
  nor_1271_nl <= NOT((NOT (fsm_output(8))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(5)) OR (fsm_output(10)));
  nor_1272_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(7)) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(9)) OR (NOT (fsm_output(5))) OR (fsm_output(10)));
  mux_104_nl <= MUX_s_1_2_2(nor_1271_nl, nor_1272_nl, fsm_output(2));
  and_795_nl <= (fsm_output(3)) AND (fsm_output(9)) AND (fsm_output(5)) AND (NOT
      (fsm_output(10)));
  nor_1273_nl <= NOT((fsm_output(3)) OR (fsm_output(9)) OR not_tmp_45);
  mux_102_nl <= MUX_s_1_2_2(and_795_nl, nor_1273_nl, fsm_output(0));
  and_794_nl <= (NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01"))))
      AND mux_102_nl;
  nor_1274_nl <= NOT((NOT (fsm_output(8))) OR (fsm_output(7)) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(5)) OR (fsm_output(10)));
  mux_103_nl <= MUX_s_1_2_2(and_794_nl, nor_1274_nl, fsm_output(2));
  mux_105_nl <= MUX_s_1_2_2(mux_104_nl, mux_103_nl, fsm_output(4));
  or_98_nl <= (NOT (fsm_output(8))) OR (NOT (fsm_output(7))) OR (fsm_output(0)) OR
      (fsm_output(3)) OR (fsm_output(9)) OR not_tmp_45;
  or_95_nl <= (NOT (fsm_output(3))) OR (fsm_output(9)) OR (fsm_output(5)) OR (NOT
      (fsm_output(10)));
  or_93_nl <= (fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(5)) OR (NOT
      (fsm_output(10)));
  mux_100_nl <= MUX_s_1_2_2(or_95_nl, or_93_nl, fsm_output(0));
  or_96_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")) OR mux_100_nl;
  mux_101_nl <= MUX_s_1_2_2(or_98_nl, or_96_nl, fsm_output(2));
  nor_1275_nl <= NOT((fsm_output(4)) OR mux_101_nl);
  mux_106_nl <= MUX_s_1_2_2(mux_105_nl, nor_1275_nl, fsm_output(6));
  mux_114_nl <= MUX_s_1_2_2(mux_113_nl, mux_106_nl, fsm_output(1));
  nor_1303_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(10)));
  mux_2862_nl <= MUX_s_1_2_2(nor_1303_nl, (fsm_output(10)), fsm_output(6));
  mux_2863_nl <= MUX_s_1_2_2((NOT mux_2862_nl), mux_tmp_2796, fsm_output(7));
  mux_2861_nl <= MUX_s_1_2_2(or_tmp_4, or_tmp_434, fsm_output(7));
  mux_2864_nl <= MUX_s_1_2_2(mux_2863_nl, mux_2861_nl, fsm_output(5));
  mux_2858_nl <= MUX_s_1_2_2(and_dcpl_109, (fsm_output(10)), and_573_cse);
  and_506_nl <= (fsm_output(6)) AND mux_2858_nl;
  and_508_nl <= (fsm_output(6)) AND (NOT nor_tmp_9);
  mux_2859_nl <= MUX_s_1_2_2(and_506_nl, and_508_nl, fsm_output(7));
  or_2643_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(3)) OR (NOT
      (fsm_output(10)));
  mux_2856_nl <= MUX_s_1_2_2(or_2643_nl, or_tmp_2253, fsm_output(6));
  mux_2855_nl <= MUX_s_1_2_2(or_tmp_21, nor_tmp_300, fsm_output(6));
  mux_2857_nl <= MUX_s_1_2_2((NOT mux_2856_nl), mux_2855_nl, fsm_output(7));
  mux_2860_nl <= MUX_s_1_2_2(mux_2859_nl, mux_2857_nl, fsm_output(5));
  mux_2865_nl <= MUX_s_1_2_2((NOT mux_2864_nl), mux_2860_nl, fsm_output(2));
  mux_2852_nl <= MUX_s_1_2_2(or_tmp_2293, or_tmp_2280, fsm_output(7));
  mux_2849_nl <= MUX_s_1_2_2(nor_tmp_6, mux_tmp_2239, nor_412_cse);
  mux_2850_nl <= MUX_s_1_2_2((NOT and_dcpl_240), mux_2849_nl, fsm_output(6));
  and_346_nl <= (fsm_output(6)) AND (and_573_cse OR (fsm_output(3)) OR (NOT (fsm_output(10))));
  mux_2851_nl <= MUX_s_1_2_2(mux_2850_nl, and_346_nl, fsm_output(7));
  mux_2853_nl <= MUX_s_1_2_2((NOT mux_2852_nl), mux_2851_nl, fsm_output(5));
  mux_2846_nl <= MUX_s_1_2_2((NOT nor_tmp_300), mux_tmp_2800, fsm_output(6));
  mux_2847_nl <= MUX_s_1_2_2(and_dcpl_243, mux_2846_nl, fsm_output(7));
  mux_2844_nl <= MUX_s_1_2_2((NOT mux_tmp_2362), nor_tmp_6, fsm_output(6));
  mux_2845_nl <= MUX_s_1_2_2(mux_2844_nl, and_tmp_16, fsm_output(7));
  mux_2848_nl <= MUX_s_1_2_2(mux_2847_nl, mux_2845_nl, fsm_output(5));
  mux_2854_nl <= MUX_s_1_2_2(mux_2853_nl, mux_2848_nl, fsm_output(2));
  mux_2866_nl <= MUX_s_1_2_2(mux_2865_nl, mux_2854_nl, fsm_output(8));
  mux_2840_nl <= MUX_s_1_2_2(not_tmp_378, mux_tmp_2813, fsm_output(7));
  or_2639_nl <= (fsm_output(6)) OR (NOT mux_tmp_2800);
  or_2638_nl <= (fsm_output(6)) OR (NOT or_tmp_2289);
  mux_2839_nl <= MUX_s_1_2_2(or_2639_nl, or_2638_nl, fsm_output(7));
  mux_2841_nl <= MUX_s_1_2_2(mux_2840_nl, mux_2839_nl, fsm_output(5));
  or_2637_nl <= (fsm_output(6)) OR (NOT and_dcpl_240);
  mux_2837_nl <= MUX_s_1_2_2(not_tmp_426, or_2637_nl, fsm_output(7));
  or_2636_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(10));
  mux_2835_nl <= MUX_s_1_2_2((NOT nand_402_cse), or_2636_nl, fsm_output(6));
  mux_2836_nl <= MUX_s_1_2_2(or_36_cse, mux_2835_nl, fsm_output(7));
  mux_2838_nl <= MUX_s_1_2_2(mux_2837_nl, mux_2836_nl, fsm_output(5));
  mux_2842_nl <= MUX_s_1_2_2(mux_2841_nl, mux_2838_nl, fsm_output(2));
  or_3347_nl <= (fsm_output(6)) OR (NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT mux_tmp_2239)));
  mux_2831_nl <= MUX_s_1_2_2((fsm_output(10)), (NOT or_tmp_2233), fsm_output(6));
  mux_2832_nl <= MUX_s_1_2_2(or_3347_nl, mux_2831_nl, fsm_output(7));
  mux_2829_nl <= MUX_s_1_2_2(or_tmp_21, mux_tmp_2254, fsm_output(6));
  or_2632_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (NOT
      nor_tmp_6);
  mux_2828_nl <= MUX_s_1_2_2(or_2632_nl, mux_tmp_2250, fsm_output(6));
  mux_2830_nl <= MUX_s_1_2_2(mux_2829_nl, mux_2828_nl, fsm_output(7));
  mux_2833_nl <= MUX_s_1_2_2(mux_2832_nl, mux_2830_nl, fsm_output(5));
  mux_2825_nl <= MUX_s_1_2_2(and_dcpl_110, or_tmp_2483, fsm_output(6));
  mux_2826_nl <= MUX_s_1_2_2(mux_2825_nl, (NOT mux_tmp_2349), fsm_output(7));
  mux_2823_nl <= MUX_s_1_2_2(and_dcpl_101, or_tmp_2266, fsm_output(6));
  mux_2824_nl <= MUX_s_1_2_2((NOT mux_2823_nl), or_tmp_4, fsm_output(7));
  mux_2827_nl <= MUX_s_1_2_2(mux_2826_nl, mux_2824_nl, fsm_output(5));
  mux_2834_nl <= MUX_s_1_2_2(mux_2833_nl, mux_2827_nl, fsm_output(2));
  mux_2843_nl <= MUX_s_1_2_2(mux_2842_nl, mux_2834_nl, fsm_output(8));
  mux_2867_nl <= MUX_s_1_2_2((NOT mux_2866_nl), mux_2843_nl, fsm_output(4));
  nor_680_nl <= NOT((fsm_output(6)) OR and_dcpl_102);
  mux_2818_nl <= MUX_s_1_2_2(nor_680_nl, or_tmp_4, fsm_output(7));
  mux_2817_nl <= MUX_s_1_2_2(or_tmp_3, or_tmp_2246, fsm_output(7));
  mux_2819_nl <= MUX_s_1_2_2(mux_2818_nl, mux_2817_nl, fsm_output(5));
  mux_2815_nl <= MUX_s_1_2_2(not_tmp_463, or_tmp_3, fsm_output(7));
  mux_2814_nl <= MUX_s_1_2_2(mux_tmp_2813, or_tmp_2474, fsm_output(7));
  mux_2816_nl <= MUX_s_1_2_2(mux_2815_nl, mux_2814_nl, fsm_output(5));
  mux_2820_nl <= MUX_s_1_2_2(mux_2819_nl, mux_2816_nl, fsm_output(2));
  or_2629_nl <= (NOT((fsm_output(3)) OR (NOT (fsm_output(1))))) OR (fsm_output(10));
  mux_2809_nl <= MUX_s_1_2_2(or_2629_nl, or_tmp_2238, fsm_output(6));
  mux_2810_nl <= MUX_s_1_2_2(or_tmp_2276, mux_2809_nl, fsm_output(7));
  nand_128_nl <= NOT((fsm_output(6)) AND (NOT((NOT((fsm_output(1)) OR (NOT (fsm_output(3)))))
      OR (fsm_output(10)))));
  mux_2808_nl <= MUX_s_1_2_2(or_tmp_14, nand_128_nl, fsm_output(7));
  mux_2811_nl <= MUX_s_1_2_2(mux_2810_nl, mux_2808_nl, fsm_output(5));
  mux_2806_nl <= MUX_s_1_2_2(or_tmp_2246, or_tmp_2474, fsm_output(7));
  mux_2805_nl <= MUX_s_1_2_2(mux_9_cse, nand_tmp_95, fsm_output(7));
  mux_2807_nl <= MUX_s_1_2_2(mux_2806_nl, mux_2805_nl, fsm_output(5));
  mux_2812_nl <= MUX_s_1_2_2(mux_2811_nl, mux_2807_nl, fsm_output(2));
  mux_2821_nl <= MUX_s_1_2_2(mux_2820_nl, mux_2812_nl, fsm_output(8));
  nand_127_nl <= NOT((fsm_output(6)) AND (NOT mux_tmp_2800));
  or_2626_nl <= (fsm_output(6)) OR (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(10));
  mux_2801_nl <= MUX_s_1_2_2(nand_127_nl, or_2626_nl, fsm_output(7));
  or_2625_nl <= (fsm_output(6)) OR (NOT nor_tmp_288);
  or_2624_nl <= (fsm_output(6)) OR (nand_237_cse AND (fsm_output(3))) OR (fsm_output(10));
  mux_2798_nl <= MUX_s_1_2_2(or_2625_nl, or_2624_nl, fsm_output(7));
  mux_2802_nl <= MUX_s_1_2_2(mux_2801_nl, mux_2798_nl, fsm_output(5));
  or_2622_nl <= (fsm_output(7)) OR mux_tmp_2796;
  or_2620_nl <= (fsm_output(0)) OR (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(10));
  mux_2794_nl <= MUX_s_1_2_2((fsm_output(10)), or_2620_nl, fsm_output(6));
  mux_2795_nl <= MUX_s_1_2_2(or_tmp_434, mux_2794_nl, fsm_output(7));
  mux_2797_nl <= MUX_s_1_2_2(or_2622_nl, mux_2795_nl, fsm_output(5));
  mux_2803_nl <= MUX_s_1_2_2(mux_2802_nl, mux_2797_nl, fsm_output(2));
  mux_2791_nl <= MUX_s_1_2_2(mux_9_cse, mux_tmp_2790, fsm_output(7));
  nand_126_nl <= NOT((fsm_output(6)) AND (NOT or_tmp_2233));
  mux_2789_nl <= MUX_s_1_2_2(mux_tmp_2788, nand_126_nl, fsm_output(7));
  mux_2792_nl <= MUX_s_1_2_2(mux_2791_nl, mux_2789_nl, fsm_output(5));
  mux_2786_nl <= MUX_s_1_2_2(or_tmp_2257, mux_7_cse, fsm_output(7));
  mux_2787_nl <= MUX_s_1_2_2(mux_2786_nl, mux_3_cse, fsm_output(5));
  mux_2793_nl <= MUX_s_1_2_2(mux_2792_nl, mux_2787_nl, fsm_output(2));
  mux_2804_nl <= MUX_s_1_2_2(mux_2803_nl, mux_2793_nl, fsm_output(8));
  mux_2822_nl <= MUX_s_1_2_2(mux_2821_nl, mux_2804_nl, fsm_output(4));
  COMP_LOOP_COMP_LOOP_and_17_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 1)=STD_LOGIC_VECTOR'("0011"));
  COMP_LOOP_1_acc_8_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_4_dfm) -
      SIGNED(modulo_result_mux_1_cse), 64));
  or_2838_nl <= (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(9))) OR (NOT
      (fsm_output(4))) OR (fsm_output(10));
  mux_3178_nl <= MUX_s_1_2_2(nand_tmp_148, or_2838_nl, fsm_output(0));
  mux_3179_nl <= MUX_s_1_2_2(or_2839_cse, mux_3178_nl, fsm_output(7));
  nor_620_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"))
      OR mux_3179_nl);
  nor_621_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(1)) OR (fsm_output(9)) OR nand_398_cse);
  nor_622_nl <= NOT((fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT
      (fsm_output(9))) OR (fsm_output(4)) OR (fsm_output(10)));
  mux_3175_nl <= MUX_s_1_2_2(and_464_cse, nor_622_nl, fsm_output(7));
  nor_623_nl <= NOT((fsm_output(7)) OR (fsm_output(0)) OR (fsm_output(3)) OR (NOT
      (fsm_output(1))) OR (fsm_output(9)) OR (fsm_output(4)) OR (fsm_output(10)));
  mux_3176_nl <= MUX_s_1_2_2(mux_3175_nl, nor_623_nl, fsm_output(5));
  mux_3177_nl <= MUX_s_1_2_2(nor_621_nl, mux_3176_nl, fsm_output(6));
  mux_3180_nl <= MUX_s_1_2_2(nor_620_nl, mux_3177_nl, fsm_output(8));
  nor_624_nl <= NOT((fsm_output(7)) OR (fsm_output(0)) OR nand_226_cse);
  or_2828_nl <= (fsm_output(1)) OR (fsm_output(9)) OR (NOT (fsm_output(4))) OR (fsm_output(10));
  or_2827_nl <= (fsm_output(1)) OR (NOT (fsm_output(9))) OR (fsm_output(4)) OR (fsm_output(10));
  mux_3170_nl <= MUX_s_1_2_2(or_2828_nl, or_2827_nl, fsm_output(3));
  mux_3171_nl <= MUX_s_1_2_2(mux_3170_nl, or_2826_cse, fsm_output(0));
  nor_625_nl <= NOT((fsm_output(7)) OR mux_3171_nl);
  mux_3172_nl <= MUX_s_1_2_2(nor_624_nl, nor_625_nl, fsm_output(5));
  mux_3169_nl <= MUX_s_1_2_2(or_2824_cse, nand_tmp_148, fsm_output(0));
  and_465_nl <= (fsm_output(5)) AND (fsm_output(7)) AND (NOT mux_3169_nl);
  mux_3173_nl <= MUX_s_1_2_2(mux_3172_nl, and_465_nl, fsm_output(6));
  or_2817_nl <= (NOT (fsm_output(0))) OR (fsm_output(3)) OR (NOT (fsm_output(1)))
      OR (fsm_output(9)) OR (fsm_output(4)) OR (fsm_output(10));
  mux_3167_nl <= MUX_s_1_2_2(or_2819_cse, or_2817_nl, fsm_output(7));
  nor_626_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10"))
      OR mux_3167_nl);
  mux_3174_nl <= MUX_s_1_2_2(mux_3173_nl, nor_626_nl, fsm_output(8));
  mux_3181_nl <= MUX_s_1_2_2(mux_3180_nl, mux_3174_nl, fsm_output(2));
  COMP_LOOP_COMP_LOOP_and_10_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_11_0(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  COMP_LOOP_1_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(COMP_LOOP_k_9_4_sva_2
      & STD_LOGIC_VECTOR'( "0000")) + SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(9
      DOWNTO 1)))) + SIGNED'( "0000000001"), 10));
  nor_nl <= NOT((fsm_output(10)) OR (fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6))
      OR and_359_cse);
  mux_3215_nl <= MUX_s_1_2_2(and_458_cse, and_459_cse, fsm_output(0));
  or_3259_nl <= (fsm_output(5)) OR ((fsm_output(4)) AND mux_3215_nl);
  nor_617_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000"))
      OR and_563_cse);
  mux_3216_nl <= MUX_s_1_2_2(or_3259_nl, nor_617_nl, fsm_output(6));
  or_2888_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000000"));
  mux_3217_nl <= MUX_s_1_2_2(mux_3216_nl, or_2888_nl, fsm_output(7));
  and_1253_nl <= (fsm_output(10)) AND ((fsm_output(8)) OR mux_3217_nl);
  mux_3223_nl <= MUX_s_1_2_2(mux_tmp_3219, nor_tmp_445, fsm_output(6));
  mux_3220_nl <= MUX_s_1_2_2(mux_tmp_3219, nor_tmp_445, or_2898_cse);
  and_452_nl <= (and_517_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")))
      AND (fsm_output(9));
  mux_3221_nl <= MUX_s_1_2_2(mux_3220_nl, and_452_nl, fsm_output(1));
  and_454_nl <= (and_528_cse OR CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")))
      AND (fsm_output(9));
  mux_3222_nl <= MUX_s_1_2_2(mux_3221_nl, and_454_nl, fsm_output(2));
  mux_3224_nl <= MUX_s_1_2_2(mux_3223_nl, mux_3222_nl, and_456_cse);
  mux_3231_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), and_528_cse, fsm_output(7));
  mux_3232_nl <= MUX_s_1_2_2(and_dcpl_268, mux_3231_nl, fsm_output(5));
  and_363_nl <= (fsm_output(6)) AND or_2902_cse;
  mux_3229_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), and_363_nl, fsm_output(7));
  mux_3230_nl <= MUX_s_1_2_2(and_dcpl_268, mux_3229_nl, fsm_output(5));
  mux_3233_nl <= MUX_s_1_2_2(mux_3232_nl, mux_3230_nl, fsm_output(2));
  nor_729_nl <= NOT((fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3)));
  mux_3226_nl <= MUX_s_1_2_2(nor_729_nl, (fsm_output(6)), fsm_output(7));
  mux_3227_nl <= MUX_s_1_2_2(and_dcpl_268, mux_3226_nl, fsm_output(5));
  mux_3225_nl <= MUX_s_1_2_2(and_dcpl_268, and_450_cse, fsm_output(5));
  mux_3228_nl <= MUX_s_1_2_2(mux_3227_nl, mux_3225_nl, fsm_output(2));
  mux_3234_nl <= MUX_s_1_2_2(mux_3233_nl, mux_3228_nl, fsm_output(4));
  mux_3239_nl <= MUX_s_1_2_2((fsm_output(7)), or_2520_cse, fsm_output(5));
  or_2906_nl <= (fsm_output(7)) OR and_528_cse;
  mux_3238_nl <= MUX_s_1_2_2(or_2906_nl, or_2520_cse, fsm_output(5));
  mux_3240_nl <= MUX_s_1_2_2(mux_3239_nl, mux_3238_nl, fsm_output(2));
  mux_3241_nl <= MUX_s_1_2_2(and_dcpl_268, mux_3240_nl, fsm_output(8));
  mux_3237_nl <= MUX_s_1_2_2((NOT mux_tmp_3236), or_2520_cse, fsm_output(8));
  mux_3242_nl <= MUX_s_1_2_2(mux_3241_nl, mux_3237_nl, fsm_output(4));
  or_3252_nl <= (fsm_output(8)) OR and_359_cse OR (fsm_output(6));
  nand_218_nl <= NOT((fsm_output(8)) AND (((CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")))
      AND CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))) OR (fsm_output(6))));
  mux_3243_nl <= MUX_s_1_2_2(or_3252_nl, nand_218_nl, fsm_output(7));
  mux_3248_nl <= MUX_s_1_2_2(mux_tmp_3244, or_tmp_2849, fsm_output(5));
  mux_3245_nl <= MUX_s_1_2_2(mux_tmp_3244, or_tmp_2849, and_563_cse);
  or_2915_nl <= (NOT((fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(7))
      OR (fsm_output(8)))) OR (fsm_output(9));
  mux_3246_nl <= MUX_s_1_2_2(mux_3245_nl, or_2915_nl, fsm_output(5));
  or_2913_nl <= (NOT(CONV_SL_1_1(fsm_output(8 DOWNTO 5)/=STD_LOGIC_VECTOR'("0000"))))
      OR (fsm_output(9));
  mux_3247_nl <= MUX_s_1_2_2(mux_3246_nl, or_2913_nl, fsm_output(3));
  mux_3249_nl <= MUX_s_1_2_2(mux_3248_nl, mux_3247_nl, fsm_output(4));
  nor_1317_nl <= NOT((fsm_output(8)) OR mux_tmp_3236);
  mux_3250_nl <= MUX_s_1_2_2(nor_1316_cse, nor_1317_nl, fsm_output(4));
  or_3346_nl <= (fsm_output(8)) OR (CONV_SL_1_1(fsm_output(7 DOWNTO 5)=STD_LOGIC_VECTOR'("111")));
  mux_3251_nl <= MUX_s_1_2_2(mux_3250_nl, or_3346_nl, fsm_output(9));
  nor_611_nl <= NOT((fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(8))
      OR (fsm_output(9)));
  mux_3253_nl <= MUX_s_1_2_2(nor_610_cse, nor_611_nl, and_456_cse);
  and_371_nl <= (fsm_output(2)) AND or_2348_cse AND CONV_SL_1_1(fsm_output(9 DOWNTO
      8)=STD_LOGIC_VECTOR'("11"));
  or_2922_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000"));
  mux_3252_nl <= MUX_s_1_2_2(and_371_nl, nor_tmp_116, or_2922_nl);
  mux_3254_nl <= MUX_s_1_2_2(mux_3253_nl, mux_3252_nl, fsm_output(6));
  mux_3255_nl <= MUX_s_1_2_2(mux_3254_nl, nor_tmp_116, fsm_output(7));
  mux_3259_nl <= MUX_s_1_2_2(mux_tmp_3256, nor_tmp_456, fsm_output(3));
  mux_3260_nl <= MUX_s_1_2_2(not_tmp_728, mux_3259_nl, fsm_output(4));
  mux_3257_nl <= MUX_s_1_2_2(not_tmp_728, mux_tmp_3256, fsm_output(3));
  mux_3258_nl <= MUX_s_1_2_2(mux_3257_nl, nor_tmp_456, fsm_output(4));
  mux_3261_nl <= MUX_s_1_2_2(mux_3260_nl, mux_3258_nl, or_2385_cse);
  mux_3262_nl <= MUX_s_1_2_2(not_tmp_728, mux_3261_nl, fsm_output(5));
  mux_3263_nl <= MUX_s_1_2_2(mux_3262_nl, nor_tmp_456, fsm_output(6));
  or_2933_nl <= CONV_SL_1_1(fsm_output(9 DOWNTO 6)/=STD_LOGIC_VECTOR'("0000"));
  mux_3265_nl <= MUX_s_1_2_2((NOT (fsm_output(10))), (fsm_output(10)), or_2933_nl);
  mux_3266_nl <= MUX_s_1_2_2(mux_3265_nl, or_tmp_2864, and_440_cse);
  mux_3267_nl <= MUX_s_1_2_2(mux_3266_nl, or_tmp_2864, fsm_output(5));
  or_2930_nl <= (NOT((fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(7)) OR (fsm_output(8)) OR (fsm_output(9)))) OR (fsm_output(10));
  mux_3264_nl <= MUX_s_1_2_2(or_tmp_2864, or_2930_nl, fsm_output(5));
  mux_3275_nl <= MUX_s_1_2_2(and_dcpl_264, (fsm_output(10)), or_2935_cse);
  mux_3271_nl <= MUX_s_1_2_2(mux_tmp_2220, (fsm_output(10)), fsm_output(7));
  mux_3272_nl <= MUX_s_1_2_2(mux_tmp_3269, mux_3271_nl, fsm_output(5));
  and_439_nl <= or_2520_cse AND (fsm_output(10));
  mux_3270_nl <= MUX_s_1_2_2(mux_tmp_3269, and_439_nl, fsm_output(5));
  mux_3273_nl <= MUX_s_1_2_2(mux_3272_nl, mux_3270_nl, fsm_output(2));
  mux_3274_nl <= MUX_s_1_2_2(mux_3273_nl, (fsm_output(10)), fsm_output(8));
  mux_3276_nl <= MUX_s_1_2_2(mux_3275_nl, mux_3274_nl, fsm_output(4));
  mux_3288_nl <= MUX_s_1_2_2(mux_tmp_3281, mux_tmp_3280, fsm_output(5));
  and_434_nl <= (fsm_output(0)) AND (fsm_output(3));
  mux_3285_nl <= MUX_s_1_2_2(mux_tmp_3281, mux_tmp_3280, and_434_nl);
  mux_3284_nl <= MUX_s_1_2_2(mux_tmp_3280, nor_tmp_461, fsm_output(3));
  mux_3286_nl <= MUX_s_1_2_2(mux_3285_nl, mux_3284_nl, fsm_output(5));
  mux_3282_nl <= MUX_s_1_2_2(mux_tmp_3281, mux_tmp_3280, fsm_output(3));
  mux_3283_nl <= MUX_s_1_2_2(mux_3282_nl, nor_tmp_461, fsm_output(5));
  mux_3287_nl <= MUX_s_1_2_2(mux_3286_nl, mux_3283_nl, or_2385_cse);
  nor_604_nl <= NOT((fsm_output(8)) OR (fsm_output(10)));
  nor_605_nl <= NOT((fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(10)));
  and_431_nl <= (fsm_output(2)) AND (fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(10));
  mux_3290_nl <= MUX_s_1_2_2(nor_605_nl, and_431_nl, fsm_output(1));
  mux_3291_nl <= MUX_s_1_2_2(nor_604_nl, mux_3290_nl, and_456_cse);
  and_433_nl <= (fsm_output(8)) AND (fsm_output(10));
  mux_3292_nl <= MUX_s_1_2_2(mux_3291_nl, and_433_nl, or_2520_cse);
  or_2947_nl <= (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(10));
  mux_3296_nl <= MUX_s_1_2_2((fsm_output(10)), or_2947_nl, and_456_cse);
  nor_603_nl <= NOT((fsm_output(8)) OR (fsm_output(6)) OR mux_3296_nl);
  and_430_nl <= (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(10));
  or_2945_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"));
  mux_3294_nl <= MUX_s_1_2_2(and_430_nl, (fsm_output(10)), or_2945_nl);
  and_374_nl <= (fsm_output(5)) AND mux_3294_nl;
  mux_3295_nl <= MUX_s_1_2_2(and_374_nl, (fsm_output(10)), fsm_output(6));
  and_375_nl <= (fsm_output(8)) AND mux_3295_nl;
  mux_3297_nl <= MUX_s_1_2_2(nor_603_nl, and_375_nl, fsm_output(7));
  or_2950_nl <= (fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(6))
      OR (fsm_output(7)) OR (fsm_output(8));
  mux_3299_nl <= MUX_s_1_2_2(or_2951_cse, or_2950_nl, and_456_cse);
  nor_1420_nl <= NOT((fsm_output(10)) OR mux_3299_nl);
  and_1254_nl <= (fsm_output(10)) AND (CONV_SL_1_1(fsm_output(8 DOWNTO 3)/=STD_LOGIC_VECTOR'("000000")));
  nor_1201_nl <= NOT((fsm_output(6)) OR (fsm_output(9)) OR (fsm_output(10)));
  mux_3302_nl <= MUX_s_1_2_2(nor_601_cse, nor_1203_cse, fsm_output(4));
  and_29_nl <= (fsm_output(2)) AND or_2348_cse AND (fsm_output(3)) AND (fsm_output(9))
      AND (fsm_output(10));
  mux_3301_nl <= MUX_s_1_2_2(and_29_nl, and_816_cse, fsm_output(4));
  mux_3303_nl <= MUX_s_1_2_2(mux_3302_nl, mux_3301_nl, fsm_output(6));
  mux_3304_nl <= MUX_s_1_2_2(nor_1201_nl, mux_3303_nl, fsm_output(5));
  COMP_LOOP_COMP_LOOP_or_15_nl <= (VEC_LOOP_j_sva_11_0(11)) OR and_850_cse OR and_857_cse
      OR and_dcpl_378 OR and_869_cse OR and_875_cse OR and_dcpl_394 OR and_886_cse
      OR and_dcpl_404 OR and_dcpl_408 OR and_dcpl_411 OR and_dcpl_415;
  COMP_LOOP_COMP_LOOP_mux_18_nl <= MUX_v_9_2_2((VEC_LOOP_j_sva_11_0(10 DOWNTO 2)),
      (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 1))), COMP_LOOP_or_60_itm);
  COMP_LOOP_or_77_nl <= (NOT and_dcpl_356) OR and_850_cse OR and_857_cse OR and_dcpl_378
      OR and_869_cse OR and_875_cse OR and_dcpl_394 OR and_886_cse OR and_dcpl_404
      OR and_dcpl_408 OR and_dcpl_411 OR and_dcpl_415;
  COMP_LOOP_COMP_LOOP_mux_19_nl <= MUX_v_5_2_2((STD_LOGIC_VECTOR'( "00") & (COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 2))), COMP_LOOP_k_9_4_sva_4_0, COMP_LOOP_or_60_itm);
  COMP_LOOP_COMP_LOOP_or_16_nl <= ((COMP_LOOP_k_9_4_sva_4_0(1)) AND (NOT(and_850_cse
      OR and_857_cse OR and_dcpl_378 OR and_869_cse OR and_875_cse))) OR and_dcpl_394
      OR and_886_cse OR and_dcpl_404 OR and_dcpl_408 OR and_dcpl_411 OR and_dcpl_415;
  COMP_LOOP_COMP_LOOP_or_17_nl <= ((COMP_LOOP_k_9_4_sva_4_0(0)) AND (NOT(and_850_cse
      OR and_857_cse OR and_dcpl_394 OR and_886_cse OR and_dcpl_404))) OR and_dcpl_378
      OR and_869_cse OR and_875_cse OR and_dcpl_408 OR and_dcpl_411 OR and_dcpl_415;
  COMP_LOOP_COMP_LOOP_or_18_nl <= (NOT(and_dcpl_356 OR and_850_cse OR and_dcpl_378
      OR and_869_cse OR and_dcpl_394 OR and_886_cse OR and_dcpl_408 OR and_dcpl_411))
      OR and_857_cse OR and_875_cse OR and_dcpl_404 OR and_dcpl_415;
  COMP_LOOP_COMP_LOOP_or_19_nl <= (NOT(and_857_cse OR and_dcpl_378 OR and_875_cse
      OR and_dcpl_394 OR and_dcpl_404 OR and_dcpl_408 OR and_dcpl_415)) OR and_dcpl_356
      OR and_850_cse OR and_869_cse OR and_886_cse OR and_dcpl_411;
  acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_15_nl
      & COMP_LOOP_COMP_LOOP_mux_18_nl & COMP_LOOP_or_77_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_mux_19_nl
      & COMP_LOOP_COMP_LOOP_or_16_nl & COMP_LOOP_COMP_LOOP_or_17_nl & COMP_LOOP_COMP_LOOP_or_18_nl
      & COMP_LOOP_COMP_LOOP_or_19_nl & '1'), 10), 11), 11));
  z_out <= acc_nl(10 DOWNTO 1);
  COMP_LOOP_mux_84_nl <= MUX_v_10_2_2((VEC_LOOP_j_sva_11_0(11 DOWNTO 2)), STAGE_LOOP_lshift_psp_sva,
      COMP_LOOP_or_24_itm);
  COMP_LOOP_COMP_LOOP_mux_20_nl <= MUX_v_5_2_2((STD_LOGIC_VECTOR'( "00") & (COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 2))), COMP_LOOP_k_9_4_sva_4_0, COMP_LOOP_or_24_itm);
  COMP_LOOP_mux_85_nl <= MUX_v_2_2_2((COMP_LOOP_k_9_4_sva_4_0(1 DOWNTO 0)), STD_LOGIC_VECTOR'(
      "01"), and_dcpl_433);
  COMP_LOOP_COMP_LOOP_or_20_nl <= MUX_v_2_2_2(COMP_LOOP_mux_85_nl, STD_LOGIC_VECTOR'("11"),
      and_dcpl_441);
  z_out_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_84_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_mux_20_nl
      & COMP_LOOP_COMP_LOOP_or_20_nl & COMP_LOOP_COMP_LOOP_or_6_cse & COMP_LOOP_COMP_LOOP_or_6_cse),
      9), 10), 10));
  and_1278_nl <= and_dcpl_353 AND (NOT (fsm_output(9))) AND (NOT (fsm_output(8)))
      AND (fsm_output(7)) AND (fsm_output(5)) AND (fsm_output(3)) AND (fsm_output(2))
      AND (fsm_output(1)) AND and_dcpl_107;
  and_1279_nl <= (NOT (fsm_output(4))) AND (NOT (fsm_output(10))) AND (NOT (fsm_output(9)))
      AND and_dcpl_373 AND (NOT (fsm_output(5))) AND (fsm_output(3)) AND (NOT (fsm_output(2)))
      AND (NOT (fsm_output(1))) AND and_dcpl_107;
  and_1280_nl <= (NOT (fsm_output(4))) AND (fsm_output(10)) AND (NOT (fsm_output(9)))
      AND and_dcpl_373 AND (fsm_output(5)) AND and_dcpl_348 AND (NOT (fsm_output(1)))
      AND (fsm_output(6)) AND (NOT (fsm_output(0)));
  COMP_LOOP_mux1h_585_nl <= MUX1HOT_v_4_4_2(STD_LOGIC_VECTOR'( "0001"), STD_LOGIC_VECTOR'(
      "0011"), STD_LOGIC_VECTOR'( "0101"), STD_LOGIC_VECTOR'( "1110"), STD_LOGIC_VECTOR'(
      and_1278_nl & and_1279_nl & (fsm_output(9)) & and_1280_nl));
  z_out_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_lshift_psp_sva) +
      CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & COMP_LOOP_mux1h_585_nl),
      9), 10), 10));
  and_1281_nl <= and_dcpl_503 AND (NOT (fsm_output(9))) AND and_dcpl_502 AND (fsm_output(3))
      AND (fsm_output(2)) AND (NOT (fsm_output(1))) AND (fsm_output(6)) AND (NOT
      (fsm_output(0)));
  COMP_LOOP_mux_86_nl <= MUX_v_2_2_2(STD_LOGIC_VECTOR'( "10"), STD_LOGIC_VECTOR'(
      "01"), and_1281_nl);
  and_1282_nl <= (NOT (fsm_output(10))) AND (NOT (fsm_output(4))) AND (NOT (fsm_output(9)))
      AND (fsm_output(8)) AND (NOT (fsm_output(7))) AND (fsm_output(5)) AND and_dcpl_480
      AND and_dcpl_99;
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl <= NOT(MUX_v_2_2_2(COMP_LOOP_mux_86_nl,
      STD_LOGIC_VECTOR'("11"), and_1282_nl));
  COMP_LOOP_or_78_nl <= MUX_v_2_2_2(COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_53_nl, STD_LOGIC_VECTOR'("11"),
      and_dcpl_511);
  z_out_3 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_lshift_psp_sva) +
      CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & COMP_LOOP_or_78_nl
      & '1' & and_dcpl_511), 9), 10), 10));
  and_1283_nl <= and_dcpl_375 AND (NOT (fsm_output(9))) AND and_dcpl_517 AND (fsm_output(3))
      AND (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(6)) AND (NOT (fsm_output(0)));
  and_1284_nl <= and_dcpl_375 AND (fsm_output(9)) AND and_dcpl_517 AND CONV_SL_1_1(fsm_output(3
      DOWNTO 1)=STD_LOGIC_VECTOR'("011")) AND nor_tmp_217;
  and_1285_nl <= and_dcpl_406 AND (fsm_output(8)) AND (NOT (fsm_output(7))) AND (fsm_output(5))
      AND (fsm_output(3)) AND (NOT (fsm_output(2))) AND (fsm_output(1)) AND nor_tmp_217;
  COMP_LOOP_mux1h_586_nl <= MUX1HOT_v_4_4_2(STD_LOGIC_VECTOR'( "0100"), STD_LOGIC_VECTOR'(
      "1001"), STD_LOGIC_VECTOR'( "1011"), STD_LOGIC_VECTOR'( "1101"), STD_LOGIC_VECTOR'(
      and_1283_nl & and_1284_nl & (NOT (fsm_output(1))) & and_1285_nl));
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_lshift_psp_sva) +
      CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & COMP_LOOP_mux1h_586_nl),
      9), 10), 10));
  COMP_LOOP_mux1h_587_nl <= MUX1HOT_v_64_3_2((STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000")
      & VEC_LOOP_j_sva_11_0), tmp_10_lpi_4_dfm, ('1' & (NOT (operator_64_false_acc_mut_63_0(62
      DOWNTO 0)))), STD_LOGIC_VECTOR'( and_dcpl_555 & (NOT mux_3724_itm) & and_dcpl_564));
  COMP_LOOP_mux1h_588_nl <= MUX1HOT_v_64_3_2((STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000")
      & COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'( "0011")), modulo_result_mux_1_cse,
      STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
      STD_LOGIC_VECTOR'( and_dcpl_555 & (NOT mux_3724_itm) & and_dcpl_564));
  z_out_5 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux1h_587_nl) + UNSIGNED(COMP_LOOP_mux1h_588_nl),
      64));
  operator_64_false_1_mux1h_2_nl <= MUX1HOT_v_64_4_2((STD_LOGIC_VECTOR'( "00000000000000000000000000000000000000000000000000000000001")
      & (NOT COMP_LOOP_k_9_4_sva_4_0)), modulo_result_rem_cmp_z, p_sva, (STD_LOGIC_VECTOR'(
      "0000000000000000000000000000000000000000000000000000") & VEC_LOOP_j_sva_11_0),
      STD_LOGIC_VECTOR'( and_dcpl_574 & (NOT mux_3788_itm) & and_dcpl_579 & and_dcpl_588));
  operator_64_false_1_mux1h_3_nl <= MUX1HOT_v_64_3_2(STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
      p_sva, (STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000")
      & STAGE_LOOP_lshift_psp_sva), STD_LOGIC_VECTOR'( and_dcpl_574 & (NOT mux_3788_itm)
      & and_dcpl_588));
  operator_64_false_1_or_1_nl <= MUX_v_64_2_2(operator_64_false_1_mux1h_3_nl, STD_LOGIC_VECTOR'("1111111111111111111111111111111111111111111111111111111111111111"),
      and_dcpl_579);
  z_out_6 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(operator_64_false_1_mux1h_2_nl),
      65) + CONV_UNSIGNED(SIGNED(operator_64_false_1_or_1_nl), 65), 65));
  COMP_LOOP_COMP_LOOP_or_21_nl <= (NOT(and_dcpl_598 OR and_850_cse OR and_857_cse
      OR and_dcpl_622 OR and_dcpl_628 OR and_869_cse OR and_875_cse OR and_dcpl_641
      OR and_dcpl_646 OR and_886_cse OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663
      OR and_dcpl_666 OR and_dcpl_669 OR and_dcpl_672 OR and_dcpl_676)) OR and_dcpl_678;
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl <= NOT((operator_66_true_div_cmp_z(63))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl <= NOT((operator_66_true_div_cmp_z(62))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl <= NOT((operator_66_true_div_cmp_z(61))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl <= NOT((operator_66_true_div_cmp_z(60))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl <= NOT((operator_66_true_div_cmp_z(59))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl <= NOT((operator_66_true_div_cmp_z(58))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl <= NOT((operator_66_true_div_cmp_z(57))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl <= NOT((operator_66_true_div_cmp_z(56))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl <= NOT((operator_66_true_div_cmp_z(55))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl <= NOT((operator_66_true_div_cmp_z(54))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl <= NOT((operator_66_true_div_cmp_z(53))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl <= NOT((operator_66_true_div_cmp_z(52))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl <= NOT((operator_66_true_div_cmp_z(51))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl <= NOT((operator_66_true_div_cmp_z(50))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl <= NOT((operator_66_true_div_cmp_z(49))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl <= NOT((operator_66_true_div_cmp_z(48))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl <= NOT((operator_66_true_div_cmp_z(47))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl <= NOT((operator_66_true_div_cmp_z(46))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl <= NOT((operator_66_true_div_cmp_z(45))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl <= NOT((operator_66_true_div_cmp_z(44))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl <= NOT((operator_66_true_div_cmp_z(43))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl <= NOT((operator_66_true_div_cmp_z(42))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl <= NOT((operator_66_true_div_cmp_z(41))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl <= NOT((operator_66_true_div_cmp_z(40))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl <= NOT((operator_66_true_div_cmp_z(39))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl <= NOT((operator_66_true_div_cmp_z(38))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl <= NOT((operator_66_true_div_cmp_z(37))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl <= NOT((operator_66_true_div_cmp_z(36))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl <= NOT((operator_66_true_div_cmp_z(35))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl <= NOT((operator_66_true_div_cmp_z(34))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl <= NOT((operator_66_true_div_cmp_z(33))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl <= NOT((operator_66_true_div_cmp_z(32))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl <= NOT((operator_66_true_div_cmp_z(31))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl <= NOT((operator_66_true_div_cmp_z(30))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl <= NOT((operator_66_true_div_cmp_z(29))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl <= NOT((operator_66_true_div_cmp_z(28))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl <= NOT((operator_66_true_div_cmp_z(27))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl <= NOT((operator_66_true_div_cmp_z(26))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl <= NOT((operator_66_true_div_cmp_z(25))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl <= NOT((operator_66_true_div_cmp_z(24))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl <= NOT((operator_66_true_div_cmp_z(23))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl <= NOT((operator_66_true_div_cmp_z(22))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl <= NOT((operator_66_true_div_cmp_z(21))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl <= NOT((operator_66_true_div_cmp_z(20))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl <= NOT((operator_66_true_div_cmp_z(19))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl <= NOT((operator_66_true_div_cmp_z(18))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl <= NOT((operator_66_true_div_cmp_z(17))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl <= NOT((operator_66_true_div_cmp_z(16))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl <= NOT((operator_66_true_div_cmp_z(15))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl <= NOT((operator_66_true_div_cmp_z(14))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_104_nl <= NOT((operator_66_true_div_cmp_z(13))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_105_nl <= NOT((operator_66_true_div_cmp_z(12))
      OR and_dcpl_598 OR and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676);
  COMP_LOOP_or_79_nl <= and_850_cse OR and_857_cse OR and_dcpl_622 OR and_dcpl_628
      OR and_869_cse OR and_875_cse OR and_dcpl_641 OR and_dcpl_646 OR and_886_cse
      OR and_dcpl_654 OR and_dcpl_659 OR and_dcpl_663 OR and_dcpl_666 OR and_dcpl_669
      OR and_dcpl_672 OR and_dcpl_676;
  COMP_LOOP_mux1h_589_nl <= MUX1HOT_v_12_3_2((STD_LOGIC_VECTOR'( "000000") & COMP_LOOP_k_9_4_sva_4_0
      & '1'), VEC_LOOP_j_sva_11_0, (NOT (operator_66_true_div_cmp_z(11 DOWNTO 0))),
      STD_LOGIC_VECTOR'( and_dcpl_598 & COMP_LOOP_or_79_nl & and_dcpl_678));
  COMP_LOOP_mux1h_590_nl <= MUX1HOT_v_7_7_2(('0' & (VEC_LOOP_j_sva_11_0(11 DOWNTO
      6))), ((z_out_9(5 DOWNTO 0)) & (STAGE_LOOP_lshift_psp_sva(3))), (z_out_2(9
      DOWNTO 3)), (z_out_3(9 DOWNTO 3)), (z_out_4(9 DOWNTO 3)), (z_out_1(9 DOWNTO
      3)), z_out_9, STD_LOGIC_VECTOR'( and_dcpl_598 & and_850_cse & COMP_LOOP_or_55_ssc
      & COMP_LOOP_or_56_ssc & COMP_LOOP_or_57_ssc & COMP_LOOP_or_58_ssc & and_886_cse));
  not_8636_nl <= NOT and_dcpl_678;
  COMP_LOOP_and_285_nl <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), COMP_LOOP_mux1h_590_nl,
      not_8636_nl);
  COMP_LOOP_or_80_nl <= and_850_cse OR and_886_cse;
  COMP_LOOP_mux1h_591_nl <= MUX1HOT_v_3_7_2((VEC_LOOP_j_sva_11_0(5 DOWNTO 3)), (STAGE_LOOP_lshift_psp_sva(2
      DOWNTO 0)), (z_out_2(2 DOWNTO 0)), (z_out_3(2 DOWNTO 0)), (z_out_4(2 DOWNTO
      0)), (z_out_1(2 DOWNTO 0)), STD_LOGIC_VECTOR'( "001"), STD_LOGIC_VECTOR'( and_dcpl_598
      & COMP_LOOP_or_80_nl & COMP_LOOP_or_55_ssc & COMP_LOOP_or_56_ssc & COMP_LOOP_or_57_ssc
      & COMP_LOOP_or_58_ssc & and_dcpl_678));
  z_out_7 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_21_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_54_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_55_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_56_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_57_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_58_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_59_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_60_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_61_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_62_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_63_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_64_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_65_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_66_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_67_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_68_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_69_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_70_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_71_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_72_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_73_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_74_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_75_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_76_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_77_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_78_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_79_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_80_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_81_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_82_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_83_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_84_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_85_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_86_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_87_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_88_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_89_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_90_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_91_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_92_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_93_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_94_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_95_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_96_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_97_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_98_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_99_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_100_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_101_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_102_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_103_nl
      & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_104_nl & COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_105_nl
      & COMP_LOOP_mux1h_589_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_and_285_nl
      & COMP_LOOP_mux1h_591_nl), 10), 65), 65));
  COMP_LOOP_mux_87_nl <= MUX_s_1_2_2((NOT modExp_exp_1_7_1_sva), (NOT COMP_LOOP_nor_134_itm),
      and_dcpl_707);
  COMP_LOOP_COMP_LOOP_or_22_nl <= COMP_LOOP_mux_87_nl OR and_dcpl_688 OR and_dcpl_698;
  COMP_LOOP_mux1h_592_nl <= MUX1HOT_s_1_3_2((NOT (STAGE_LOOP_lshift_psp_sva(9))),
      (NOT modExp_exp_1_6_1_sva), (NOT modExp_exp_1_7_1_sva), STD_LOGIC_VECTOR'(
      COMP_LOOP_or_67_itm & not_tmp_980 & and_dcpl_707));
  COMP_LOOP_mux1h_593_nl <= MUX1HOT_s_1_3_2((NOT (STAGE_LOOP_lshift_psp_sva(8))),
      (NOT modExp_exp_1_5_1_sva), (NOT modExp_exp_1_6_1_sva), STD_LOGIC_VECTOR'(
      COMP_LOOP_or_67_itm & not_tmp_980 & and_dcpl_707));
  COMP_LOOP_mux1h_594_nl <= MUX1HOT_s_1_3_2((NOT (STAGE_LOOP_lshift_psp_sva(7))),
      (NOT modExp_exp_1_4_1_sva), (NOT modExp_exp_1_5_1_sva), STD_LOGIC_VECTOR'(
      COMP_LOOP_or_67_itm & not_tmp_980 & and_dcpl_707));
  COMP_LOOP_mux1h_595_nl <= MUX1HOT_s_1_3_2((NOT (STAGE_LOOP_lshift_psp_sva(6))),
      (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm), (NOT modExp_exp_1_4_1_sva), STD_LOGIC_VECTOR'(
      COMP_LOOP_or_67_itm & not_tmp_980 & and_dcpl_707));
  COMP_LOOP_mux1h_596_nl <= MUX1HOT_s_1_3_2((NOT (STAGE_LOOP_lshift_psp_sva(5))),
      (NOT COMP_LOOP_nor_137_itm), (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm), STD_LOGIC_VECTOR'(
      COMP_LOOP_or_67_itm & not_tmp_980 & and_dcpl_707));
  COMP_LOOP_mux1h_597_nl <= MUX1HOT_s_1_3_2((NOT (STAGE_LOOP_lshift_psp_sva(4))),
      (NOT COMP_LOOP_nor_134_itm), (NOT COMP_LOOP_nor_137_itm), STD_LOGIC_VECTOR'(
      COMP_LOOP_or_67_itm & not_tmp_980 & and_dcpl_707));
  COMP_LOOP_or_81_nl <= not_tmp_980 OR and_dcpl_707;
  COMP_LOOP_COMP_LOOP_mux_21_nl <= MUX_s_1_2_2((NOT (STAGE_LOOP_lshift_psp_sva(3))),
      (NOT COMP_LOOP_nor_12_itm), COMP_LOOP_or_81_nl);
  COMP_LOOP_or_82_nl <= COMP_LOOP_nor_680_itm OR and_dcpl_688 OR and_dcpl_698;
  COMP_LOOP_COMP_LOOP_and_990_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), COMP_LOOP_k_9_4_sva_4_0,
      COMP_LOOP_nor_680_itm);
  COMP_LOOP_COMP_LOOP_or_23_nl <= (NOT(and_dcpl_688 OR not_tmp_980 OR and_dcpl_707))
      OR and_dcpl_698;
  acc_8_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( COMP_LOOP_COMP_LOOP_or_9_cse
      & COMP_LOOP_COMP_LOOP_or_22_nl & COMP_LOOP_mux1h_592_nl & COMP_LOOP_mux1h_593_nl
      & COMP_LOOP_mux1h_594_nl & COMP_LOOP_mux1h_595_nl & COMP_LOOP_mux1h_596_nl
      & COMP_LOOP_mux1h_597_nl & COMP_LOOP_COMP_LOOP_mux_21_nl & COMP_LOOP_or_82_nl)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_and_990_nl & COMP_LOOP_COMP_LOOP_or_23_nl
      & COMP_LOOP_COMP_LOOP_or_9_cse & '1'), 8), 10), 10));
  z_out_8_8_7 <= acc_8_nl(9 DOWNTO 8);
  COMP_LOOP_COMP_LOOP_or_24_nl <= ((STAGE_LOOP_lshift_psp_sva(9)) AND (NOT(and_dcpl_727
      OR and_dcpl_734))) OR and_dcpl_717;
  COMP_LOOP_mux1h_598_nl <= MUX1HOT_v_6_4_2((NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO
      4))), ('1' & (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 5)))), (STAGE_LOOP_lshift_psp_sva(9
      DOWNTO 4)), (STAGE_LOOP_lshift_psp_sva(8 DOWNTO 3)), STD_LOGIC_VECTOR'( and_dcpl_717
      & and_dcpl_727 & and_dcpl_734 & and_dcpl_741));
  COMP_LOOP_or_83_nl <= (NOT(and_dcpl_734 OR and_dcpl_741)) OR and_dcpl_717 OR and_dcpl_727;
  COMP_LOOP_or_84_nl <= and_dcpl_727 OR and_dcpl_734;
  COMP_LOOP_COMP_LOOP_mux_22_nl <= MUX_v_5_2_2(COMP_LOOP_k_9_4_sva_4_0, ('0' & (COMP_LOOP_k_9_4_sva_4_0(4
      DOWNTO 1))), COMP_LOOP_or_84_nl);
  COMP_LOOP_COMP_LOOP_or_25_nl <= ((COMP_LOOP_k_9_4_sva_4_0(0)) AND (NOT and_dcpl_717))
      OR and_dcpl_741;
  acc_9_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_24_nl
      & COMP_LOOP_mux1h_598_nl & COMP_LOOP_or_83_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_mux_22_nl
      & COMP_LOOP_COMP_LOOP_or_25_nl & '1'), 7), 8), 8));
  z_out_9 <= acc_9_nl(7 DOWNTO 1);
  nor_1463_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(6)));
  nor_1464_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(2))
      OR (fsm_output(3)) OR nand_257_cse);
  mux_3958_nl <= MUX_s_1_2_2(nor_1463_nl, nor_1464_nl, fsm_output(1));
  nor_1465_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(6)));
  mux_3957_nl <= MUX_s_1_2_2(mux_3958_nl, nor_1465_nl, fsm_output(4));
  nor_1466_nl <= NOT((fsm_output(1)) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (fsm_output(3)) OR nand_257_cse);
  nor_1467_nl <= NOT((fsm_output(5)) OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT
      (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(6)));
  nor_1468_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (fsm_output(3)) OR (fsm_output(8)) OR (NOT (fsm_output(6))));
  mux_3960_nl <= MUX_s_1_2_2(nor_1467_nl, nor_1468_nl, fsm_output(1));
  mux_3959_nl <= MUX_s_1_2_2(nor_1466_nl, mux_3960_nl, fsm_output(4));
  mux_3956_nl <= MUX_s_1_2_2(mux_3957_nl, mux_3959_nl, fsm_output(7));
  nor_1469_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(6)));
  nor_1470_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR (fsm_output(2)) OR (NOT((fsm_output(3)) AND (fsm_output(8)) AND (fsm_output(6)))));
  mux_3962_nl <= MUX_s_1_2_2(nor_1469_nl, nor_1470_nl, fsm_output(4));
  nor_1471_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)) OR (fsm_output(9))
      OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR nand_257_cse);
  or_3612_nl <= (NOT (fsm_output(9))) OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(8))
      OR (fsm_output(6));
  or_3613_nl <= (fsm_output(9)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))
      OR (fsm_output(8)) OR (NOT (fsm_output(6)));
  mux_3964_nl <= MUX_s_1_2_2(or_3612_nl, or_3613_nl, fsm_output(5));
  nor_1472_nl <= NOT((fsm_output(1)) OR mux_3964_nl);
  mux_3963_nl <= MUX_s_1_2_2(nor_1471_nl, nor_1472_nl, fsm_output(4));
  mux_3961_nl <= MUX_s_1_2_2(mux_3962_nl, mux_3963_nl, fsm_output(7));
  mux_3955_nl <= MUX_s_1_2_2(mux_3956_nl, mux_3961_nl, fsm_output(0));
  nor_1473_nl <= NOT((fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(2)))
      OR (fsm_output(3)) OR nand_257_cse);
  nor_1474_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(9))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(3))) OR (fsm_output(8)) OR (fsm_output(6)));
  mux_3967_nl <= MUX_s_1_2_2(nor_1473_nl, nor_1474_nl, fsm_output(1));
  and_1286_nl <= (fsm_output(4)) AND mux_3967_nl;
  nor_1475_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(1))) OR (fsm_output(5))
      OR (fsm_output(9)) OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (fsm_output(8))
      OR (fsm_output(6)));
  mux_3966_nl <= MUX_s_1_2_2(and_1286_nl, nor_1475_nl, fsm_output(7));
  nor_1476_nl <= NOT((fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR (NOT (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(8))
      OR (fsm_output(6)));
  and_1287_nl <= (fsm_output(1)) AND (fsm_output(5)) AND (NOT (fsm_output(9))) AND
      (fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(8))) AND (fsm_output(6));
  nor_1477_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (fsm_output(2)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(8))) OR (fsm_output(6)));
  mux_3969_nl <= MUX_s_1_2_2(and_1287_nl, nor_1477_nl, fsm_output(4));
  mux_3968_nl <= MUX_s_1_2_2(nor_1476_nl, mux_3969_nl, fsm_output(7));
  mux_3965_nl <= MUX_s_1_2_2(mux_3966_nl, mux_3968_nl, fsm_output(0));
  mux_3954_nl <= MUX_s_1_2_2(mux_3955_nl, mux_3965_nl, fsm_output(10));
  modExp_while_if_mux_1_nl <= MUX_v_64_2_2(modExp_result_sva, COMP_LOOP_10_mul_mut,
      mux_3954_nl);
  z_out_10 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(modExp_while_if_mux_1_nl)
      * SIGNED(COMP_LOOP_10_mul_mut)), 64));
END v43;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_0_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_wea : OUT STD_LOGIC;
    vec_rsc_0_0_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_1_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_wea : OUT STD_LOGIC;
    vec_rsc_0_1_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_2_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_wea : OUT STD_LOGIC;
    vec_rsc_0_2_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_3_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_wea : OUT STD_LOGIC;
    vec_rsc_0_3_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_4_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_wea : OUT STD_LOGIC;
    vec_rsc_0_4_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_5_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_wea : OUT STD_LOGIC;
    vec_rsc_0_5_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_6_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_wea : OUT STD_LOGIC;
    vec_rsc_0_6_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_7_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_wea : OUT STD_LOGIC;
    vec_rsc_0_7_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_8_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_wea : OUT STD_LOGIC;
    vec_rsc_0_8_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_9_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_wea : OUT STD_LOGIC;
    vec_rsc_0_9_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_10_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_wea : OUT STD_LOGIC;
    vec_rsc_0_10_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_11_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_wea : OUT STD_LOGIC;
    vec_rsc_0_11_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_12_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_wea : OUT STD_LOGIC;
    vec_rsc_0_12_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_13_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_wea : OUT STD_LOGIC;
    vec_rsc_0_13_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_14_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_wea : OUT STD_LOGIC;
    vec_rsc_0_14_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    vec_rsc_0_15_da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_wea : OUT STD_LOGIC;
    vec_rsc_0_15_qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC
  );
END inPlaceNTT_DIT;

ARCHITECTURE v43 OF inPlaceNTT_DIT IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_adra_d_iff : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_wea_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_wea_d_iff : STD_LOGIC;

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_8_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_9_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_10_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_11_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_12_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_13_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_14_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_15_i_qa : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_da : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_adra : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      r_rsc_triosy_lz : OUT STD_LOGIC;
      vec_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      vec_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
      vec_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_r_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff : STD_LOGIC_VECTOR (7
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO
      0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_0_i_qa,
      wea => vec_rsc_0_0_wea,
      da => vec_rsc_0_0_i_da,
      adra => vec_rsc_0_0_i_adra,
      adra_d => vec_rsc_0_0_i_adra_d,
      da_d => vec_rsc_0_0_i_da_d,
      qa_d => vec_rsc_0_0_i_qa_d_1,
      wea_d => vec_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_wea_d_iff
    );
  vec_rsc_0_0_i_qa <= vec_rsc_0_0_qa;
  vec_rsc_0_0_da <= vec_rsc_0_0_i_da;
  vec_rsc_0_0_adra <= vec_rsc_0_0_i_adra;
  vec_rsc_0_0_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_0_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d_1;

  vec_rsc_0_1_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_1_i_qa,
      wea => vec_rsc_0_1_wea,
      da => vec_rsc_0_1_i_da,
      adra => vec_rsc_0_1_i_adra,
      adra_d => vec_rsc_0_1_i_adra_d,
      da_d => vec_rsc_0_1_i_da_d,
      qa_d => vec_rsc_0_1_i_qa_d_1,
      wea_d => vec_rsc_0_1_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_wea_d_iff
    );
  vec_rsc_0_1_i_qa <= vec_rsc_0_1_qa;
  vec_rsc_0_1_da <= vec_rsc_0_1_i_da;
  vec_rsc_0_1_adra <= vec_rsc_0_1_i_adra;
  vec_rsc_0_1_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_1_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d_1;

  vec_rsc_0_2_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_2_i_qa,
      wea => vec_rsc_0_2_wea,
      da => vec_rsc_0_2_i_da,
      adra => vec_rsc_0_2_i_adra,
      adra_d => vec_rsc_0_2_i_adra_d,
      da_d => vec_rsc_0_2_i_da_d,
      qa_d => vec_rsc_0_2_i_qa_d_1,
      wea_d => vec_rsc_0_2_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_wea_d_iff
    );
  vec_rsc_0_2_i_qa <= vec_rsc_0_2_qa;
  vec_rsc_0_2_da <= vec_rsc_0_2_i_da;
  vec_rsc_0_2_adra <= vec_rsc_0_2_i_adra;
  vec_rsc_0_2_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_2_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d_1;

  vec_rsc_0_3_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_3_i_qa,
      wea => vec_rsc_0_3_wea,
      da => vec_rsc_0_3_i_da,
      adra => vec_rsc_0_3_i_adra,
      adra_d => vec_rsc_0_3_i_adra_d,
      da_d => vec_rsc_0_3_i_da_d,
      qa_d => vec_rsc_0_3_i_qa_d_1,
      wea_d => vec_rsc_0_3_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_wea_d_iff
    );
  vec_rsc_0_3_i_qa <= vec_rsc_0_3_qa;
  vec_rsc_0_3_da <= vec_rsc_0_3_i_da;
  vec_rsc_0_3_adra <= vec_rsc_0_3_i_adra;
  vec_rsc_0_3_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_3_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d_1;

  vec_rsc_0_4_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_4_i_qa,
      wea => vec_rsc_0_4_wea,
      da => vec_rsc_0_4_i_da,
      adra => vec_rsc_0_4_i_adra,
      adra_d => vec_rsc_0_4_i_adra_d,
      da_d => vec_rsc_0_4_i_da_d,
      qa_d => vec_rsc_0_4_i_qa_d_1,
      wea_d => vec_rsc_0_4_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_wea_d_iff
    );
  vec_rsc_0_4_i_qa <= vec_rsc_0_4_qa;
  vec_rsc_0_4_da <= vec_rsc_0_4_i_da;
  vec_rsc_0_4_adra <= vec_rsc_0_4_i_adra;
  vec_rsc_0_4_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_4_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d_1;

  vec_rsc_0_5_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_5_i_qa,
      wea => vec_rsc_0_5_wea,
      da => vec_rsc_0_5_i_da,
      adra => vec_rsc_0_5_i_adra,
      adra_d => vec_rsc_0_5_i_adra_d,
      da_d => vec_rsc_0_5_i_da_d,
      qa_d => vec_rsc_0_5_i_qa_d_1,
      wea_d => vec_rsc_0_5_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_wea_d_iff
    );
  vec_rsc_0_5_i_qa <= vec_rsc_0_5_qa;
  vec_rsc_0_5_da <= vec_rsc_0_5_i_da;
  vec_rsc_0_5_adra <= vec_rsc_0_5_i_adra;
  vec_rsc_0_5_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_5_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d_1;

  vec_rsc_0_6_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_6_i_qa,
      wea => vec_rsc_0_6_wea,
      da => vec_rsc_0_6_i_da,
      adra => vec_rsc_0_6_i_adra,
      adra_d => vec_rsc_0_6_i_adra_d,
      da_d => vec_rsc_0_6_i_da_d,
      qa_d => vec_rsc_0_6_i_qa_d_1,
      wea_d => vec_rsc_0_6_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_wea_d_iff
    );
  vec_rsc_0_6_i_qa <= vec_rsc_0_6_qa;
  vec_rsc_0_6_da <= vec_rsc_0_6_i_da;
  vec_rsc_0_6_adra <= vec_rsc_0_6_i_adra;
  vec_rsc_0_6_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_6_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d_1;

  vec_rsc_0_7_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_7_i_qa,
      wea => vec_rsc_0_7_wea,
      da => vec_rsc_0_7_i_da,
      adra => vec_rsc_0_7_i_adra,
      adra_d => vec_rsc_0_7_i_adra_d,
      da_d => vec_rsc_0_7_i_da_d,
      qa_d => vec_rsc_0_7_i_qa_d_1,
      wea_d => vec_rsc_0_7_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_wea_d_iff
    );
  vec_rsc_0_7_i_qa <= vec_rsc_0_7_qa;
  vec_rsc_0_7_da <= vec_rsc_0_7_i_da;
  vec_rsc_0_7_adra <= vec_rsc_0_7_i_adra;
  vec_rsc_0_7_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_7_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d_1;

  vec_rsc_0_8_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_8_i_qa,
      wea => vec_rsc_0_8_wea,
      da => vec_rsc_0_8_i_da,
      adra => vec_rsc_0_8_i_adra,
      adra_d => vec_rsc_0_8_i_adra_d,
      da_d => vec_rsc_0_8_i_da_d,
      qa_d => vec_rsc_0_8_i_qa_d_1,
      wea_d => vec_rsc_0_8_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_8_i_wea_d_iff
    );
  vec_rsc_0_8_i_qa <= vec_rsc_0_8_qa;
  vec_rsc_0_8_da <= vec_rsc_0_8_i_da;
  vec_rsc_0_8_adra <= vec_rsc_0_8_i_adra;
  vec_rsc_0_8_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_8_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_8_i_qa_d <= vec_rsc_0_8_i_qa_d_1;

  vec_rsc_0_9_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_9_i_qa,
      wea => vec_rsc_0_9_wea,
      da => vec_rsc_0_9_i_da,
      adra => vec_rsc_0_9_i_adra,
      adra_d => vec_rsc_0_9_i_adra_d,
      da_d => vec_rsc_0_9_i_da_d,
      qa_d => vec_rsc_0_9_i_qa_d_1,
      wea_d => vec_rsc_0_9_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_9_i_wea_d_iff
    );
  vec_rsc_0_9_i_qa <= vec_rsc_0_9_qa;
  vec_rsc_0_9_da <= vec_rsc_0_9_i_da;
  vec_rsc_0_9_adra <= vec_rsc_0_9_i_adra;
  vec_rsc_0_9_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_9_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_9_i_qa_d <= vec_rsc_0_9_i_qa_d_1;

  vec_rsc_0_10_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_10_i_qa,
      wea => vec_rsc_0_10_wea,
      da => vec_rsc_0_10_i_da,
      adra => vec_rsc_0_10_i_adra,
      adra_d => vec_rsc_0_10_i_adra_d,
      da_d => vec_rsc_0_10_i_da_d,
      qa_d => vec_rsc_0_10_i_qa_d_1,
      wea_d => vec_rsc_0_10_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_10_i_wea_d_iff
    );
  vec_rsc_0_10_i_qa <= vec_rsc_0_10_qa;
  vec_rsc_0_10_da <= vec_rsc_0_10_i_da;
  vec_rsc_0_10_adra <= vec_rsc_0_10_i_adra;
  vec_rsc_0_10_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_10_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_10_i_qa_d <= vec_rsc_0_10_i_qa_d_1;

  vec_rsc_0_11_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_11_i_qa,
      wea => vec_rsc_0_11_wea,
      da => vec_rsc_0_11_i_da,
      adra => vec_rsc_0_11_i_adra,
      adra_d => vec_rsc_0_11_i_adra_d,
      da_d => vec_rsc_0_11_i_da_d,
      qa_d => vec_rsc_0_11_i_qa_d_1,
      wea_d => vec_rsc_0_11_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_11_i_wea_d_iff
    );
  vec_rsc_0_11_i_qa <= vec_rsc_0_11_qa;
  vec_rsc_0_11_da <= vec_rsc_0_11_i_da;
  vec_rsc_0_11_adra <= vec_rsc_0_11_i_adra;
  vec_rsc_0_11_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_11_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_11_i_qa_d <= vec_rsc_0_11_i_qa_d_1;

  vec_rsc_0_12_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_12_i_qa,
      wea => vec_rsc_0_12_wea,
      da => vec_rsc_0_12_i_da,
      adra => vec_rsc_0_12_i_adra,
      adra_d => vec_rsc_0_12_i_adra_d,
      da_d => vec_rsc_0_12_i_da_d,
      qa_d => vec_rsc_0_12_i_qa_d_1,
      wea_d => vec_rsc_0_12_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_12_i_wea_d_iff
    );
  vec_rsc_0_12_i_qa <= vec_rsc_0_12_qa;
  vec_rsc_0_12_da <= vec_rsc_0_12_i_da;
  vec_rsc_0_12_adra <= vec_rsc_0_12_i_adra;
  vec_rsc_0_12_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_12_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_12_i_qa_d <= vec_rsc_0_12_i_qa_d_1;

  vec_rsc_0_13_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_13_i_qa,
      wea => vec_rsc_0_13_wea,
      da => vec_rsc_0_13_i_da,
      adra => vec_rsc_0_13_i_adra,
      adra_d => vec_rsc_0_13_i_adra_d,
      da_d => vec_rsc_0_13_i_da_d,
      qa_d => vec_rsc_0_13_i_qa_d_1,
      wea_d => vec_rsc_0_13_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_13_i_wea_d_iff
    );
  vec_rsc_0_13_i_qa <= vec_rsc_0_13_qa;
  vec_rsc_0_13_da <= vec_rsc_0_13_i_da;
  vec_rsc_0_13_adra <= vec_rsc_0_13_i_adra;
  vec_rsc_0_13_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_13_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_13_i_qa_d <= vec_rsc_0_13_i_qa_d_1;

  vec_rsc_0_14_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_14_i_qa,
      wea => vec_rsc_0_14_wea,
      da => vec_rsc_0_14_i_da,
      adra => vec_rsc_0_14_i_adra,
      adra_d => vec_rsc_0_14_i_adra_d,
      da_d => vec_rsc_0_14_i_da_d,
      qa_d => vec_rsc_0_14_i_qa_d_1,
      wea_d => vec_rsc_0_14_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_14_i_wea_d_iff
    );
  vec_rsc_0_14_i_qa <= vec_rsc_0_14_qa;
  vec_rsc_0_14_da <= vec_rsc_0_14_i_da;
  vec_rsc_0_14_adra <= vec_rsc_0_14_i_adra;
  vec_rsc_0_14_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_14_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_14_i_qa_d <= vec_rsc_0_14_i_qa_d_1;

  vec_rsc_0_15_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    PORT MAP(
      qa => vec_rsc_0_15_i_qa,
      wea => vec_rsc_0_15_wea,
      da => vec_rsc_0_15_i_da,
      adra => vec_rsc_0_15_i_adra,
      adra_d => vec_rsc_0_15_i_adra_d,
      da_d => vec_rsc_0_15_i_da_d,
      qa_d => vec_rsc_0_15_i_qa_d_1,
      wea_d => vec_rsc_0_15_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => vec_rsc_0_15_i_wea_d_iff
    );
  vec_rsc_0_15_i_qa <= vec_rsc_0_15_qa;
  vec_rsc_0_15_da <= vec_rsc_0_15_i_da;
  vec_rsc_0_15_adra <= vec_rsc_0_15_i_adra;
  vec_rsc_0_15_i_adra_d <= vec_rsc_0_0_i_adra_d_iff;
  vec_rsc_0_15_i_da_d <= vec_rsc_0_0_i_da_d_iff;
  vec_rsc_0_15_i_qa_d <= vec_rsc_0_15_i_qa_d_1;

  inPlaceNTT_DIT_core_inst : inPlaceNTT_DIT_core
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      vec_rsc_triosy_0_8_lz => vec_rsc_triosy_0_8_lz,
      vec_rsc_triosy_0_9_lz => vec_rsc_triosy_0_9_lz,
      vec_rsc_triosy_0_10_lz => vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz => vec_rsc_triosy_0_11_lz,
      vec_rsc_triosy_0_12_lz => vec_rsc_triosy_0_12_lz,
      vec_rsc_triosy_0_13_lz => vec_rsc_triosy_0_13_lz,
      vec_rsc_triosy_0_14_lz => vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz => vec_rsc_triosy_0_15_lz,
      p_rsc_dat => inPlaceNTT_DIT_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_dat => inPlaceNTT_DIT_core_inst_r_rsc_dat,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d,
      vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d,
      vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d,
      vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d,
      vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d,
      vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_8_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_qa_d,
      vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_qa_d,
      vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_10_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_qa_d,
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_11_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_qa_d,
      vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_qa_d,
      vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_13_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_qa_d,
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_14_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_qa_d,
      vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_qa_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_qa_d,
      vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_adra_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff,
      vec_rsc_0_0_i_wea_d_pff => vec_rsc_0_0_i_wea_d_iff,
      vec_rsc_0_1_i_wea_d_pff => vec_rsc_0_1_i_wea_d_iff,
      vec_rsc_0_2_i_wea_d_pff => vec_rsc_0_2_i_wea_d_iff,
      vec_rsc_0_3_i_wea_d_pff => vec_rsc_0_3_i_wea_d_iff,
      vec_rsc_0_4_i_wea_d_pff => vec_rsc_0_4_i_wea_d_iff,
      vec_rsc_0_5_i_wea_d_pff => vec_rsc_0_5_i_wea_d_iff,
      vec_rsc_0_6_i_wea_d_pff => vec_rsc_0_6_i_wea_d_iff,
      vec_rsc_0_7_i_wea_d_pff => vec_rsc_0_7_i_wea_d_iff,
      vec_rsc_0_8_i_wea_d_pff => vec_rsc_0_8_i_wea_d_iff,
      vec_rsc_0_9_i_wea_d_pff => vec_rsc_0_9_i_wea_d_iff,
      vec_rsc_0_10_i_wea_d_pff => vec_rsc_0_10_i_wea_d_iff,
      vec_rsc_0_11_i_wea_d_pff => vec_rsc_0_11_i_wea_d_iff,
      vec_rsc_0_12_i_wea_d_pff => vec_rsc_0_12_i_wea_d_iff,
      vec_rsc_0_13_i_wea_d_pff => vec_rsc_0_13_i_wea_d_iff,
      vec_rsc_0_14_i_wea_d_pff => vec_rsc_0_14_i_wea_d_iff,
      vec_rsc_0_15_i_wea_d_pff => vec_rsc_0_15_i_wea_d_iff
    );
  inPlaceNTT_DIT_core_inst_p_rsc_dat <= p_rsc_dat;
  inPlaceNTT_DIT_core_inst_r_rsc_dat <= r_rsc_dat;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_qa_d <= vec_rsc_0_0_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_qa_d <= vec_rsc_0_1_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_qa_d <= vec_rsc_0_2_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_qa_d <= vec_rsc_0_3_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_qa_d <= vec_rsc_0_4_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_qa_d <= vec_rsc_0_5_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_qa_d <= vec_rsc_0_6_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_qa_d <= vec_rsc_0_7_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_qa_d <= vec_rsc_0_8_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_qa_d <= vec_rsc_0_9_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_qa_d <= vec_rsc_0_10_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_qa_d <= vec_rsc_0_11_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_qa_d <= vec_rsc_0_12_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_qa_d <= vec_rsc_0_13_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_qa_d <= vec_rsc_0_14_i_qa_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_qa_d <= vec_rsc_0_15_i_qa_d;
  vec_rsc_0_0_i_adra_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_adra_d_pff;
  vec_rsc_0_0_i_da_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_da_d_pff;

END v43;



