
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Wed May 19 22:57:49 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_8_tr0, modExp_while_C_38_tr0, VEC_LOOP_1_COMP_LOOP_C_1_tr0,
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38_tr0, VEC_LOOP_1_COMP_LOOP_C_62_tr0,
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38_tr0, VEC_LOOP_1_COMP_LOOP_C_124_tr0,
      VEC_LOOP_C_0_tr0, VEC_LOOP_2_COMP_LOOP_C_1_tr0, VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38_tr0,
      VEC_LOOP_2_COMP_LOOP_C_62_tr0, VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38_tr0,
      VEC_LOOP_2_COMP_LOOP_C_124_tr0, VEC_LOOP_C_1_tr0, STAGE_LOOP_C_9_tr0
);
  input clk;
  input rst;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input STAGE_LOOP_C_8_tr0;
  input modExp_while_C_38_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_1_tr0;
  input VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_62_tr0;
  input VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_124_tr0;
  input VEC_LOOP_C_0_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_1_tr0;
  input VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_62_tr0;
  input VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_124_tr0;
  input VEC_LOOP_C_1_tr0;
  input STAGE_LOOP_C_9_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 9'd0,
    STAGE_LOOP_C_0 = 9'd1,
    STAGE_LOOP_C_1 = 9'd2,
    STAGE_LOOP_C_2 = 9'd3,
    STAGE_LOOP_C_3 = 9'd4,
    STAGE_LOOP_C_4 = 9'd5,
    STAGE_LOOP_C_5 = 9'd6,
    STAGE_LOOP_C_6 = 9'd7,
    STAGE_LOOP_C_7 = 9'd8,
    STAGE_LOOP_C_8 = 9'd9,
    modExp_while_C_0 = 9'd10,
    modExp_while_C_1 = 9'd11,
    modExp_while_C_2 = 9'd12,
    modExp_while_C_3 = 9'd13,
    modExp_while_C_4 = 9'd14,
    modExp_while_C_5 = 9'd15,
    modExp_while_C_6 = 9'd16,
    modExp_while_C_7 = 9'd17,
    modExp_while_C_8 = 9'd18,
    modExp_while_C_9 = 9'd19,
    modExp_while_C_10 = 9'd20,
    modExp_while_C_11 = 9'd21,
    modExp_while_C_12 = 9'd22,
    modExp_while_C_13 = 9'd23,
    modExp_while_C_14 = 9'd24,
    modExp_while_C_15 = 9'd25,
    modExp_while_C_16 = 9'd26,
    modExp_while_C_17 = 9'd27,
    modExp_while_C_18 = 9'd28,
    modExp_while_C_19 = 9'd29,
    modExp_while_C_20 = 9'd30,
    modExp_while_C_21 = 9'd31,
    modExp_while_C_22 = 9'd32,
    modExp_while_C_23 = 9'd33,
    modExp_while_C_24 = 9'd34,
    modExp_while_C_25 = 9'd35,
    modExp_while_C_26 = 9'd36,
    modExp_while_C_27 = 9'd37,
    modExp_while_C_28 = 9'd38,
    modExp_while_C_29 = 9'd39,
    modExp_while_C_30 = 9'd40,
    modExp_while_C_31 = 9'd41,
    modExp_while_C_32 = 9'd42,
    modExp_while_C_33 = 9'd43,
    modExp_while_C_34 = 9'd44,
    modExp_while_C_35 = 9'd45,
    modExp_while_C_36 = 9'd46,
    modExp_while_C_37 = 9'd47,
    modExp_while_C_38 = 9'd48,
    VEC_LOOP_1_COMP_LOOP_C_0 = 9'd49,
    VEC_LOOP_1_COMP_LOOP_C_1 = 9'd50,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0 = 9'd51,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1 = 9'd52,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2 = 9'd53,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3 = 9'd54,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4 = 9'd55,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5 = 9'd56,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6 = 9'd57,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7 = 9'd58,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8 = 9'd59,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9 = 9'd60,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10 = 9'd61,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11 = 9'd62,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12 = 9'd63,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13 = 9'd64,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14 = 9'd65,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15 = 9'd66,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16 = 9'd67,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17 = 9'd68,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18 = 9'd69,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19 = 9'd70,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20 = 9'd71,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21 = 9'd72,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22 = 9'd73,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23 = 9'd74,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24 = 9'd75,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_25 = 9'd76,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_26 = 9'd77,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_27 = 9'd78,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_28 = 9'd79,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_29 = 9'd80,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_30 = 9'd81,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_31 = 9'd82,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_32 = 9'd83,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_33 = 9'd84,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_34 = 9'd85,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_35 = 9'd86,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_36 = 9'd87,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_37 = 9'd88,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38 = 9'd89,
    VEC_LOOP_1_COMP_LOOP_C_2 = 9'd90,
    VEC_LOOP_1_COMP_LOOP_C_3 = 9'd91,
    VEC_LOOP_1_COMP_LOOP_C_4 = 9'd92,
    VEC_LOOP_1_COMP_LOOP_C_5 = 9'd93,
    VEC_LOOP_1_COMP_LOOP_C_6 = 9'd94,
    VEC_LOOP_1_COMP_LOOP_C_7 = 9'd95,
    VEC_LOOP_1_COMP_LOOP_C_8 = 9'd96,
    VEC_LOOP_1_COMP_LOOP_C_9 = 9'd97,
    VEC_LOOP_1_COMP_LOOP_C_10 = 9'd98,
    VEC_LOOP_1_COMP_LOOP_C_11 = 9'd99,
    VEC_LOOP_1_COMP_LOOP_C_12 = 9'd100,
    VEC_LOOP_1_COMP_LOOP_C_13 = 9'd101,
    VEC_LOOP_1_COMP_LOOP_C_14 = 9'd102,
    VEC_LOOP_1_COMP_LOOP_C_15 = 9'd103,
    VEC_LOOP_1_COMP_LOOP_C_16 = 9'd104,
    VEC_LOOP_1_COMP_LOOP_C_17 = 9'd105,
    VEC_LOOP_1_COMP_LOOP_C_18 = 9'd106,
    VEC_LOOP_1_COMP_LOOP_C_19 = 9'd107,
    VEC_LOOP_1_COMP_LOOP_C_20 = 9'd108,
    VEC_LOOP_1_COMP_LOOP_C_21 = 9'd109,
    VEC_LOOP_1_COMP_LOOP_C_22 = 9'd110,
    VEC_LOOP_1_COMP_LOOP_C_23 = 9'd111,
    VEC_LOOP_1_COMP_LOOP_C_24 = 9'd112,
    VEC_LOOP_1_COMP_LOOP_C_25 = 9'd113,
    VEC_LOOP_1_COMP_LOOP_C_26 = 9'd114,
    VEC_LOOP_1_COMP_LOOP_C_27 = 9'd115,
    VEC_LOOP_1_COMP_LOOP_C_28 = 9'd116,
    VEC_LOOP_1_COMP_LOOP_C_29 = 9'd117,
    VEC_LOOP_1_COMP_LOOP_C_30 = 9'd118,
    VEC_LOOP_1_COMP_LOOP_C_31 = 9'd119,
    VEC_LOOP_1_COMP_LOOP_C_32 = 9'd120,
    VEC_LOOP_1_COMP_LOOP_C_33 = 9'd121,
    VEC_LOOP_1_COMP_LOOP_C_34 = 9'd122,
    VEC_LOOP_1_COMP_LOOP_C_35 = 9'd123,
    VEC_LOOP_1_COMP_LOOP_C_36 = 9'd124,
    VEC_LOOP_1_COMP_LOOP_C_37 = 9'd125,
    VEC_LOOP_1_COMP_LOOP_C_38 = 9'd126,
    VEC_LOOP_1_COMP_LOOP_C_39 = 9'd127,
    VEC_LOOP_1_COMP_LOOP_C_40 = 9'd128,
    VEC_LOOP_1_COMP_LOOP_C_41 = 9'd129,
    VEC_LOOP_1_COMP_LOOP_C_42 = 9'd130,
    VEC_LOOP_1_COMP_LOOP_C_43 = 9'd131,
    VEC_LOOP_1_COMP_LOOP_C_44 = 9'd132,
    VEC_LOOP_1_COMP_LOOP_C_45 = 9'd133,
    VEC_LOOP_1_COMP_LOOP_C_46 = 9'd134,
    VEC_LOOP_1_COMP_LOOP_C_47 = 9'd135,
    VEC_LOOP_1_COMP_LOOP_C_48 = 9'd136,
    VEC_LOOP_1_COMP_LOOP_C_49 = 9'd137,
    VEC_LOOP_1_COMP_LOOP_C_50 = 9'd138,
    VEC_LOOP_1_COMP_LOOP_C_51 = 9'd139,
    VEC_LOOP_1_COMP_LOOP_C_52 = 9'd140,
    VEC_LOOP_1_COMP_LOOP_C_53 = 9'd141,
    VEC_LOOP_1_COMP_LOOP_C_54 = 9'd142,
    VEC_LOOP_1_COMP_LOOP_C_55 = 9'd143,
    VEC_LOOP_1_COMP_LOOP_C_56 = 9'd144,
    VEC_LOOP_1_COMP_LOOP_C_57 = 9'd145,
    VEC_LOOP_1_COMP_LOOP_C_58 = 9'd146,
    VEC_LOOP_1_COMP_LOOP_C_59 = 9'd147,
    VEC_LOOP_1_COMP_LOOP_C_60 = 9'd148,
    VEC_LOOP_1_COMP_LOOP_C_61 = 9'd149,
    VEC_LOOP_1_COMP_LOOP_C_62 = 9'd150,
    VEC_LOOP_1_COMP_LOOP_C_63 = 9'd151,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0 = 9'd152,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1 = 9'd153,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2 = 9'd154,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3 = 9'd155,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4 = 9'd156,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5 = 9'd157,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6 = 9'd158,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7 = 9'd159,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8 = 9'd160,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9 = 9'd161,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10 = 9'd162,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11 = 9'd163,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12 = 9'd164,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13 = 9'd165,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14 = 9'd166,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15 = 9'd167,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16 = 9'd168,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17 = 9'd169,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18 = 9'd170,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19 = 9'd171,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20 = 9'd172,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21 = 9'd173,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22 = 9'd174,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23 = 9'd175,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24 = 9'd176,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_25 = 9'd177,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_26 = 9'd178,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_27 = 9'd179,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_28 = 9'd180,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_29 = 9'd181,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_30 = 9'd182,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_31 = 9'd183,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_32 = 9'd184,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_33 = 9'd185,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_34 = 9'd186,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_35 = 9'd187,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_36 = 9'd188,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_37 = 9'd189,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38 = 9'd190,
    VEC_LOOP_1_COMP_LOOP_C_64 = 9'd191,
    VEC_LOOP_1_COMP_LOOP_C_65 = 9'd192,
    VEC_LOOP_1_COMP_LOOP_C_66 = 9'd193,
    VEC_LOOP_1_COMP_LOOP_C_67 = 9'd194,
    VEC_LOOP_1_COMP_LOOP_C_68 = 9'd195,
    VEC_LOOP_1_COMP_LOOP_C_69 = 9'd196,
    VEC_LOOP_1_COMP_LOOP_C_70 = 9'd197,
    VEC_LOOP_1_COMP_LOOP_C_71 = 9'd198,
    VEC_LOOP_1_COMP_LOOP_C_72 = 9'd199,
    VEC_LOOP_1_COMP_LOOP_C_73 = 9'd200,
    VEC_LOOP_1_COMP_LOOP_C_74 = 9'd201,
    VEC_LOOP_1_COMP_LOOP_C_75 = 9'd202,
    VEC_LOOP_1_COMP_LOOP_C_76 = 9'd203,
    VEC_LOOP_1_COMP_LOOP_C_77 = 9'd204,
    VEC_LOOP_1_COMP_LOOP_C_78 = 9'd205,
    VEC_LOOP_1_COMP_LOOP_C_79 = 9'd206,
    VEC_LOOP_1_COMP_LOOP_C_80 = 9'd207,
    VEC_LOOP_1_COMP_LOOP_C_81 = 9'd208,
    VEC_LOOP_1_COMP_LOOP_C_82 = 9'd209,
    VEC_LOOP_1_COMP_LOOP_C_83 = 9'd210,
    VEC_LOOP_1_COMP_LOOP_C_84 = 9'd211,
    VEC_LOOP_1_COMP_LOOP_C_85 = 9'd212,
    VEC_LOOP_1_COMP_LOOP_C_86 = 9'd213,
    VEC_LOOP_1_COMP_LOOP_C_87 = 9'd214,
    VEC_LOOP_1_COMP_LOOP_C_88 = 9'd215,
    VEC_LOOP_1_COMP_LOOP_C_89 = 9'd216,
    VEC_LOOP_1_COMP_LOOP_C_90 = 9'd217,
    VEC_LOOP_1_COMP_LOOP_C_91 = 9'd218,
    VEC_LOOP_1_COMP_LOOP_C_92 = 9'd219,
    VEC_LOOP_1_COMP_LOOP_C_93 = 9'd220,
    VEC_LOOP_1_COMP_LOOP_C_94 = 9'd221,
    VEC_LOOP_1_COMP_LOOP_C_95 = 9'd222,
    VEC_LOOP_1_COMP_LOOP_C_96 = 9'd223,
    VEC_LOOP_1_COMP_LOOP_C_97 = 9'd224,
    VEC_LOOP_1_COMP_LOOP_C_98 = 9'd225,
    VEC_LOOP_1_COMP_LOOP_C_99 = 9'd226,
    VEC_LOOP_1_COMP_LOOP_C_100 = 9'd227,
    VEC_LOOP_1_COMP_LOOP_C_101 = 9'd228,
    VEC_LOOP_1_COMP_LOOP_C_102 = 9'd229,
    VEC_LOOP_1_COMP_LOOP_C_103 = 9'd230,
    VEC_LOOP_1_COMP_LOOP_C_104 = 9'd231,
    VEC_LOOP_1_COMP_LOOP_C_105 = 9'd232,
    VEC_LOOP_1_COMP_LOOP_C_106 = 9'd233,
    VEC_LOOP_1_COMP_LOOP_C_107 = 9'd234,
    VEC_LOOP_1_COMP_LOOP_C_108 = 9'd235,
    VEC_LOOP_1_COMP_LOOP_C_109 = 9'd236,
    VEC_LOOP_1_COMP_LOOP_C_110 = 9'd237,
    VEC_LOOP_1_COMP_LOOP_C_111 = 9'd238,
    VEC_LOOP_1_COMP_LOOP_C_112 = 9'd239,
    VEC_LOOP_1_COMP_LOOP_C_113 = 9'd240,
    VEC_LOOP_1_COMP_LOOP_C_114 = 9'd241,
    VEC_LOOP_1_COMP_LOOP_C_115 = 9'd242,
    VEC_LOOP_1_COMP_LOOP_C_116 = 9'd243,
    VEC_LOOP_1_COMP_LOOP_C_117 = 9'd244,
    VEC_LOOP_1_COMP_LOOP_C_118 = 9'd245,
    VEC_LOOP_1_COMP_LOOP_C_119 = 9'd246,
    VEC_LOOP_1_COMP_LOOP_C_120 = 9'd247,
    VEC_LOOP_1_COMP_LOOP_C_121 = 9'd248,
    VEC_LOOP_1_COMP_LOOP_C_122 = 9'd249,
    VEC_LOOP_1_COMP_LOOP_C_123 = 9'd250,
    VEC_LOOP_1_COMP_LOOP_C_124 = 9'd251,
    VEC_LOOP_C_0 = 9'd252,
    VEC_LOOP_2_COMP_LOOP_C_0 = 9'd253,
    VEC_LOOP_2_COMP_LOOP_C_1 = 9'd254,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0 = 9'd255,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1 = 9'd256,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2 = 9'd257,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3 = 9'd258,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4 = 9'd259,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5 = 9'd260,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6 = 9'd261,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7 = 9'd262,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8 = 9'd263,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9 = 9'd264,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10 = 9'd265,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11 = 9'd266,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12 = 9'd267,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13 = 9'd268,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14 = 9'd269,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15 = 9'd270,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16 = 9'd271,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17 = 9'd272,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18 = 9'd273,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19 = 9'd274,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20 = 9'd275,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21 = 9'd276,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22 = 9'd277,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23 = 9'd278,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24 = 9'd279,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_25 = 9'd280,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_26 = 9'd281,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_27 = 9'd282,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_28 = 9'd283,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_29 = 9'd284,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_30 = 9'd285,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_31 = 9'd286,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_32 = 9'd287,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_33 = 9'd288,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_34 = 9'd289,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_35 = 9'd290,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_36 = 9'd291,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_37 = 9'd292,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38 = 9'd293,
    VEC_LOOP_2_COMP_LOOP_C_2 = 9'd294,
    VEC_LOOP_2_COMP_LOOP_C_3 = 9'd295,
    VEC_LOOP_2_COMP_LOOP_C_4 = 9'd296,
    VEC_LOOP_2_COMP_LOOP_C_5 = 9'd297,
    VEC_LOOP_2_COMP_LOOP_C_6 = 9'd298,
    VEC_LOOP_2_COMP_LOOP_C_7 = 9'd299,
    VEC_LOOP_2_COMP_LOOP_C_8 = 9'd300,
    VEC_LOOP_2_COMP_LOOP_C_9 = 9'd301,
    VEC_LOOP_2_COMP_LOOP_C_10 = 9'd302,
    VEC_LOOP_2_COMP_LOOP_C_11 = 9'd303,
    VEC_LOOP_2_COMP_LOOP_C_12 = 9'd304,
    VEC_LOOP_2_COMP_LOOP_C_13 = 9'd305,
    VEC_LOOP_2_COMP_LOOP_C_14 = 9'd306,
    VEC_LOOP_2_COMP_LOOP_C_15 = 9'd307,
    VEC_LOOP_2_COMP_LOOP_C_16 = 9'd308,
    VEC_LOOP_2_COMP_LOOP_C_17 = 9'd309,
    VEC_LOOP_2_COMP_LOOP_C_18 = 9'd310,
    VEC_LOOP_2_COMP_LOOP_C_19 = 9'd311,
    VEC_LOOP_2_COMP_LOOP_C_20 = 9'd312,
    VEC_LOOP_2_COMP_LOOP_C_21 = 9'd313,
    VEC_LOOP_2_COMP_LOOP_C_22 = 9'd314,
    VEC_LOOP_2_COMP_LOOP_C_23 = 9'd315,
    VEC_LOOP_2_COMP_LOOP_C_24 = 9'd316,
    VEC_LOOP_2_COMP_LOOP_C_25 = 9'd317,
    VEC_LOOP_2_COMP_LOOP_C_26 = 9'd318,
    VEC_LOOP_2_COMP_LOOP_C_27 = 9'd319,
    VEC_LOOP_2_COMP_LOOP_C_28 = 9'd320,
    VEC_LOOP_2_COMP_LOOP_C_29 = 9'd321,
    VEC_LOOP_2_COMP_LOOP_C_30 = 9'd322,
    VEC_LOOP_2_COMP_LOOP_C_31 = 9'd323,
    VEC_LOOP_2_COMP_LOOP_C_32 = 9'd324,
    VEC_LOOP_2_COMP_LOOP_C_33 = 9'd325,
    VEC_LOOP_2_COMP_LOOP_C_34 = 9'd326,
    VEC_LOOP_2_COMP_LOOP_C_35 = 9'd327,
    VEC_LOOP_2_COMP_LOOP_C_36 = 9'd328,
    VEC_LOOP_2_COMP_LOOP_C_37 = 9'd329,
    VEC_LOOP_2_COMP_LOOP_C_38 = 9'd330,
    VEC_LOOP_2_COMP_LOOP_C_39 = 9'd331,
    VEC_LOOP_2_COMP_LOOP_C_40 = 9'd332,
    VEC_LOOP_2_COMP_LOOP_C_41 = 9'd333,
    VEC_LOOP_2_COMP_LOOP_C_42 = 9'd334,
    VEC_LOOP_2_COMP_LOOP_C_43 = 9'd335,
    VEC_LOOP_2_COMP_LOOP_C_44 = 9'd336,
    VEC_LOOP_2_COMP_LOOP_C_45 = 9'd337,
    VEC_LOOP_2_COMP_LOOP_C_46 = 9'd338,
    VEC_LOOP_2_COMP_LOOP_C_47 = 9'd339,
    VEC_LOOP_2_COMP_LOOP_C_48 = 9'd340,
    VEC_LOOP_2_COMP_LOOP_C_49 = 9'd341,
    VEC_LOOP_2_COMP_LOOP_C_50 = 9'd342,
    VEC_LOOP_2_COMP_LOOP_C_51 = 9'd343,
    VEC_LOOP_2_COMP_LOOP_C_52 = 9'd344,
    VEC_LOOP_2_COMP_LOOP_C_53 = 9'd345,
    VEC_LOOP_2_COMP_LOOP_C_54 = 9'd346,
    VEC_LOOP_2_COMP_LOOP_C_55 = 9'd347,
    VEC_LOOP_2_COMP_LOOP_C_56 = 9'd348,
    VEC_LOOP_2_COMP_LOOP_C_57 = 9'd349,
    VEC_LOOP_2_COMP_LOOP_C_58 = 9'd350,
    VEC_LOOP_2_COMP_LOOP_C_59 = 9'd351,
    VEC_LOOP_2_COMP_LOOP_C_60 = 9'd352,
    VEC_LOOP_2_COMP_LOOP_C_61 = 9'd353,
    VEC_LOOP_2_COMP_LOOP_C_62 = 9'd354,
    VEC_LOOP_2_COMP_LOOP_C_63 = 9'd355,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0 = 9'd356,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1 = 9'd357,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2 = 9'd358,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3 = 9'd359,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4 = 9'd360,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5 = 9'd361,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6 = 9'd362,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7 = 9'd363,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8 = 9'd364,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9 = 9'd365,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10 = 9'd366,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11 = 9'd367,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12 = 9'd368,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13 = 9'd369,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14 = 9'd370,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15 = 9'd371,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16 = 9'd372,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17 = 9'd373,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18 = 9'd374,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19 = 9'd375,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20 = 9'd376,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21 = 9'd377,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22 = 9'd378,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23 = 9'd379,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24 = 9'd380,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_25 = 9'd381,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_26 = 9'd382,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_27 = 9'd383,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_28 = 9'd384,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_29 = 9'd385,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_30 = 9'd386,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_31 = 9'd387,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_32 = 9'd388,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_33 = 9'd389,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_34 = 9'd390,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_35 = 9'd391,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_36 = 9'd392,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_37 = 9'd393,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38 = 9'd394,
    VEC_LOOP_2_COMP_LOOP_C_64 = 9'd395,
    VEC_LOOP_2_COMP_LOOP_C_65 = 9'd396,
    VEC_LOOP_2_COMP_LOOP_C_66 = 9'd397,
    VEC_LOOP_2_COMP_LOOP_C_67 = 9'd398,
    VEC_LOOP_2_COMP_LOOP_C_68 = 9'd399,
    VEC_LOOP_2_COMP_LOOP_C_69 = 9'd400,
    VEC_LOOP_2_COMP_LOOP_C_70 = 9'd401,
    VEC_LOOP_2_COMP_LOOP_C_71 = 9'd402,
    VEC_LOOP_2_COMP_LOOP_C_72 = 9'd403,
    VEC_LOOP_2_COMP_LOOP_C_73 = 9'd404,
    VEC_LOOP_2_COMP_LOOP_C_74 = 9'd405,
    VEC_LOOP_2_COMP_LOOP_C_75 = 9'd406,
    VEC_LOOP_2_COMP_LOOP_C_76 = 9'd407,
    VEC_LOOP_2_COMP_LOOP_C_77 = 9'd408,
    VEC_LOOP_2_COMP_LOOP_C_78 = 9'd409,
    VEC_LOOP_2_COMP_LOOP_C_79 = 9'd410,
    VEC_LOOP_2_COMP_LOOP_C_80 = 9'd411,
    VEC_LOOP_2_COMP_LOOP_C_81 = 9'd412,
    VEC_LOOP_2_COMP_LOOP_C_82 = 9'd413,
    VEC_LOOP_2_COMP_LOOP_C_83 = 9'd414,
    VEC_LOOP_2_COMP_LOOP_C_84 = 9'd415,
    VEC_LOOP_2_COMP_LOOP_C_85 = 9'd416,
    VEC_LOOP_2_COMP_LOOP_C_86 = 9'd417,
    VEC_LOOP_2_COMP_LOOP_C_87 = 9'd418,
    VEC_LOOP_2_COMP_LOOP_C_88 = 9'd419,
    VEC_LOOP_2_COMP_LOOP_C_89 = 9'd420,
    VEC_LOOP_2_COMP_LOOP_C_90 = 9'd421,
    VEC_LOOP_2_COMP_LOOP_C_91 = 9'd422,
    VEC_LOOP_2_COMP_LOOP_C_92 = 9'd423,
    VEC_LOOP_2_COMP_LOOP_C_93 = 9'd424,
    VEC_LOOP_2_COMP_LOOP_C_94 = 9'd425,
    VEC_LOOP_2_COMP_LOOP_C_95 = 9'd426,
    VEC_LOOP_2_COMP_LOOP_C_96 = 9'd427,
    VEC_LOOP_2_COMP_LOOP_C_97 = 9'd428,
    VEC_LOOP_2_COMP_LOOP_C_98 = 9'd429,
    VEC_LOOP_2_COMP_LOOP_C_99 = 9'd430,
    VEC_LOOP_2_COMP_LOOP_C_100 = 9'd431,
    VEC_LOOP_2_COMP_LOOP_C_101 = 9'd432,
    VEC_LOOP_2_COMP_LOOP_C_102 = 9'd433,
    VEC_LOOP_2_COMP_LOOP_C_103 = 9'd434,
    VEC_LOOP_2_COMP_LOOP_C_104 = 9'd435,
    VEC_LOOP_2_COMP_LOOP_C_105 = 9'd436,
    VEC_LOOP_2_COMP_LOOP_C_106 = 9'd437,
    VEC_LOOP_2_COMP_LOOP_C_107 = 9'd438,
    VEC_LOOP_2_COMP_LOOP_C_108 = 9'd439,
    VEC_LOOP_2_COMP_LOOP_C_109 = 9'd440,
    VEC_LOOP_2_COMP_LOOP_C_110 = 9'd441,
    VEC_LOOP_2_COMP_LOOP_C_111 = 9'd442,
    VEC_LOOP_2_COMP_LOOP_C_112 = 9'd443,
    VEC_LOOP_2_COMP_LOOP_C_113 = 9'd444,
    VEC_LOOP_2_COMP_LOOP_C_114 = 9'd445,
    VEC_LOOP_2_COMP_LOOP_C_115 = 9'd446,
    VEC_LOOP_2_COMP_LOOP_C_116 = 9'd447,
    VEC_LOOP_2_COMP_LOOP_C_117 = 9'd448,
    VEC_LOOP_2_COMP_LOOP_C_118 = 9'd449,
    VEC_LOOP_2_COMP_LOOP_C_119 = 9'd450,
    VEC_LOOP_2_COMP_LOOP_C_120 = 9'd451,
    VEC_LOOP_2_COMP_LOOP_C_121 = 9'd452,
    VEC_LOOP_2_COMP_LOOP_C_122 = 9'd453,
    VEC_LOOP_2_COMP_LOOP_C_123 = 9'd454,
    VEC_LOOP_2_COMP_LOOP_C_124 = 9'd455,
    VEC_LOOP_C_1 = 9'd456,
    STAGE_LOOP_C_9 = 9'd457,
    main_C_1 = 9'd458;

  reg [8:0] state_var;
  reg [8:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 9'b000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 9'b000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 9'b000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 9'b000000100;
        state_var_NS = STAGE_LOOP_C_4;
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 9'b000000101;
        state_var_NS = STAGE_LOOP_C_5;
      end
      STAGE_LOOP_C_5 : begin
        fsm_output = 9'b000000110;
        state_var_NS = STAGE_LOOP_C_6;
      end
      STAGE_LOOP_C_6 : begin
        fsm_output = 9'b000000111;
        state_var_NS = STAGE_LOOP_C_7;
      end
      STAGE_LOOP_C_7 : begin
        fsm_output = 9'b000001000;
        state_var_NS = STAGE_LOOP_C_8;
      end
      STAGE_LOOP_C_8 : begin
        fsm_output = 9'b000001001;
        if ( STAGE_LOOP_C_8_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      modExp_while_C_0 : begin
        fsm_output = 9'b000001010;
        state_var_NS = modExp_while_C_1;
      end
      modExp_while_C_1 : begin
        fsm_output = 9'b000001011;
        state_var_NS = modExp_while_C_2;
      end
      modExp_while_C_2 : begin
        fsm_output = 9'b000001100;
        state_var_NS = modExp_while_C_3;
      end
      modExp_while_C_3 : begin
        fsm_output = 9'b000001101;
        state_var_NS = modExp_while_C_4;
      end
      modExp_while_C_4 : begin
        fsm_output = 9'b000001110;
        state_var_NS = modExp_while_C_5;
      end
      modExp_while_C_5 : begin
        fsm_output = 9'b000001111;
        state_var_NS = modExp_while_C_6;
      end
      modExp_while_C_6 : begin
        fsm_output = 9'b000010000;
        state_var_NS = modExp_while_C_7;
      end
      modExp_while_C_7 : begin
        fsm_output = 9'b000010001;
        state_var_NS = modExp_while_C_8;
      end
      modExp_while_C_8 : begin
        fsm_output = 9'b000010010;
        state_var_NS = modExp_while_C_9;
      end
      modExp_while_C_9 : begin
        fsm_output = 9'b000010011;
        state_var_NS = modExp_while_C_10;
      end
      modExp_while_C_10 : begin
        fsm_output = 9'b000010100;
        state_var_NS = modExp_while_C_11;
      end
      modExp_while_C_11 : begin
        fsm_output = 9'b000010101;
        state_var_NS = modExp_while_C_12;
      end
      modExp_while_C_12 : begin
        fsm_output = 9'b000010110;
        state_var_NS = modExp_while_C_13;
      end
      modExp_while_C_13 : begin
        fsm_output = 9'b000010111;
        state_var_NS = modExp_while_C_14;
      end
      modExp_while_C_14 : begin
        fsm_output = 9'b000011000;
        state_var_NS = modExp_while_C_15;
      end
      modExp_while_C_15 : begin
        fsm_output = 9'b000011001;
        state_var_NS = modExp_while_C_16;
      end
      modExp_while_C_16 : begin
        fsm_output = 9'b000011010;
        state_var_NS = modExp_while_C_17;
      end
      modExp_while_C_17 : begin
        fsm_output = 9'b000011011;
        state_var_NS = modExp_while_C_18;
      end
      modExp_while_C_18 : begin
        fsm_output = 9'b000011100;
        state_var_NS = modExp_while_C_19;
      end
      modExp_while_C_19 : begin
        fsm_output = 9'b000011101;
        state_var_NS = modExp_while_C_20;
      end
      modExp_while_C_20 : begin
        fsm_output = 9'b000011110;
        state_var_NS = modExp_while_C_21;
      end
      modExp_while_C_21 : begin
        fsm_output = 9'b000011111;
        state_var_NS = modExp_while_C_22;
      end
      modExp_while_C_22 : begin
        fsm_output = 9'b000100000;
        state_var_NS = modExp_while_C_23;
      end
      modExp_while_C_23 : begin
        fsm_output = 9'b000100001;
        state_var_NS = modExp_while_C_24;
      end
      modExp_while_C_24 : begin
        fsm_output = 9'b000100010;
        state_var_NS = modExp_while_C_25;
      end
      modExp_while_C_25 : begin
        fsm_output = 9'b000100011;
        state_var_NS = modExp_while_C_26;
      end
      modExp_while_C_26 : begin
        fsm_output = 9'b000100100;
        state_var_NS = modExp_while_C_27;
      end
      modExp_while_C_27 : begin
        fsm_output = 9'b000100101;
        state_var_NS = modExp_while_C_28;
      end
      modExp_while_C_28 : begin
        fsm_output = 9'b000100110;
        state_var_NS = modExp_while_C_29;
      end
      modExp_while_C_29 : begin
        fsm_output = 9'b000100111;
        state_var_NS = modExp_while_C_30;
      end
      modExp_while_C_30 : begin
        fsm_output = 9'b000101000;
        state_var_NS = modExp_while_C_31;
      end
      modExp_while_C_31 : begin
        fsm_output = 9'b000101001;
        state_var_NS = modExp_while_C_32;
      end
      modExp_while_C_32 : begin
        fsm_output = 9'b000101010;
        state_var_NS = modExp_while_C_33;
      end
      modExp_while_C_33 : begin
        fsm_output = 9'b000101011;
        state_var_NS = modExp_while_C_34;
      end
      modExp_while_C_34 : begin
        fsm_output = 9'b000101100;
        state_var_NS = modExp_while_C_35;
      end
      modExp_while_C_35 : begin
        fsm_output = 9'b000101101;
        state_var_NS = modExp_while_C_36;
      end
      modExp_while_C_36 : begin
        fsm_output = 9'b000101110;
        state_var_NS = modExp_while_C_37;
      end
      modExp_while_C_37 : begin
        fsm_output = 9'b000101111;
        state_var_NS = modExp_while_C_38;
      end
      modExp_while_C_38 : begin
        fsm_output = 9'b000110000;
        if ( modExp_while_C_38_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_0 : begin
        fsm_output = 9'b000110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_C_1 : begin
        fsm_output = 9'b000110010;
        if ( VEC_LOOP_1_COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 9'b000110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 9'b000110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 9'b000110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 9'b000110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 9'b000110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 9'b000111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 9'b000111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 9'b000111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 9'b000111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 9'b000111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 9'b000111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 9'b000111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 9'b000111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 9'b001000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 9'b001000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 9'b001000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 9'b001000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 9'b001000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 9'b001000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 9'b001000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 9'b001000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 9'b001001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 9'b001001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 9'b001001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 9'b001001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_25;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 9'b001001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_26;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 9'b001001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_27;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 9'b001001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_28;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 9'b001001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_29;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 9'b001010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_30;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 9'b001010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_31;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 9'b001010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_32;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 9'b001010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_33;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 9'b001010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_34;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 9'b001010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_35;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 9'b001010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_36;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 9'b001010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_37;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 9'b001011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 9'b001011001;
        if ( VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_2 : begin
        fsm_output = 9'b001011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_C_3 : begin
        fsm_output = 9'b001011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_C_4 : begin
        fsm_output = 9'b001011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_C_5 : begin
        fsm_output = 9'b001011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_C_6 : begin
        fsm_output = 9'b001011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_C_7 : begin
        fsm_output = 9'b001011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_C_8 : begin
        fsm_output = 9'b001100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_C_9 : begin
        fsm_output = 9'b001100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_C_10 : begin
        fsm_output = 9'b001100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_C_11 : begin
        fsm_output = 9'b001100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_C_12 : begin
        fsm_output = 9'b001100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_C_13 : begin
        fsm_output = 9'b001100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_C_14 : begin
        fsm_output = 9'b001100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_C_15 : begin
        fsm_output = 9'b001100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_C_16 : begin
        fsm_output = 9'b001101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_C_17 : begin
        fsm_output = 9'b001101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_C_18 : begin
        fsm_output = 9'b001101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_C_19 : begin
        fsm_output = 9'b001101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_C_20 : begin
        fsm_output = 9'b001101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_C_21 : begin
        fsm_output = 9'b001101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_C_22 : begin
        fsm_output = 9'b001101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_C_23 : begin
        fsm_output = 9'b001101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_C_24 : begin
        fsm_output = 9'b001110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_25;
      end
      VEC_LOOP_1_COMP_LOOP_C_25 : begin
        fsm_output = 9'b001110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_26;
      end
      VEC_LOOP_1_COMP_LOOP_C_26 : begin
        fsm_output = 9'b001110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_27;
      end
      VEC_LOOP_1_COMP_LOOP_C_27 : begin
        fsm_output = 9'b001110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_28;
      end
      VEC_LOOP_1_COMP_LOOP_C_28 : begin
        fsm_output = 9'b001110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_29;
      end
      VEC_LOOP_1_COMP_LOOP_C_29 : begin
        fsm_output = 9'b001110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_30;
      end
      VEC_LOOP_1_COMP_LOOP_C_30 : begin
        fsm_output = 9'b001110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_31;
      end
      VEC_LOOP_1_COMP_LOOP_C_31 : begin
        fsm_output = 9'b001110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_32;
      end
      VEC_LOOP_1_COMP_LOOP_C_32 : begin
        fsm_output = 9'b001111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_33;
      end
      VEC_LOOP_1_COMP_LOOP_C_33 : begin
        fsm_output = 9'b001111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_34;
      end
      VEC_LOOP_1_COMP_LOOP_C_34 : begin
        fsm_output = 9'b001111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_35;
      end
      VEC_LOOP_1_COMP_LOOP_C_35 : begin
        fsm_output = 9'b001111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_36;
      end
      VEC_LOOP_1_COMP_LOOP_C_36 : begin
        fsm_output = 9'b001111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_37;
      end
      VEC_LOOP_1_COMP_LOOP_C_37 : begin
        fsm_output = 9'b001111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_38;
      end
      VEC_LOOP_1_COMP_LOOP_C_38 : begin
        fsm_output = 9'b001111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_39;
      end
      VEC_LOOP_1_COMP_LOOP_C_39 : begin
        fsm_output = 9'b001111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_40;
      end
      VEC_LOOP_1_COMP_LOOP_C_40 : begin
        fsm_output = 9'b010000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_41;
      end
      VEC_LOOP_1_COMP_LOOP_C_41 : begin
        fsm_output = 9'b010000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_42;
      end
      VEC_LOOP_1_COMP_LOOP_C_42 : begin
        fsm_output = 9'b010000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_43;
      end
      VEC_LOOP_1_COMP_LOOP_C_43 : begin
        fsm_output = 9'b010000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_44;
      end
      VEC_LOOP_1_COMP_LOOP_C_44 : begin
        fsm_output = 9'b010000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_45;
      end
      VEC_LOOP_1_COMP_LOOP_C_45 : begin
        fsm_output = 9'b010000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_46;
      end
      VEC_LOOP_1_COMP_LOOP_C_46 : begin
        fsm_output = 9'b010000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_47;
      end
      VEC_LOOP_1_COMP_LOOP_C_47 : begin
        fsm_output = 9'b010000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_48;
      end
      VEC_LOOP_1_COMP_LOOP_C_48 : begin
        fsm_output = 9'b010001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_49;
      end
      VEC_LOOP_1_COMP_LOOP_C_49 : begin
        fsm_output = 9'b010001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_50;
      end
      VEC_LOOP_1_COMP_LOOP_C_50 : begin
        fsm_output = 9'b010001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_51;
      end
      VEC_LOOP_1_COMP_LOOP_C_51 : begin
        fsm_output = 9'b010001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_52;
      end
      VEC_LOOP_1_COMP_LOOP_C_52 : begin
        fsm_output = 9'b010001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_53;
      end
      VEC_LOOP_1_COMP_LOOP_C_53 : begin
        fsm_output = 9'b010001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_54;
      end
      VEC_LOOP_1_COMP_LOOP_C_54 : begin
        fsm_output = 9'b010001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_55;
      end
      VEC_LOOP_1_COMP_LOOP_C_55 : begin
        fsm_output = 9'b010001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_56;
      end
      VEC_LOOP_1_COMP_LOOP_C_56 : begin
        fsm_output = 9'b010010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_57;
      end
      VEC_LOOP_1_COMP_LOOP_C_57 : begin
        fsm_output = 9'b010010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_58;
      end
      VEC_LOOP_1_COMP_LOOP_C_58 : begin
        fsm_output = 9'b010010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_59;
      end
      VEC_LOOP_1_COMP_LOOP_C_59 : begin
        fsm_output = 9'b010010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_60;
      end
      VEC_LOOP_1_COMP_LOOP_C_60 : begin
        fsm_output = 9'b010010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_61;
      end
      VEC_LOOP_1_COMP_LOOP_C_61 : begin
        fsm_output = 9'b010010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_62;
      end
      VEC_LOOP_1_COMP_LOOP_C_62 : begin
        fsm_output = 9'b010010110;
        if ( VEC_LOOP_1_COMP_LOOP_C_62_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_63;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_63 : begin
        fsm_output = 9'b010010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 9'b010011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 9'b010011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 9'b010011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 9'b010011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 9'b010011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 9'b010011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 9'b010011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 9'b010011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 9'b010100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 9'b010100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 9'b010100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 9'b010100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 9'b010100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 9'b010100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 9'b010100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 9'b010100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 9'b010101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 9'b010101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 9'b010101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 9'b010101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 9'b010101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 9'b010101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 9'b010101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 9'b010101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 9'b010110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_25;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 9'b010110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_26;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 9'b010110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_27;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 9'b010110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_28;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 9'b010110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_29;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 9'b010110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_30;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 9'b010110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_31;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 9'b010110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_32;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 9'b010111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_33;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 9'b010111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_34;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 9'b010111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_35;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 9'b010111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_36;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 9'b010111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_37;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 9'b010111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 9'b010111110;
        if ( VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_64;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_64 : begin
        fsm_output = 9'b010111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_65;
      end
      VEC_LOOP_1_COMP_LOOP_C_65 : begin
        fsm_output = 9'b011000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_66;
      end
      VEC_LOOP_1_COMP_LOOP_C_66 : begin
        fsm_output = 9'b011000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_67;
      end
      VEC_LOOP_1_COMP_LOOP_C_67 : begin
        fsm_output = 9'b011000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_68;
      end
      VEC_LOOP_1_COMP_LOOP_C_68 : begin
        fsm_output = 9'b011000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_69;
      end
      VEC_LOOP_1_COMP_LOOP_C_69 : begin
        fsm_output = 9'b011000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_70;
      end
      VEC_LOOP_1_COMP_LOOP_C_70 : begin
        fsm_output = 9'b011000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_71;
      end
      VEC_LOOP_1_COMP_LOOP_C_71 : begin
        fsm_output = 9'b011000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_72;
      end
      VEC_LOOP_1_COMP_LOOP_C_72 : begin
        fsm_output = 9'b011000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_73;
      end
      VEC_LOOP_1_COMP_LOOP_C_73 : begin
        fsm_output = 9'b011001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_74;
      end
      VEC_LOOP_1_COMP_LOOP_C_74 : begin
        fsm_output = 9'b011001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_75;
      end
      VEC_LOOP_1_COMP_LOOP_C_75 : begin
        fsm_output = 9'b011001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_76;
      end
      VEC_LOOP_1_COMP_LOOP_C_76 : begin
        fsm_output = 9'b011001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_77;
      end
      VEC_LOOP_1_COMP_LOOP_C_77 : begin
        fsm_output = 9'b011001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_78;
      end
      VEC_LOOP_1_COMP_LOOP_C_78 : begin
        fsm_output = 9'b011001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_79;
      end
      VEC_LOOP_1_COMP_LOOP_C_79 : begin
        fsm_output = 9'b011001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_80;
      end
      VEC_LOOP_1_COMP_LOOP_C_80 : begin
        fsm_output = 9'b011001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_81;
      end
      VEC_LOOP_1_COMP_LOOP_C_81 : begin
        fsm_output = 9'b011010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_82;
      end
      VEC_LOOP_1_COMP_LOOP_C_82 : begin
        fsm_output = 9'b011010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_83;
      end
      VEC_LOOP_1_COMP_LOOP_C_83 : begin
        fsm_output = 9'b011010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_84;
      end
      VEC_LOOP_1_COMP_LOOP_C_84 : begin
        fsm_output = 9'b011010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_85;
      end
      VEC_LOOP_1_COMP_LOOP_C_85 : begin
        fsm_output = 9'b011010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_86;
      end
      VEC_LOOP_1_COMP_LOOP_C_86 : begin
        fsm_output = 9'b011010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_87;
      end
      VEC_LOOP_1_COMP_LOOP_C_87 : begin
        fsm_output = 9'b011010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_88;
      end
      VEC_LOOP_1_COMP_LOOP_C_88 : begin
        fsm_output = 9'b011010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_89;
      end
      VEC_LOOP_1_COMP_LOOP_C_89 : begin
        fsm_output = 9'b011011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_90;
      end
      VEC_LOOP_1_COMP_LOOP_C_90 : begin
        fsm_output = 9'b011011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_91;
      end
      VEC_LOOP_1_COMP_LOOP_C_91 : begin
        fsm_output = 9'b011011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_92;
      end
      VEC_LOOP_1_COMP_LOOP_C_92 : begin
        fsm_output = 9'b011011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_93;
      end
      VEC_LOOP_1_COMP_LOOP_C_93 : begin
        fsm_output = 9'b011011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_94;
      end
      VEC_LOOP_1_COMP_LOOP_C_94 : begin
        fsm_output = 9'b011011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_95;
      end
      VEC_LOOP_1_COMP_LOOP_C_95 : begin
        fsm_output = 9'b011011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_96;
      end
      VEC_LOOP_1_COMP_LOOP_C_96 : begin
        fsm_output = 9'b011011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_97;
      end
      VEC_LOOP_1_COMP_LOOP_C_97 : begin
        fsm_output = 9'b011100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_98;
      end
      VEC_LOOP_1_COMP_LOOP_C_98 : begin
        fsm_output = 9'b011100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_99;
      end
      VEC_LOOP_1_COMP_LOOP_C_99 : begin
        fsm_output = 9'b011100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_100;
      end
      VEC_LOOP_1_COMP_LOOP_C_100 : begin
        fsm_output = 9'b011100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_101;
      end
      VEC_LOOP_1_COMP_LOOP_C_101 : begin
        fsm_output = 9'b011100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_102;
      end
      VEC_LOOP_1_COMP_LOOP_C_102 : begin
        fsm_output = 9'b011100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_103;
      end
      VEC_LOOP_1_COMP_LOOP_C_103 : begin
        fsm_output = 9'b011100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_104;
      end
      VEC_LOOP_1_COMP_LOOP_C_104 : begin
        fsm_output = 9'b011100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_105;
      end
      VEC_LOOP_1_COMP_LOOP_C_105 : begin
        fsm_output = 9'b011101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_106;
      end
      VEC_LOOP_1_COMP_LOOP_C_106 : begin
        fsm_output = 9'b011101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_107;
      end
      VEC_LOOP_1_COMP_LOOP_C_107 : begin
        fsm_output = 9'b011101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_108;
      end
      VEC_LOOP_1_COMP_LOOP_C_108 : begin
        fsm_output = 9'b011101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_109;
      end
      VEC_LOOP_1_COMP_LOOP_C_109 : begin
        fsm_output = 9'b011101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_110;
      end
      VEC_LOOP_1_COMP_LOOP_C_110 : begin
        fsm_output = 9'b011101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_111;
      end
      VEC_LOOP_1_COMP_LOOP_C_111 : begin
        fsm_output = 9'b011101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_112;
      end
      VEC_LOOP_1_COMP_LOOP_C_112 : begin
        fsm_output = 9'b011101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_113;
      end
      VEC_LOOP_1_COMP_LOOP_C_113 : begin
        fsm_output = 9'b011110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_114;
      end
      VEC_LOOP_1_COMP_LOOP_C_114 : begin
        fsm_output = 9'b011110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_115;
      end
      VEC_LOOP_1_COMP_LOOP_C_115 : begin
        fsm_output = 9'b011110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_116;
      end
      VEC_LOOP_1_COMP_LOOP_C_116 : begin
        fsm_output = 9'b011110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_117;
      end
      VEC_LOOP_1_COMP_LOOP_C_117 : begin
        fsm_output = 9'b011110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_118;
      end
      VEC_LOOP_1_COMP_LOOP_C_118 : begin
        fsm_output = 9'b011110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_119;
      end
      VEC_LOOP_1_COMP_LOOP_C_119 : begin
        fsm_output = 9'b011110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_120;
      end
      VEC_LOOP_1_COMP_LOOP_C_120 : begin
        fsm_output = 9'b011110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_121;
      end
      VEC_LOOP_1_COMP_LOOP_C_121 : begin
        fsm_output = 9'b011111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_122;
      end
      VEC_LOOP_1_COMP_LOOP_C_122 : begin
        fsm_output = 9'b011111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_123;
      end
      VEC_LOOP_1_COMP_LOOP_C_123 : begin
        fsm_output = 9'b011111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_124;
      end
      VEC_LOOP_1_COMP_LOOP_C_124 : begin
        fsm_output = 9'b011111011;
        if ( VEC_LOOP_1_COMP_LOOP_C_124_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 9'b011111100;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_9;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_0 : begin
        fsm_output = 9'b011111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_C_1 : begin
        fsm_output = 9'b011111110;
        if ( VEC_LOOP_2_COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 9'b011111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 9'b100000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 9'b100000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 9'b100000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 9'b100000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 9'b100000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 9'b100000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 9'b100000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 9'b100000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 9'b100001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 9'b100001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 9'b100001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 9'b100001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 9'b100001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 9'b100001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 9'b100001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 9'b100001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 9'b100010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 9'b100010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 9'b100010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 9'b100010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 9'b100010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 9'b100010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 9'b100010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 9'b100010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_25;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 9'b100011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_26;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 9'b100011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_27;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 9'b100011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_28;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 9'b100011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_29;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 9'b100011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_30;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 9'b100011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_31;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 9'b100011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_32;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 9'b100011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_33;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 9'b100100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_34;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 9'b100100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_35;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 9'b100100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_36;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 9'b100100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_37;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 9'b100100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 9'b100100101;
        if ( VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_2 : begin
        fsm_output = 9'b100100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_C_3 : begin
        fsm_output = 9'b100100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_C_4 : begin
        fsm_output = 9'b100101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_C_5 : begin
        fsm_output = 9'b100101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_C_6 : begin
        fsm_output = 9'b100101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_C_7 : begin
        fsm_output = 9'b100101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_C_8 : begin
        fsm_output = 9'b100101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_C_9 : begin
        fsm_output = 9'b100101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_C_10 : begin
        fsm_output = 9'b100101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_C_11 : begin
        fsm_output = 9'b100101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_C_12 : begin
        fsm_output = 9'b100110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_C_13 : begin
        fsm_output = 9'b100110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_C_14 : begin
        fsm_output = 9'b100110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_C_15 : begin
        fsm_output = 9'b100110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_C_16 : begin
        fsm_output = 9'b100110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_C_17 : begin
        fsm_output = 9'b100110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_C_18 : begin
        fsm_output = 9'b100110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_C_19 : begin
        fsm_output = 9'b100110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_C_20 : begin
        fsm_output = 9'b100111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_C_21 : begin
        fsm_output = 9'b100111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_C_22 : begin
        fsm_output = 9'b100111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_C_23 : begin
        fsm_output = 9'b100111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_C_24 : begin
        fsm_output = 9'b100111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_25;
      end
      VEC_LOOP_2_COMP_LOOP_C_25 : begin
        fsm_output = 9'b100111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_26;
      end
      VEC_LOOP_2_COMP_LOOP_C_26 : begin
        fsm_output = 9'b100111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_27;
      end
      VEC_LOOP_2_COMP_LOOP_C_27 : begin
        fsm_output = 9'b100111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_28;
      end
      VEC_LOOP_2_COMP_LOOP_C_28 : begin
        fsm_output = 9'b101000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_29;
      end
      VEC_LOOP_2_COMP_LOOP_C_29 : begin
        fsm_output = 9'b101000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_30;
      end
      VEC_LOOP_2_COMP_LOOP_C_30 : begin
        fsm_output = 9'b101000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_31;
      end
      VEC_LOOP_2_COMP_LOOP_C_31 : begin
        fsm_output = 9'b101000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_32;
      end
      VEC_LOOP_2_COMP_LOOP_C_32 : begin
        fsm_output = 9'b101000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_33;
      end
      VEC_LOOP_2_COMP_LOOP_C_33 : begin
        fsm_output = 9'b101000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_34;
      end
      VEC_LOOP_2_COMP_LOOP_C_34 : begin
        fsm_output = 9'b101000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_35;
      end
      VEC_LOOP_2_COMP_LOOP_C_35 : begin
        fsm_output = 9'b101000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_36;
      end
      VEC_LOOP_2_COMP_LOOP_C_36 : begin
        fsm_output = 9'b101001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_37;
      end
      VEC_LOOP_2_COMP_LOOP_C_37 : begin
        fsm_output = 9'b101001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_38;
      end
      VEC_LOOP_2_COMP_LOOP_C_38 : begin
        fsm_output = 9'b101001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_39;
      end
      VEC_LOOP_2_COMP_LOOP_C_39 : begin
        fsm_output = 9'b101001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_40;
      end
      VEC_LOOP_2_COMP_LOOP_C_40 : begin
        fsm_output = 9'b101001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_41;
      end
      VEC_LOOP_2_COMP_LOOP_C_41 : begin
        fsm_output = 9'b101001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_42;
      end
      VEC_LOOP_2_COMP_LOOP_C_42 : begin
        fsm_output = 9'b101001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_43;
      end
      VEC_LOOP_2_COMP_LOOP_C_43 : begin
        fsm_output = 9'b101001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_44;
      end
      VEC_LOOP_2_COMP_LOOP_C_44 : begin
        fsm_output = 9'b101010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_45;
      end
      VEC_LOOP_2_COMP_LOOP_C_45 : begin
        fsm_output = 9'b101010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_46;
      end
      VEC_LOOP_2_COMP_LOOP_C_46 : begin
        fsm_output = 9'b101010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_47;
      end
      VEC_LOOP_2_COMP_LOOP_C_47 : begin
        fsm_output = 9'b101010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_48;
      end
      VEC_LOOP_2_COMP_LOOP_C_48 : begin
        fsm_output = 9'b101010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_49;
      end
      VEC_LOOP_2_COMP_LOOP_C_49 : begin
        fsm_output = 9'b101010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_50;
      end
      VEC_LOOP_2_COMP_LOOP_C_50 : begin
        fsm_output = 9'b101010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_51;
      end
      VEC_LOOP_2_COMP_LOOP_C_51 : begin
        fsm_output = 9'b101010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_52;
      end
      VEC_LOOP_2_COMP_LOOP_C_52 : begin
        fsm_output = 9'b101011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_53;
      end
      VEC_LOOP_2_COMP_LOOP_C_53 : begin
        fsm_output = 9'b101011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_54;
      end
      VEC_LOOP_2_COMP_LOOP_C_54 : begin
        fsm_output = 9'b101011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_55;
      end
      VEC_LOOP_2_COMP_LOOP_C_55 : begin
        fsm_output = 9'b101011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_56;
      end
      VEC_LOOP_2_COMP_LOOP_C_56 : begin
        fsm_output = 9'b101011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_57;
      end
      VEC_LOOP_2_COMP_LOOP_C_57 : begin
        fsm_output = 9'b101011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_58;
      end
      VEC_LOOP_2_COMP_LOOP_C_58 : begin
        fsm_output = 9'b101011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_59;
      end
      VEC_LOOP_2_COMP_LOOP_C_59 : begin
        fsm_output = 9'b101011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_60;
      end
      VEC_LOOP_2_COMP_LOOP_C_60 : begin
        fsm_output = 9'b101100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_61;
      end
      VEC_LOOP_2_COMP_LOOP_C_61 : begin
        fsm_output = 9'b101100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_62;
      end
      VEC_LOOP_2_COMP_LOOP_C_62 : begin
        fsm_output = 9'b101100010;
        if ( VEC_LOOP_2_COMP_LOOP_C_62_tr0 ) begin
          state_var_NS = VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_63;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_63 : begin
        fsm_output = 9'b101100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 9'b101100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 9'b101100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 9'b101100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 9'b101100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 9'b101101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 9'b101101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 9'b101101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 9'b101101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 9'b101101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 9'b101101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 9'b101101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 9'b101101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 9'b101110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 9'b101110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 9'b101110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 9'b101110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 9'b101110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 9'b101110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 9'b101110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 9'b101110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 9'b101111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 9'b101111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 9'b101111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 9'b101111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 9'b101111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_25;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 9'b101111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_26;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 9'b101111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_27;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 9'b101111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_28;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 9'b110000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_29;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 9'b110000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_30;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 9'b110000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_31;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 9'b110000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_32;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 9'b110000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_33;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 9'b110000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_34;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 9'b110000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_35;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 9'b110000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_36;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 9'b110001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_37;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 9'b110001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 9'b110001010;
        if ( VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_64;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_64 : begin
        fsm_output = 9'b110001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_65;
      end
      VEC_LOOP_2_COMP_LOOP_C_65 : begin
        fsm_output = 9'b110001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_66;
      end
      VEC_LOOP_2_COMP_LOOP_C_66 : begin
        fsm_output = 9'b110001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_67;
      end
      VEC_LOOP_2_COMP_LOOP_C_67 : begin
        fsm_output = 9'b110001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_68;
      end
      VEC_LOOP_2_COMP_LOOP_C_68 : begin
        fsm_output = 9'b110001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_69;
      end
      VEC_LOOP_2_COMP_LOOP_C_69 : begin
        fsm_output = 9'b110010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_70;
      end
      VEC_LOOP_2_COMP_LOOP_C_70 : begin
        fsm_output = 9'b110010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_71;
      end
      VEC_LOOP_2_COMP_LOOP_C_71 : begin
        fsm_output = 9'b110010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_72;
      end
      VEC_LOOP_2_COMP_LOOP_C_72 : begin
        fsm_output = 9'b110010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_73;
      end
      VEC_LOOP_2_COMP_LOOP_C_73 : begin
        fsm_output = 9'b110010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_74;
      end
      VEC_LOOP_2_COMP_LOOP_C_74 : begin
        fsm_output = 9'b110010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_75;
      end
      VEC_LOOP_2_COMP_LOOP_C_75 : begin
        fsm_output = 9'b110010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_76;
      end
      VEC_LOOP_2_COMP_LOOP_C_76 : begin
        fsm_output = 9'b110010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_77;
      end
      VEC_LOOP_2_COMP_LOOP_C_77 : begin
        fsm_output = 9'b110011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_78;
      end
      VEC_LOOP_2_COMP_LOOP_C_78 : begin
        fsm_output = 9'b110011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_79;
      end
      VEC_LOOP_2_COMP_LOOP_C_79 : begin
        fsm_output = 9'b110011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_80;
      end
      VEC_LOOP_2_COMP_LOOP_C_80 : begin
        fsm_output = 9'b110011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_81;
      end
      VEC_LOOP_2_COMP_LOOP_C_81 : begin
        fsm_output = 9'b110011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_82;
      end
      VEC_LOOP_2_COMP_LOOP_C_82 : begin
        fsm_output = 9'b110011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_83;
      end
      VEC_LOOP_2_COMP_LOOP_C_83 : begin
        fsm_output = 9'b110011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_84;
      end
      VEC_LOOP_2_COMP_LOOP_C_84 : begin
        fsm_output = 9'b110011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_85;
      end
      VEC_LOOP_2_COMP_LOOP_C_85 : begin
        fsm_output = 9'b110100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_86;
      end
      VEC_LOOP_2_COMP_LOOP_C_86 : begin
        fsm_output = 9'b110100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_87;
      end
      VEC_LOOP_2_COMP_LOOP_C_87 : begin
        fsm_output = 9'b110100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_88;
      end
      VEC_LOOP_2_COMP_LOOP_C_88 : begin
        fsm_output = 9'b110100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_89;
      end
      VEC_LOOP_2_COMP_LOOP_C_89 : begin
        fsm_output = 9'b110100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_90;
      end
      VEC_LOOP_2_COMP_LOOP_C_90 : begin
        fsm_output = 9'b110100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_91;
      end
      VEC_LOOP_2_COMP_LOOP_C_91 : begin
        fsm_output = 9'b110100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_92;
      end
      VEC_LOOP_2_COMP_LOOP_C_92 : begin
        fsm_output = 9'b110100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_93;
      end
      VEC_LOOP_2_COMP_LOOP_C_93 : begin
        fsm_output = 9'b110101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_94;
      end
      VEC_LOOP_2_COMP_LOOP_C_94 : begin
        fsm_output = 9'b110101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_95;
      end
      VEC_LOOP_2_COMP_LOOP_C_95 : begin
        fsm_output = 9'b110101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_96;
      end
      VEC_LOOP_2_COMP_LOOP_C_96 : begin
        fsm_output = 9'b110101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_97;
      end
      VEC_LOOP_2_COMP_LOOP_C_97 : begin
        fsm_output = 9'b110101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_98;
      end
      VEC_LOOP_2_COMP_LOOP_C_98 : begin
        fsm_output = 9'b110101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_99;
      end
      VEC_LOOP_2_COMP_LOOP_C_99 : begin
        fsm_output = 9'b110101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_100;
      end
      VEC_LOOP_2_COMP_LOOP_C_100 : begin
        fsm_output = 9'b110101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_101;
      end
      VEC_LOOP_2_COMP_LOOP_C_101 : begin
        fsm_output = 9'b110110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_102;
      end
      VEC_LOOP_2_COMP_LOOP_C_102 : begin
        fsm_output = 9'b110110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_103;
      end
      VEC_LOOP_2_COMP_LOOP_C_103 : begin
        fsm_output = 9'b110110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_104;
      end
      VEC_LOOP_2_COMP_LOOP_C_104 : begin
        fsm_output = 9'b110110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_105;
      end
      VEC_LOOP_2_COMP_LOOP_C_105 : begin
        fsm_output = 9'b110110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_106;
      end
      VEC_LOOP_2_COMP_LOOP_C_106 : begin
        fsm_output = 9'b110110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_107;
      end
      VEC_LOOP_2_COMP_LOOP_C_107 : begin
        fsm_output = 9'b110110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_108;
      end
      VEC_LOOP_2_COMP_LOOP_C_108 : begin
        fsm_output = 9'b110110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_109;
      end
      VEC_LOOP_2_COMP_LOOP_C_109 : begin
        fsm_output = 9'b110111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_110;
      end
      VEC_LOOP_2_COMP_LOOP_C_110 : begin
        fsm_output = 9'b110111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_111;
      end
      VEC_LOOP_2_COMP_LOOP_C_111 : begin
        fsm_output = 9'b110111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_112;
      end
      VEC_LOOP_2_COMP_LOOP_C_112 : begin
        fsm_output = 9'b110111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_113;
      end
      VEC_LOOP_2_COMP_LOOP_C_113 : begin
        fsm_output = 9'b110111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_114;
      end
      VEC_LOOP_2_COMP_LOOP_C_114 : begin
        fsm_output = 9'b110111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_115;
      end
      VEC_LOOP_2_COMP_LOOP_C_115 : begin
        fsm_output = 9'b110111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_116;
      end
      VEC_LOOP_2_COMP_LOOP_C_116 : begin
        fsm_output = 9'b110111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_117;
      end
      VEC_LOOP_2_COMP_LOOP_C_117 : begin
        fsm_output = 9'b111000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_118;
      end
      VEC_LOOP_2_COMP_LOOP_C_118 : begin
        fsm_output = 9'b111000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_119;
      end
      VEC_LOOP_2_COMP_LOOP_C_119 : begin
        fsm_output = 9'b111000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_120;
      end
      VEC_LOOP_2_COMP_LOOP_C_120 : begin
        fsm_output = 9'b111000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_121;
      end
      VEC_LOOP_2_COMP_LOOP_C_121 : begin
        fsm_output = 9'b111000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_122;
      end
      VEC_LOOP_2_COMP_LOOP_C_122 : begin
        fsm_output = 9'b111000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_123;
      end
      VEC_LOOP_2_COMP_LOOP_C_123 : begin
        fsm_output = 9'b111000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_124;
      end
      VEC_LOOP_2_COMP_LOOP_C_124 : begin
        fsm_output = 9'b111000111;
        if ( VEC_LOOP_2_COMP_LOOP_C_124_tr0 ) begin
          state_var_NS = VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_1 : begin
        fsm_output = 9'b111001000;
        if ( VEC_LOOP_C_1_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_9;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_9 : begin
        fsm_output = 9'b111001001;
        if ( STAGE_LOOP_C_9_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 9'b111001010;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 9'b000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff, vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff, vec_rsc_0_2_i_wea_d_pff,
      vec_rsc_0_3_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_qa_d;
  output vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_qa_d;
  output vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;
  output vec_rsc_0_2_i_wea_d_pff;
  output vec_rsc_0_3_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  reg [63:0] modulo_result_rem_cmp_a;
  reg [63:0] modulo_result_rem_cmp_b;
  wire [63:0] modulo_result_rem_cmp_z;
  reg [64:0] operator_66_true_div_cmp_a;
  wire [64:0] operator_66_true_div_cmp_z;
  reg [9:0] operator_66_true_div_cmp_b_9_0;
  wire [8:0] fsm_output;
  wire not_tmp_20;
  wire not_tmp_38;
  wire mux_tmp_40;
  wire or_tmp_69;
  wire or_tmp_93;
  wire and_tmp_7;
  wire mux_tmp_94;
  wire mux_tmp_95;
  wire and_dcpl_10;
  wire and_dcpl_11;
  wire and_dcpl_12;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_19;
  wire and_dcpl_21;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_29;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_37;
  wire and_dcpl_40;
  wire mux_tmp_103;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire and_dcpl_49;
  wire not_tmp_92;
  wire not_tmp_109;
  wire nor_tmp_48;
  wire and_dcpl_62;
  wire or_tmp_242;
  wire nor_tmp_51;
  wire or_tmp_244;
  wire mux_tmp_168;
  wire or_tmp_245;
  wire or_tmp_247;
  wire mux_tmp_174;
  wire mux_tmp_175;
  wire or_tmp_249;
  wire mux_tmp_179;
  wire mux_tmp_180;
  wire and_tmp_10;
  wire or_tmp_251;
  wire mux_tmp_184;
  wire mux_tmp_195;
  wire or_tmp_254;
  wire or_tmp_255;
  wire or_tmp_277;
  wire not_tmp_156;
  wire and_dcpl_64;
  wire and_dcpl_68;
  wire and_dcpl_72;
  wire or_tmp_305;
  wire and_dcpl_73;
  wire mux_tmp_296;
  wire or_tmp_351;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire not_tmp_197;
  wire and_dcpl_78;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire mux_tmp_315;
  wire and_dcpl_86;
  wire not_tmp_208;
  wire or_tmp_398;
  wire mux_tmp_341;
  wire nor_tmp_97;
  wire and_dcpl_97;
  wire not_tmp_236;
  wire or_tmp_417;
  wire nor_tmp_103;
  wire and_dcpl_105;
  wire and_dcpl_112;
  wire and_dcpl_121;
  wire and_dcpl_123;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire mux_tmp_387;
  wire not_tmp_252;
  wire and_dcpl_127;
  wire nor_tmp_118;
  wire and_dcpl_130;
  wire and_dcpl_132;
  wire and_dcpl_139;
  wire or_tmp_523;
  wire or_tmp_524;
  wire mux_tmp_466;
  wire mux_tmp_476;
  wire not_tmp_310;
  reg exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva;
  reg VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  reg [11:0] VEC_LOOP_j_1_12_0_sva_11_0;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg modExp_exp_1_0_1_sva;
  reg [11:0] COMP_LOOP_acc_10_cse_12_1_1_sva;
  reg [10:0] COMP_LOOP_acc_psp_1_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_2_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_2_sva;
  reg [7:0] COMP_LOOP_k_9_1_1_sva_7_0;
  reg [63:0] tmp_2_lpi_4_dfm;
  reg [11:0] reg_VEC_LOOP_1_acc_1_psp_ftd_1;
  wire and_123_m1c;
  wire and_138_m1c;
  wire and_98_m1c;
  wire and_102_m1c;
  wire and_251_cse;
  wire nor_259_cse;
  reg reg_vec_rsc_triosy_0_3_obj_ld_cse;
  wire or_605_cse;
  wire and_231_cse;
  wire or_610_cse;
  wire nor_217_cse;
  wire and_230_cse;
  wire nor_161_cse;
  wire and_273_cse;
  wire or_621_cse;
  wire and_206_cse;
  wire and_187_cse;
  wire or_603_cse;
  wire and_182_cse;
  wire or_604_cse;
  wire and_224_cse;
  wire or_619_cse;
  wire and_196_cse;
  wire and_266_cse;
  wire mux_106_cse;
  wire mux_136_cse;
  wire or_298_cse;
  wire and_215_cse;
  wire or_95_cse;
  wire or_581_cse;
  wire mux_63_cse;
  wire mux_68_cse;
  wire or_280_cse;
  wire [63:0] COMP_LOOP_mux1h_1_itm_mx1;
  wire mux_96_itm;
  wire and_dcpl_150;
  wire [9:0] z_out;
  wire or_tmp_550;
  wire not_tmp_321;
  wire and_dcpl_155;
  wire and_dcpl_156;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_169;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire and_dcpl_181;
  wire and_dcpl_184;
  wire and_dcpl_187;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_195;
  wire and_dcpl_197;
  wire and_dcpl_199;
  wire [64:0] z_out_1;
  wire [10:0] z_out_2;
  wire [11:0] nl_z_out_2;
  wire [8:0] z_out_4;
  wire [9:0] nl_z_out_4;
  wire nor_tmp_146;
  wire not_tmp_368;
  wire [63:0] z_out_5;
  wire [127:0] nl_z_out_5;
  reg [63:0] p_sva;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [63:0] modExp_result_sva;
  reg modExp_exp_1_7_1_sva;
  reg modExp_exp_1_6_1_sva;
  reg modExp_exp_1_5_1_sva;
  reg modExp_exp_1_4_1_sva;
  reg modExp_exp_1_3_1_sva;
  reg modExp_exp_1_2_1_sva;
  reg modExp_exp_1_1_1_sva;
  reg modExp_exp_1_0_1_sva_1;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_mul_itm;
  reg [63:0] COMP_LOOP_mux1h_1_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [63:0] VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w5;
  wire [64:0] nl_VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w5;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire VEC_LOOP_j_1_12_0_sva_11_0_mx0c1;
  wire modExp_result_sva_mx0c0;
  wire [62:0] operator_64_false_slc_modExp_exp_63_1_3;
  wire [63:0] modulo_qr_sva_1_mx0w11;
  wire [64:0] nl_modulo_qr_sva_1_mx0w11;
  wire VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c0;
  wire VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c1;
  wire modExp_while_and_3;
  wire modExp_while_and_5;
  wire modExp_result_and_rgt;
  wire modExp_result_and_1_rgt;
  wire and_379_ssc;
  wire and_387_ssc;
  wire and_392_ssc;
  wire and_396_ssc;
  wire COMP_LOOP_or_cse;
  wire COMP_LOOP_or_1_cse;
  wire mux_462_cse;
  wire nand_86_cse;
  wire and_220_cse;
  wire or_303_cse;
  wire nor_tmp;
  wire or_tmp_586;
  wire or_tmp_598;
  wire or_tmp_600;
  wire [64:0] operator_64_false_mux1h_2_rgt;
  wire not_tmp_395;
  reg operator_64_false_acc_mut_64;
  reg [63:0] operator_64_false_acc_mut_63_0;
  wire and_226_cse;
  wire or_674_cse;
  wire COMP_LOOP_nor_3_itm;
  wire COMP_LOOP_or_24_itm;
  wire COMP_LOOP_or_25_itm;
  wire and_434_cse;

  wire[0:0] modulo_result_or_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] nor_212_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] nand_89_nl;
  wire[0:0] or_294_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] nor_213_nl;
  wire[0:0] nor_214_nl;
  wire[0:0] and_228_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] nor_215_nl;
  wire[0:0] and_284_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] nor_219_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] or_269_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] or_266_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] or_286_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] and_229_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] or_284_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] or_281_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] or_279_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] or_314_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] and_221_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] nand_101_nl;
  wire[0:0] or_308_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] or_306_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] or_304_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] mux_252_nl;
  wire[63:0] modExp_while_if_mux1h_nl;
  wire[0:0] modExp_while_if_or_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] nor_154_nl;
  wire[0:0] nor_155_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] or_588_nl;
  wire[0:0] nand_45_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] nor_156_nl;
  wire[0:0] modExp_while_if_and_nl;
  wire[0:0] modExp_while_if_and_1_nl;
  wire[0:0] and_80_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] or_628_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] nor_328_nl;
  wire[0:0] or_629_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] or_471_nl;
  wire[0:0] and_85_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] or_339_nl;
  wire[0:0] or_338_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] nor_201_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] or_474_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] nor_202_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] and_214_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] or_19_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] or_329_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] mux_530_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] or_684_nl;
  wire[0:0] and_425_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] nand_128_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] and_426_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] and_427_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] and_428_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] and_429_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] and_430_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] or_676_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] and_431_nl;
  wire[0:0] mux_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] nand_125_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] and_421_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] or_700_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] and_422_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] or_697_nl;
  wire[0:0] and_423_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] and_415_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] and_424_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] nand_118_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] mux_535_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] or_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] nand_25_nl;
  wire[0:0] or_372_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] and_417_nl;
  wire[0:0] mux_551_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] and_418_nl;
  wire[0:0] and_419_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] and_100_nl;
  wire[0:0] r_or_nl;
  wire[0:0] r_or_1_nl;
  wire[0:0] and_105_nl;
  wire[0:0] and_107_nl;
  wire[0:0] and_109_nl;
  wire[0:0] and_111_nl;
  wire[0:0] nor_301_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nand_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] nor_302_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] or_620_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] or_32_nl;
  wire[0:0] or_30_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] or_593_nl;
  wire[0:0] or_594_nl;
  wire[0:0] nand_51_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] nand_52_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] or_595_nl;
  wire[0:0] nand_53_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] nand_54_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] nand_55_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] nor_181_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] nor_182_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] or_426_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] or_424_nl;
  wire[0:0] or_104_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] nand_87_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] or_418_nl;
  wire[0:0] COMP_LOOP_or_3_nl;
  wire[0:0] COMP_LOOP_or_4_nl;
  wire[0:0] COMP_LOOP_or_5_nl;
  wire[0:0] COMP_LOOP_or_6_nl;
  wire[0:0] mux_379_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] and_189_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] nor_174_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] nor_175_nl;
  wire[0:0] and_191_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] or_440_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] COMP_LOOP_mux1h_11_nl;
  wire[0:0] COMP_LOOP_and_11_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] and_288_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] or_592_nl;
  wire[0:0] nor_165_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] nor_167_nl;
  wire[0:0] and_186_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] mux_393_nl;
  wire[0:0] or_463_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] nor_168_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] or_459_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] or_458_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] or_457_nl;
  wire[0:0] or_455_nl;
  wire[0:0] nand_49_nl;
  wire[9:0] VEC_LOOP_1_COMP_LOOP_1_acc_11_nl;
  wire[10:0] nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl;
  wire[0:0] nor_330_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] or_506_nl;
  wire[0:0] or_505_nl;
  wire[0:0] or_504_nl;
  wire[0:0] nor_331_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] or_501_nl;
  wire[0:0] or_499_nl;
  wire[11:0] COMP_LOOP_mux_88_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] and_175_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] and_177_nl;
  wire[0:0] and_179_nl;
  wire[0:0] nor_146_nl;
  wire[0:0] nor_147_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] and_172_nl;
  wire[0:0] nor_148_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] or_544_nl;
  wire[0:0] or_542_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] nor_326_nl;
  wire[0:0] and_286_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] or_538_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] and_287_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] nor_316_nl;
  wire[0:0] nor_317_nl;
  wire[0:0] nor_318_nl;
  wire[0:0] and_283_nl;
  wire[0:0] COMP_LOOP_mux1h_20_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] nand_38_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] or_558_nl;
  wire[0:0] mux_473_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] and_162_nl;
  wire[0:0] or_556_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] or_555_nl;
  wire[0:0] COMP_LOOP_mux1h_37_nl;
  wire[0:0] nor_277_nl;
  wire[0:0] and_18_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] and_17_nl;
  wire[0:0] or_135_nl;
  wire[0:0] or_133_nl;
  wire[0:0] or_145_nl;
  wire[0:0] or_143_nl;
  wire[0:0] nor_242_nl;
  wire[0:0] nor_243_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] or_271_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] and_216_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] and_217_nl;
  wire[0:0] nor_208_nl;
  wire[0:0] and_218_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] or_626_nl;
  wire[0:0] or_627_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] nor_205_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] nor_203_nl;
  wire[0:0] nor_204_nl;
  wire[0:0] or_373_nl;
  wire[0:0] or_392_nl;
  wire[0:0] or_390_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] nor_275_nl;
  wire[0:0] nor_276_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] mux_317_nl;
  wire[0:0] or_607_nl;
  wire[0:0] nand_74_nl;
  wire[0:0] or_396_nl;
  wire[0:0] nor_186_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] or_407_nl;
  wire[0:0] or_406_nl;
  wire[0:0] nor_187_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] or_403_nl;
  wire[0:0] or_401_nl;
  wire[0:0] nor_178_nl;
  wire[0:0] nor_179_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] nor_173_nl;
  wire[0:0] and_188_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] nor_171_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] or_452_nl;
  wire[0:0] or_451_nl;
  wire[0:0] nor_172_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] or_552_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] nand_73_nl;
  wire[0:0] nand_40_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] mux_491_nl;
  wire[0:0] nand_37_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] and_168_nl;
  wire[0:0] nor_143_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] mux_486_nl;
  wire[0:0] mux_485_nl;
  wire[0:0] nor_144_nl;
  wire[0:0] nor_145_nl;
  wire[0:0] mux_484_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] mux_482_nl;
  wire[0:0] nor_190_nl;
  wire[0:0] and_94_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] or_394_nl;
  wire[0:0] and_49_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] nor_273_nl;
  wire[0:0] nor_274_nl;
  wire[0:0] mux_101_nl;
  wire[0:0] and_253_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] nor_270_nl;
  wire[0:0] nor_271_nl;
  wire[0:0] nor_272_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] or_124_nl;
  wire[0:0] or_122_nl;
  wire[0:0] and_51_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] nor_268_nl;
  wire[0:0] nor_269_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] and_252_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] nor_263_nl;
  wire[0:0] nor_264_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] nor_265_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] or_150_nl;
  wire[0:0] or_149_nl;
  wire[0:0] nor_266_nl;
  wire[0:0] nor_267_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] or_140_nl;
  wire[0:0] or_138_nl;
  wire[0:0] and_250_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] nor_256_nl;
  wire[0:0] nor_257_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] nor_258_nl;
  wire[0:0] nor_260_nl;
  wire[0:0] or_160_nl;
  wire[0:0] nor_261_nl;
  wire[0:0] nor_262_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] or_157_nl;
  wire[0:0] or_156_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] and_249_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] nor_251_nl;
  wire[0:0] nor_252_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] nor_253_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] or_184_nl;
  wire[0:0] or_183_nl;
  wire[0:0] nor_254_nl;
  wire[0:0] nor_255_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] or_174_nl;
  wire[0:0] or_172_nl;
  wire[0:0] and_246_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] nor_245_nl;
  wire[0:0] and_247_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] nor_246_nl;
  wire[0:0] nor_248_nl;
  wire[0:0] or_195_nl;
  wire[0:0] nor_249_nl;
  wire[0:0] nor_250_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] or_192_nl;
  wire[0:0] or_190_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] and_244_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] nor_239_nl;
  wire[0:0] nor_240_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] nor_241_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] or_216_nl;
  wire[0:0] or_215_nl;
  wire[0:0] and_245_nl;
  wire[0:0] nor_244_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] or_209_nl;
  wire[0:0] or_207_nl;
  wire[0:0] and_241_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] nor_233_nl;
  wire[0:0] and_242_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] nor_234_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] nor_235_nl;
  wire[0:0] nor_45_nl;
  wire[0:0] nor_237_nl;
  wire[0:0] nor_238_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] or_223_nl;
  wire[0:0] or_222_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] and_238_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] nor_226_nl;
  wire[0:0] nor_227_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] nor_228_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] nor_229_nl;
  wire[0:0] and_239_nl;
  wire[0:0] nor_232_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] or_239_nl;
  wire[0:0] nand_90_nl;
  wire[0:0] and_234_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] nor_220_nl;
  wire[0:0] and_235_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] nor_221_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] nor_222_nl;
  wire[0:0] and_237_nl;
  wire[0:0] nor_224_nl;
  wire[0:0] nor_225_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] or_253_nl;
  wire[0:0] nand_64_nl;
  wire[0:0] nor_343_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] or_642_nl;
  wire[0:0] nor_344_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] or_638_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] nor_nl;
  wire[0:0] mux_503_nl;
  wire[0:0] nor_352_nl;
  wire[0:0] nor_353_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] nand_112_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] or_708_nl;
  wire[0:0] nand_127_nl;
  wire[0:0] and_420_nl;
  wire[0:0] nor_388_nl;
  wire[10:0] acc_nl;
  wire[11:0] nl_acc_nl;
  wire[9:0] COMP_LOOP_mux_85_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nand_1_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] nor_401_nl;
  wire[65:0] acc_1_nl;
  wire[66:0] nl_acc_1_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_53_nl;
  wire[0:0] COMP_LOOP_mux_86_nl;
  wire[50:0] COMP_LOOP_or_32_nl;
  wire[50:0] COMP_LOOP_and_70_nl;
  wire[50:0] COMP_LOOP_mux1h_67_nl;
  wire[1:0] COMP_LOOP_or_33_nl;
  wire[1:0] COMP_LOOP_and_71_nl;
  wire[1:0] COMP_LOOP_mux1h_68_nl;
  wire[0:0] COMP_LOOP_nor_59_nl;
  wire[9:0] COMP_LOOP_mux1h_69_nl;
  wire[8:0] COMP_LOOP_acc_33_nl;
  wire[9:0] nl_COMP_LOOP_acc_33_nl;
  wire[0:0] COMP_LOOP_or_34_nl;
  wire[0:0] COMP_LOOP_or_35_nl;
  wire[0:0] COMP_LOOP_or_36_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_54_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_55_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_56_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_57_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_58_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_59_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_60_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_61_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_62_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_63_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_64_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_65_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_66_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_67_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_68_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_69_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_70_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_71_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_72_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_73_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_74_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_75_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_76_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_77_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_78_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_79_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_80_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_81_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_82_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_83_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_84_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_85_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_86_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_87_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_88_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_89_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_90_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_91_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_92_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_93_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_94_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_95_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_96_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_97_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_98_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_99_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_100_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_101_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_102_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_103_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_104_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_105_nl;
  wire[1:0] COMP_LOOP_or_37_nl;
  wire[1:0] COMP_LOOP_and_72_nl;
  wire[1:0] COMP_LOOP_mux1h_70_nl;
  wire[0:0] COMP_LOOP_nor_61_nl;
  wire[9:0] COMP_LOOP_or_38_nl;
  wire[9:0] COMP_LOOP_mux1h_71_nl;
  wire[0:0] COMP_LOOP_or_39_nl;
  wire[0:0] COMP_LOOP_or_40_nl;
  wire[10:0] COMP_LOOP_mux_87_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_1_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_nor_4_nl;
  wire[0:0] operator_64_false_1_mux1h_9_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_nor_5_nl;
  wire[0:0] operator_64_false_1_mux1h_10_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_nor_6_nl;
  wire[0:0] operator_64_false_1_mux1h_11_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_nor_7_nl;
  wire[0:0] operator_64_false_1_mux1h_12_nl;
  wire[0:0] operator_64_false_1_mux1h_13_nl;
  wire[0:0] operator_64_false_1_mux1h_14_nl;
  wire[0:0] operator_64_false_1_mux1h_15_nl;
  wire[0:0] operator_64_false_1_mux1h_16_nl;
  wire[0:0] operator_64_false_1_or_2_nl;
  wire[63:0] modExp_while_if_mux1h_2_nl;
  wire[0:0] and_436_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] nand_129_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] or_713_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] or_714_nl;
  wire[0:0] or_715_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] mux_564_nl;
  wire[0:0] or_716_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] or_717_nl;
  wire[0:0] or_718_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] and_437_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_operator_66_true_div_cmp_b;
  assign nl_operator_66_true_div_cmp_b = {1'b0, operator_66_true_div_cmp_b_9_0};
  wire[64:0] operator_64_false_acc_1_nl;
  wire[65:0] nl_operator_64_false_acc_1_nl;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0;
  assign nl_operator_64_false_acc_1_nl = ({1'b1 , (~ (operator_66_true_div_cmp_z[63:0]))})
      + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_acc_1_nl = nl_operator_64_false_acc_1_nl[64:0];
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 = ~ (readslicef_65_1_64(operator_64_false_acc_1_nl));
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0 = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_62_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_62_tr0 = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_1[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0 = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_62_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_62_tr0 = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0 = z_out_1[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 = ~ (z_out_1[2]);
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd1)) modulo_result_rem_cmp (
      .a(modulo_result_rem_cmp_a),
      .b(modulo_result_rem_cmp_b),
      .z(modulo_result_rem_cmp_z)
    );
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(nl_operator_66_true_div_cmp_b[10:0]),
      .z(operator_66_true_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_8_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0[0:0]),
      .modExp_while_C_38_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_1_COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_1_COMP_LOOP_C_62_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_62_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_C_124_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_2_COMP_LOOP_C_62_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_62_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_C_124_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0[0:0]),
      .STAGE_LOOP_C_9_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0[0:0])
    );
  assign and_251_cse = (fsm_output[2]) & (fsm_output[7]) & (fsm_output[4]) & (~ (fsm_output[8]));
  assign nor_259_cse = ~((~ (fsm_output[5])) | (fsm_output[2]) | (fsm_output[7])
      | (fsm_output[4]) | (~ (fsm_output[8])));
  assign or_605_cse = (fsm_output[1:0]!=2'b00);
  assign and_231_cse = (fsm_output[1:0]==2'b11);
  assign or_603_cse = (fsm_output[4:3]!=2'b00);
  assign nor_217_cse = ~((fsm_output[2:1]!=2'b00));
  assign and_230_cse = (fsm_output[2:0]==3'b111);
  assign or_604_cse = (fsm_output[3]) | (fsm_output[7]);
  assign and_224_cse = (fsm_output[3]) & (fsm_output[7]);
  assign or_298_cse = (fsm_output[7:6]!=2'b00);
  assign or_280_cse = and_231_cse | (fsm_output[2]);
  assign and_220_cse = (fsm_output[3]) & (fsm_output[7]) & (fsm_output[6]);
  assign or_303_cse = (fsm_output[3]) | (fsm_output[7]) | (fsm_output[6]);
  assign and_226_cse = (fsm_output[1]) & (fsm_output[3]);
  assign or_610_cse = (fsm_output[5:4]!=2'b00);
  assign and_215_cse = (fsm_output[8:6]==3'b111);
  assign nor_161_cse = ~((fsm_output[1:0]!=2'b00));
  assign and_182_cse = (fsm_output[8:7]==2'b11);
  assign nor_154_nl = ~((~ (fsm_output[8])) | (fsm_output[3]) | (fsm_output[7]) |
      (fsm_output[1]) | (~ nor_tmp_118));
  assign or_588_nl = (fsm_output[7]) | (~ (fsm_output[1])) | (~ (fsm_output[5]))
      | (fsm_output[2]) | (fsm_output[6]);
  assign nor_156_nl = ~((fsm_output[5]) | (fsm_output[2]) | (fsm_output[6]));
  assign mux_429_nl = MUX_s_1_2_2(nor_156_nl, nor_tmp_118, fsm_output[1]);
  assign nand_45_nl = ~((fsm_output[7]) & mux_429_nl);
  assign mux_430_nl = MUX_s_1_2_2(or_588_nl, nand_45_nl, fsm_output[3]);
  assign nor_155_nl = ~((fsm_output[8]) | mux_430_nl);
  assign mux_431_nl = MUX_s_1_2_2(nor_154_nl, nor_155_nl, fsm_output[4]);
  assign modExp_while_if_or_nl = and_dcpl_62 | (mux_431_nl & modExp_exp_1_0_1_sva
      & (fsm_output[0]));
  assign modExp_while_if_and_nl = modExp_while_and_3 & and_dcpl_125;
  assign modExp_while_if_and_1_nl = modExp_while_and_5 & and_dcpl_125;
  assign modExp_while_if_mux1h_nl = MUX1HOT_v_64_5_2(z_out_5, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w11, (z_out_1[63:0]), {modExp_while_if_or_nl
      , and_dcpl_86 , modExp_while_if_and_nl , modExp_while_if_and_1_nl , not_tmp_156});
  assign and_80_nl = and_dcpl_15 & and_dcpl_24;
  assign or_628_nl = (fsm_output[4]) | (fsm_output[8]);
  assign nor_328_nl = ~(nor_217_cse | (fsm_output[8]));
  assign mux_269_nl = MUX_s_1_2_2((fsm_output[8]), nor_328_nl, fsm_output[4]);
  assign mux_270_nl = MUX_s_1_2_2(or_628_nl, mux_269_nl, fsm_output[5]);
  assign or_629_nl = (fsm_output[5:4]!=2'b10) | (or_280_cse & (fsm_output[8]));
  assign mux_271_nl = MUX_s_1_2_2(mux_270_nl, or_629_nl, fsm_output[6]);
  assign or_471_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[8]);
  assign mux_266_nl = MUX_s_1_2_2(or_471_nl, or_tmp_305, fsm_output[4]);
  assign and_85_nl = (fsm_output[4]) & (and_231_cse | (fsm_output[2]) | (~ (fsm_output[8])));
  assign mux_267_nl = MUX_s_1_2_2(mux_266_nl, and_85_nl, fsm_output[5]);
  assign or_339_nl = (~ (fsm_output[4])) | (~ (fsm_output[2])) | (fsm_output[8]);
  assign or_338_nl = (fsm_output[4]) | and_230_cse | (fsm_output[8]);
  assign mux_265_nl = MUX_s_1_2_2(or_339_nl, or_338_nl, fsm_output[5]);
  assign mux_268_nl = MUX_s_1_2_2(mux_267_nl, mux_265_nl, fsm_output[6]);
  assign mux_272_nl = MUX_s_1_2_2(mux_271_nl, mux_268_nl, fsm_output[3]);
  assign nor_201_nl = ~((fsm_output[5]) | (~((fsm_output[4]) & (((~((fsm_output[1:0]==2'b11)))
      & (fsm_output[2])) | (fsm_output[8])))));
  assign or_474_nl = (fsm_output[2]) | (~ (fsm_output[8]));
  assign mux_260_nl = MUX_s_1_2_2((~ or_tmp_305), or_474_nl, or_605_cse);
  assign mux_261_nl = MUX_s_1_2_2(mux_260_nl, or_tmp_305, fsm_output[4]);
  assign mux_262_nl = MUX_s_1_2_2(mux_261_nl, (fsm_output[8]), fsm_output[5]);
  assign mux_263_nl = MUX_s_1_2_2(nor_201_nl, mux_262_nl, fsm_output[6]);
  assign and_214_nl = or_605_cse & (fsm_output[2]) & (fsm_output[8]);
  assign mux_258_nl = MUX_s_1_2_2(and_214_nl, (fsm_output[8]), fsm_output[4]);
  assign nor_202_nl = ~((fsm_output[5]) | (~ mux_258_nl));
  assign or_19_nl = (~ (fsm_output[4])) | (fsm_output[8]);
  assign or_329_nl = (fsm_output[0]) | (fsm_output[2]) | (fsm_output[8]);
  assign mux_255_nl = MUX_s_1_2_2(or_329_nl, or_tmp_305, fsm_output[1]);
  assign mux_256_nl = MUX_s_1_2_2((fsm_output[8]), mux_255_nl, fsm_output[4]);
  assign mux_257_nl = MUX_s_1_2_2(or_19_nl, mux_256_nl, fsm_output[5]);
  assign mux_259_nl = MUX_s_1_2_2(nor_202_nl, mux_257_nl, fsm_output[6]);
  assign mux_264_nl = MUX_s_1_2_2(mux_263_nl, mux_259_nl, fsm_output[3]);
  assign mux_273_nl = MUX_s_1_2_2(mux_272_nl, (~ mux_264_nl), fsm_output[7]);
  assign operator_64_false_mux1h_2_rgt = MUX1HOT_v_65_3_2(z_out_1, ({2'b00 , operator_64_false_slc_modExp_exp_63_1_3}),
      ({1'b0 , modExp_while_if_mux1h_nl}), {and_80_nl , and_dcpl_72 , mux_273_nl});
  assign or_674_cse = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[3]);
  assign and_206_cse = (fsm_output[5:4]==2'b11);
  assign and_98_m1c = and_dcpl_33 & (fsm_output[2]) & and_dcpl_12 & and_dcpl_78;
  assign modExp_result_and_rgt = (~ modExp_while_and_5) & and_98_m1c;
  assign modExp_result_and_1_rgt = modExp_while_and_5 & and_98_m1c;
  assign and_196_cse = (fsm_output[0]) & (fsm_output[3]);
  assign or_95_cse = (fsm_output[4]) | (fsm_output[7]);
  assign mux_63_cse = MUX_s_1_2_2((~ or_604_cse), (fsm_output[7]), fsm_output[4]);
  assign mux_68_cse = MUX_s_1_2_2(or_95_cse, or_tmp_69, fsm_output[5]);
  assign or_621_cse = (fsm_output[3:2]!=2'b00);
  assign and_273_cse = (fsm_output[2:1]==2'b11);
  assign and_187_cse = (fsm_output[5]) & (fsm_output[1]) & (fsm_output[2]);
  assign or_619_cse = (fsm_output[2:1]!=2'b00);
  assign COMP_LOOP_or_cse = (and_dcpl_27 & and_dcpl_24) | (and_dcpl_44 & and_dcpl_12
      & and_dcpl_19);
  assign and_266_cse = (fsm_output[7:6]==2'b11);
  assign nor_146_nl = ~((fsm_output[5]) | (fsm_output[4]) | (~ (fsm_output[8])));
  assign nor_147_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_462_cse = MUX_s_1_2_2(nor_146_nl, nor_147_nl, fsm_output[2]);
  assign COMP_LOOP_or_1_cse = (and_dcpl_33 & (~ (fsm_output[2])) & and_dcpl_32 &
      (fsm_output[7:6]==2'b01) & and_dcpl_29) | (and_dcpl_45 & and_dcpl_43) | ((fsm_output[5])
      & (~ (fsm_output[4])) & (fsm_output[2]) & and_dcpl_49 & and_dcpl_11) | (and_dcpl_14
      & and_dcpl_49 & and_dcpl_43);
  assign nl_VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w5 = tmp_2_lpi_4_dfm + COMP_LOOP_mux1h_1_itm_mx1;
  assign VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w5 = nl_VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w5[63:0];
  assign operator_64_false_slc_modExp_exp_63_1_3 = MUX_v_63_2_2((operator_66_true_div_cmp_z[63:1]),
      (tmp_2_lpi_4_dfm[63:1]), and_dcpl_82);
  assign nl_modulo_qr_sva_1_mx0w11 = modulo_result_rem_cmp_z + p_sva;
  assign modulo_qr_sva_1_mx0w11 = nl_modulo_qr_sva_1_mx0w11[63:0];
  assign COMP_LOOP_mux1h_1_itm_mx1 = MUX_v_64_2_2(modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w11,
      modulo_result_rem_cmp_z[63]);
  assign modExp_while_and_3 = (~ (modulo_result_rem_cmp_z[63])) & modExp_exp_1_0_1_sva;
  assign modExp_while_and_5 = (modulo_result_rem_cmp_z[63]) & modExp_exp_1_0_1_sva;
  assign not_tmp_20 = ~((fsm_output[0]) & (fsm_output[7]));
  assign not_tmp_38 = ~((fsm_output[8:7]!=2'b00));
  assign mux_tmp_40 = MUX_s_1_2_2(not_tmp_38, and_182_cse, fsm_output[6]);
  assign or_tmp_69 = (~ (fsm_output[4])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_tmp_93 = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[5]);
  assign and_tmp_7 = (fsm_output[8:6]==3'b111) & or_tmp_93;
  assign nor_277_nl = ~((fsm_output[6]) | (fsm_output[8]) | (fsm_output[1]) | (fsm_output[2])
      | (fsm_output[4]) | (fsm_output[5]));
  assign and_18_nl = (fsm_output[6]) & (fsm_output[8]) & or_610_cse;
  assign mux_tmp_94 = MUX_s_1_2_2(nor_277_nl, and_18_nl, fsm_output[7]);
  assign mux_tmp_95 = MUX_s_1_2_2(mux_tmp_94, and_tmp_7, fsm_output[3]);
  assign and_17_nl = (fsm_output[8:6]==3'b111) & or_610_cse;
  assign mux_93_nl = MUX_s_1_2_2(and_17_nl, and_tmp_7, fsm_output[3]);
  assign mux_96_itm = MUX_s_1_2_2(mux_tmp_95, mux_93_nl, fsm_output[0]);
  assign and_dcpl_10 = ~((fsm_output[7:6]!=2'b00));
  assign and_dcpl_11 = and_dcpl_10 & (~ (fsm_output[3])) & (~ (fsm_output[0]));
  assign and_dcpl_12 = ~((fsm_output[1]) | (fsm_output[8]));
  assign and_dcpl_13 = ~((fsm_output[5:4]!=2'b00));
  assign and_dcpl_14 = and_dcpl_13 & (~ (fsm_output[2]));
  assign and_dcpl_15 = and_dcpl_14 & and_dcpl_12;
  assign and_dcpl_19 = and_266_cse & and_196_cse;
  assign and_dcpl_21 = and_dcpl_14 & (~ (fsm_output[1])) & (fsm_output[8]);
  assign and_dcpl_23 = (~ (fsm_output[3])) & (fsm_output[0]);
  assign and_dcpl_24 = and_dcpl_10 & and_dcpl_23;
  assign and_dcpl_26 = and_206_cse & (~ (fsm_output[2]));
  assign and_dcpl_27 = and_dcpl_26 & and_dcpl_12;
  assign and_dcpl_29 = (fsm_output[3]) & (~ (fsm_output[0]));
  assign and_dcpl_32 = (fsm_output[1]) & (~ (fsm_output[8]));
  assign and_dcpl_33 = (fsm_output[5:4]==2'b01);
  assign and_dcpl_37 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_40 = (fsm_output[1]) & (~ (fsm_output[3]));
  assign or_135_nl = (~ (fsm_output[6])) | (~ (fsm_output[8])) | (fsm_output[2])
      | (fsm_output[4]) | (~ (fsm_output[5]));
  assign or_133_nl = (fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[2])) | (~
      (fsm_output[4])) | (fsm_output[5]);
  assign mux_tmp_103 = MUX_s_1_2_2(or_135_nl, or_133_nl, fsm_output[7]);
  assign and_dcpl_42 = (fsm_output[7:6]==2'b10);
  assign and_dcpl_43 = and_dcpl_42 & and_196_cse;
  assign and_dcpl_44 = and_206_cse & (fsm_output[2]);
  assign and_dcpl_45 = and_dcpl_44 & and_dcpl_32;
  assign and_dcpl_49 = (fsm_output[1]) & (fsm_output[8]);
  assign not_tmp_92 = ~((fsm_output[8]) & (fsm_output[6]));
  assign or_145_nl = (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign or_143_nl = (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[6]);
  assign mux_106_cse = MUX_s_1_2_2(or_145_nl, or_143_nl, fsm_output[4]);
  assign not_tmp_109 = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[1]) & (fsm_output[8]) &
      (fsm_output[6]));
  assign nor_242_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[6])));
  assign nor_243_nl = ~((fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[6]));
  assign mux_136_cse = MUX_s_1_2_2(nor_242_nl, nor_243_nl, fsm_output[4]);
  assign nor_tmp_48 = (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b11) & (fsm_output[8])
      & (fsm_output[6]);
  assign and_dcpl_62 = and_dcpl_14 & and_dcpl_32 & and_dcpl_10 & and_dcpl_29;
  assign or_tmp_242 = (fsm_output[3]) | (fsm_output[8]);
  assign nor_tmp_51 = (fsm_output[3]) & (fsm_output[8]);
  assign or_tmp_244 = (~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[8]);
  assign mux_167_nl = MUX_s_1_2_2((~ nor_tmp_51), or_tmp_242, fsm_output[7]);
  assign mux_tmp_168 = MUX_s_1_2_2(or_tmp_244, mux_167_nl, fsm_output[4]);
  assign or_tmp_245 = (fsm_output[8:7]!=2'b10);
  assign or_tmp_247 = (~ (fsm_output[3])) | (fsm_output[8]);
  assign mux_tmp_174 = MUX_s_1_2_2((~ or_tmp_242), nor_tmp_51, fsm_output[7]);
  assign or_271_nl = (fsm_output[7]) | (fsm_output[3]) | (fsm_output[8]);
  assign mux_tmp_175 = MUX_s_1_2_2(mux_tmp_174, or_271_nl, fsm_output[4]);
  assign or_tmp_249 = (fsm_output[3]) | (~ (fsm_output[8]));
  assign mux_178_nl = MUX_s_1_2_2(or_tmp_242, or_tmp_249, fsm_output[7]);
  assign mux_tmp_179 = MUX_s_1_2_2(mux_178_nl, or_tmp_245, fsm_output[4]);
  assign mux_tmp_180 = MUX_s_1_2_2(mux_tmp_179, mux_tmp_168, fsm_output[5]);
  assign mux_182_nl = MUX_s_1_2_2((~ or_tmp_247), or_tmp_249, fsm_output[7]);
  assign and_tmp_10 = (fsm_output[4]) & mux_182_nl;
  assign or_tmp_251 = and_224_cse | (fsm_output[8]);
  assign mux_tmp_184 = MUX_s_1_2_2(mux_tmp_174, or_tmp_251, fsm_output[4]);
  assign mux_tmp_195 = MUX_s_1_2_2((~ nor_tmp_51), (fsm_output[8]), fsm_output[7]);
  assign or_tmp_254 = (fsm_output[7:6]!=2'b10);
  assign or_tmp_255 = (fsm_output[7:6]!=2'b01);
  assign or_tmp_277 = (~((fsm_output[3]) | (fsm_output[7]))) | (fsm_output[6]);
  assign and_217_nl = (fsm_output[4]) & (fsm_output[2]) & (fsm_output[6]) & (~ (fsm_output[8]));
  assign nor_208_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[6]) | (~
      (fsm_output[8])));
  assign mux_247_nl = MUX_s_1_2_2(and_217_nl, nor_208_nl, fsm_output[5]);
  assign and_216_nl = (~((fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[7]))))
      & mux_247_nl;
  assign and_218_nl = (fsm_output[1]) & (fsm_output[3]) & (~ (fsm_output[7])) & (fsm_output[5])
      & mux_136_cse;
  assign not_tmp_156 = MUX_s_1_2_2(and_216_nl, and_218_nl, fsm_output[0]);
  assign or_626_nl = (fsm_output[7]) | (~ (fsm_output[6])) | (~ (fsm_output[8]))
      | (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[5]));
  assign or_627_nl = (~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[2])
      | (~ (fsm_output[4])) | (fsm_output[5]);
  assign mux_249_nl = MUX_s_1_2_2(or_626_nl, or_627_nl, fsm_output[3]);
  assign and_dcpl_64 = ~(mux_249_nl | (fsm_output[1:0]!=2'b00));
  assign mux_250_nl = MUX_s_1_2_2(or_619_cse, (~ or_619_cse), fsm_output[3]);
  assign nor_205_nl = ~((fsm_output[3]) | (~ or_619_cse));
  assign mux_251_nl = MUX_s_1_2_2(mux_250_nl, nor_205_nl, fsm_output[0]);
  assign and_dcpl_68 = mux_251_nl & (~ (fsm_output[5])) & (~ (fsm_output[4])) & (~
      (fsm_output[8])) & and_dcpl_10;
  assign nor_203_nl = ~((fsm_output[3]) | (~ and_206_cse));
  assign nor_204_nl = ~((fsm_output[5:3]!=3'b001));
  assign mux_254_nl = MUX_s_1_2_2(nor_203_nl, nor_204_nl, fsm_output[0]);
  assign and_dcpl_72 = mux_254_nl & (~ (fsm_output[2])) & and_dcpl_12 & and_dcpl_10;
  assign or_tmp_305 = (~ (fsm_output[2])) | (fsm_output[8]);
  assign and_dcpl_73 = and_266_cse & and_dcpl_29;
  assign or_373_nl = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[5]);
  assign mux_tmp_296 = MUX_s_1_2_2((~ and_dcpl_44), or_373_nl, fsm_output[8]);
  assign or_tmp_351 = (fsm_output[7]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[2])
      | (~ and_206_cse);
  assign and_dcpl_76 = (~ mux_tmp_296) & (fsm_output[1]);
  assign and_dcpl_77 = and_dcpl_76 & and_dcpl_43;
  assign not_tmp_197 = ~((fsm_output[8:6]!=3'b000));
  assign and_dcpl_78 = and_dcpl_10 & and_196_cse;
  assign and_dcpl_82 = and_dcpl_27 & and_dcpl_11;
  assign and_dcpl_84 = ~((fsm_output[1]) | (fsm_output[7]));
  assign or_392_nl = (fsm_output[6]) | (~ (fsm_output[8])) | (~ (fsm_output[2]))
      | (fsm_output[4]) | (~ (fsm_output[5]));
  assign or_390_nl = (~ (fsm_output[6])) | (fsm_output[8]) | (fsm_output[2]) | (~
      (fsm_output[4])) | (fsm_output[5]);
  assign mux_tmp_315 = MUX_s_1_2_2(or_392_nl, or_390_nl, fsm_output[3]);
  assign nor_275_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[0])) | (~ (fsm_output[6]))
      | (fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[2]) | (fsm_output[7]));
  assign or_607_nl = (fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[2]) | (fsm_output[7]);
  assign nand_74_nl = ~((fsm_output[3]) & (fsm_output[5]) & (fsm_output[2]) & (fsm_output[7]));
  assign mux_317_nl = MUX_s_1_2_2(or_607_nl, nand_74_nl, fsm_output[6]);
  assign or_396_nl = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[5]) | (~((fsm_output[2])
      & (fsm_output[7])));
  assign mux_318_nl = MUX_s_1_2_2(mux_317_nl, or_396_nl, fsm_output[0]);
  assign nor_276_nl = ~((fsm_output[8]) | mux_318_nl);
  assign mux_319_nl = MUX_s_1_2_2(nor_275_nl, nor_276_nl, fsm_output[4]);
  assign and_dcpl_86 = mux_319_nl & (fsm_output[1]);
  assign or_407_nl = (~ (fsm_output[6])) | (fsm_output[8]) | (fsm_output[3]);
  assign or_406_nl = (fsm_output[6]) | (~((fsm_output[8]) & (fsm_output[3])));
  assign mux_321_nl = MUX_s_1_2_2(or_407_nl, or_406_nl, fsm_output[2]);
  assign nor_186_nl = ~((fsm_output[1]) | (~ (fsm_output[7])) | (fsm_output[5]) |
      (fsm_output[4]) | mux_321_nl);
  assign or_403_nl = (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[6]))
      | (fsm_output[8]) | (~ (fsm_output[3]));
  assign or_401_nl = (fsm_output[4]) | (~ (fsm_output[2])) | (fsm_output[6]) | (~
      (fsm_output[8])) | (fsm_output[3]);
  assign mux_320_nl = MUX_s_1_2_2(or_403_nl, or_401_nl, fsm_output[5]);
  assign nor_187_nl = ~((~ (fsm_output[1])) | (fsm_output[7]) | mux_320_nl);
  assign not_tmp_208 = MUX_s_1_2_2(nor_186_nl, nor_187_nl, fsm_output[0]);
  assign nand_86_cse = ~((fsm_output[0]) & (fsm_output[3]));
  assign or_tmp_398 = ~(nand_86_cse & (fsm_output[7]));
  assign mux_tmp_341 = MUX_s_1_2_2(and_224_cse, or_604_cse, fsm_output[0]);
  assign nor_tmp_97 = or_603_cse & (fsm_output[7]);
  assign and_dcpl_97 = (fsm_output[5]) & (fsm_output[1]);
  assign nor_178_nl = ~((fsm_output[7]) | (~((fsm_output[6]) & (fsm_output[8]) &
      (fsm_output[2]) & (fsm_output[4]))));
  assign nor_179_nl = ~((~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[8]) |
      (fsm_output[2]) | (fsm_output[4]));
  assign not_tmp_236 = MUX_s_1_2_2(nor_178_nl, nor_179_nl, fsm_output[3]);
  assign or_tmp_417 = (fsm_output[7]) | (~ (fsm_output[4]));
  assign nor_tmp_103 = (fsm_output[7]) & (fsm_output[4]);
  assign and_dcpl_105 = (fsm_output[1]) & (~ (COMP_LOOP_acc_1_cse_2_sva[1]));
  assign and_dcpl_112 = (fsm_output[1]) & (COMP_LOOP_acc_1_cse_2_sva[1]);
  assign and_dcpl_121 = (fsm_output[4]) & (fsm_output[1]);
  assign nor_173_nl = ~((fsm_output[7]) | (fsm_output[6]) | (fsm_output[2]));
  assign and_188_nl = (fsm_output[7]) & (fsm_output[6]) & (fsm_output[2]);
  assign mux_381_nl = MUX_s_1_2_2(nor_173_nl, and_188_nl, fsm_output[3]);
  assign and_dcpl_123 = mux_381_nl & (fsm_output[5]);
  assign and_dcpl_124 = and_dcpl_123 & and_dcpl_121 & (~ (fsm_output[8])) & (~ (fsm_output[0]));
  assign or_452_nl = (~ (fsm_output[8])) | (fsm_output[2]) | (~ (fsm_output[4]))
      | (fsm_output[5]);
  assign or_451_nl = (fsm_output[8]) | (~ (fsm_output[2])) | (fsm_output[4]) | (fsm_output[5]);
  assign mux_382_nl = MUX_s_1_2_2(or_452_nl, or_451_nl, fsm_output[6]);
  assign nor_171_nl = ~((fsm_output[7]) | mux_382_nl);
  assign nor_172_nl = ~((fsm_output[7:6]!=2'b10) | mux_tmp_296);
  assign mux_383_nl = MUX_s_1_2_2(nor_171_nl, nor_172_nl, fsm_output[3]);
  assign and_dcpl_125 = mux_383_nl & and_dcpl_37;
  assign mux_tmp_387 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[5]);
  assign not_tmp_252 = ~((fsm_output[1]) | (fsm_output[2]) | (fsm_output[8]));
  assign and_dcpl_127 = (~ mux_tmp_103) & and_dcpl_40 & (fsm_output[0]);
  assign nor_tmp_118 = (fsm_output[5]) & (fsm_output[2]) & (fsm_output[6]);
  assign and_dcpl_130 = (~ (fsm_output[8])) & (fsm_output[0]);
  assign and_dcpl_132 = and_dcpl_123 & and_dcpl_121 & and_dcpl_130;
  assign or_552_nl = (~ (fsm_output[3])) | (~ (fsm_output[7])) | (fsm_output[6])
      | mux_tmp_296;
  assign nand_73_nl = ~((fsm_output[8:6]==3'b011) & and_dcpl_44);
  assign mux_464_nl = MUX_s_1_2_2(or_tmp_351, nand_73_nl, fsm_output[3]);
  assign mux_465_nl = MUX_s_1_2_2(or_552_nl, mux_464_nl, fsm_output[0]);
  assign and_dcpl_139 = (~ mux_465_nl) & (fsm_output[1]);
  assign or_tmp_523 = (fsm_output[7]) | (~ (fsm_output[5]));
  assign or_tmp_524 = (fsm_output[7]) | (fsm_output[5]);
  assign mux_tmp_466 = MUX_s_1_2_2(or_tmp_524, or_tmp_523, fsm_output[6]);
  assign nand_40_nl = ~((fsm_output[7]) & (fsm_output[5]));
  assign mux_tmp_476 = MUX_s_1_2_2(nand_40_nl, or_tmp_524, fsm_output[6]);
  assign or_581_cse = (fsm_output[2]) | (fsm_output[4]);
  assign nand_37_nl = ~((and_273_cse | (fsm_output[4])) & (fsm_output[5]));
  assign mux_491_nl = MUX_s_1_2_2(and_dcpl_44, nand_37_nl, fsm_output[8]);
  assign and_168_nl = or_581_cse & (fsm_output[5]);
  assign mux_490_nl = MUX_s_1_2_2((~ (fsm_output[5])), and_168_nl, fsm_output[8]);
  assign mux_492_nl = MUX_s_1_2_2(mux_491_nl, mux_490_nl, fsm_output[6]);
  assign mux_489_nl = MUX_s_1_2_2((~ (fsm_output[5])), or_610_cse, fsm_output[8]);
  assign nor_143_nl = ~((fsm_output[6]) | mux_489_nl);
  assign mux_493_nl = MUX_s_1_2_2(mux_492_nl, nor_143_nl, fsm_output[7]);
  assign mux_486_nl = MUX_s_1_2_2(and_206_cse, (~ (fsm_output[5])), fsm_output[8]);
  assign nor_144_nl = ~((or_619_cse & (fsm_output[4])) | (fsm_output[5]));
  assign mux_485_nl = MUX_s_1_2_2(nor_144_nl, (fsm_output[5]), fsm_output[8]);
  assign mux_487_nl = MUX_s_1_2_2(mux_486_nl, mux_485_nl, fsm_output[6]);
  assign mux_482_nl = MUX_s_1_2_2((~ (fsm_output[5])), (fsm_output[5]), fsm_output[4]);
  assign mux_483_nl = MUX_s_1_2_2(and_dcpl_13, mux_482_nl, and_273_cse);
  assign mux_484_nl = MUX_s_1_2_2(mux_483_nl, or_tmp_93, fsm_output[8]);
  assign nor_145_nl = ~((fsm_output[6]) | mux_484_nl);
  assign mux_488_nl = MUX_s_1_2_2(mux_487_nl, nor_145_nl, fsm_output[7]);
  assign not_tmp_310 = MUX_s_1_2_2(mux_493_nl, mux_488_nl, fsm_output[3]);
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_21 & and_dcpl_19;
  assign VEC_LOOP_j_1_12_0_sva_11_0_mx0c1 = and_dcpl_21 & and_dcpl_73;
  assign nor_190_nl = ~((fsm_output[8:7]!=2'b00) | (or_619_cse & (fsm_output[3]))
      | (fsm_output[5:4]!=2'b00));
  assign and_94_nl = (fsm_output[8:7]==2'b11) & ((((fsm_output[2:0]!=3'b000)) & (fsm_output[3]))
      | (fsm_output[5:4]!=2'b00));
  assign modExp_result_sva_mx0c0 = MUX_s_1_2_2(nor_190_nl, and_94_nl, fsm_output[6]);
  assign VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c0
      = and_dcpl_123 & (fsm_output[4]) & (~ (fsm_output[1])) & and_dcpl_130;
  assign VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c1
      = ~(mux_tmp_315 | (~ (fsm_output[1])) | (fsm_output[7]) | (fsm_output[0]));
  assign or_394_nl = (fsm_output[3]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[2])
      | (~ and_206_cse);
  assign mux_316_nl = MUX_s_1_2_2(or_394_nl, mux_tmp_315, fsm_output[0]);
  assign and_102_m1c = (~ mux_316_nl) & and_dcpl_84;
  assign and_123_m1c = and_dcpl_26 & and_dcpl_32 & and_dcpl_11;
  assign and_138_m1c = and_dcpl_45 & and_dcpl_73;
  assign nor_273_nl = ~((~ (fsm_output[7])) | (fsm_output[6]) | (fsm_output[8]) |
      (fsm_output[2]));
  assign nor_274_nl = ~((fsm_output[7]) | (~((fsm_output[6]) & (fsm_output[8]) &
      (fsm_output[2]))));
  assign mux_98_nl = MUX_s_1_2_2(nor_273_nl, nor_274_nl, fsm_output[3]);
  assign and_49_nl = mux_98_nl & and_dcpl_13 & and_dcpl_37;
  assign nor_270_nl = ~((~ (fsm_output[2])) | (fsm_output[5]) | (fsm_output[4]) |
      (~ (fsm_output[8])));
  assign nor_271_nl = ~((fsm_output[2]) | (~ (fsm_output[5])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_100_nl = MUX_s_1_2_2(nor_270_nl, nor_271_nl, fsm_output[3]);
  assign and_253_nl = (fsm_output[1]) & (fsm_output[7]) & (fsm_output[6]) & mux_100_nl;
  assign or_124_nl = (~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[2]) | (~
      (fsm_output[5])) | (fsm_output[4]) | (~ (fsm_output[8]));
  assign or_122_nl = (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[2])) | (fsm_output[5])
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_99_nl = MUX_s_1_2_2(or_124_nl, or_122_nl, fsm_output[7]);
  assign nor_272_nl = ~((fsm_output[1]) | mux_99_nl);
  assign mux_101_nl = MUX_s_1_2_2(and_253_nl, nor_272_nl, fsm_output[0]);
  assign nor_268_nl = ~((~ (fsm_output[8])) | (fsm_output[2]) | (~ and_206_cse));
  assign nor_269_nl = ~((fsm_output[8]) | (~ (fsm_output[2])) | (fsm_output[4]) |
      (~ (fsm_output[5])));
  assign mux_102_nl = MUX_s_1_2_2(nor_268_nl, nor_269_nl, fsm_output[6]);
  assign nand_6_nl = ~((fsm_output[7]) & mux_102_nl);
  assign mux_104_nl = MUX_s_1_2_2(mux_tmp_103, nand_6_nl, fsm_output[0]);
  assign and_51_nl = (~ mux_104_nl) & and_dcpl_40;
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_10_5_2((z_out_2[10:1]), (z_out_1[12:3]),
      (COMP_LOOP_acc_psp_1_sva[10:1]), (COMP_LOOP_acc_10_cse_12_1_1_sva[11:2]), (COMP_LOOP_acc_1_cse_2_sva[11:2]),
      {COMP_LOOP_or_cse , COMP_LOOP_or_1_cse , and_49_nl , mux_101_nl , and_51_nl});
  assign vec_rsc_0_0_i_da_d_pff = COMP_LOOP_mux1h_1_itm_mx1;
  assign nor_263_nl = ~((~ (fsm_output[5])) | (fsm_output[4]) | (fsm_output[2]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00) | not_tmp_92);
  assign nor_264_nl = ~((fsm_output[5]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00) | (fsm_output[8]) | (fsm_output[6]));
  assign mux_109_nl = MUX_s_1_2_2(nor_263_nl, nor_264_nl, fsm_output[7]);
  assign and_252_nl = (fsm_output[0]) & mux_109_nl;
  assign or_150_nl = (COMP_LOOP_acc_psp_1_sva[0]) | (VEC_LOOP_j_1_12_0_sva_11_0[0])
      | (fsm_output[8]) | (fsm_output[6]);
  assign or_149_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00) | not_tmp_92;
  assign mux_107_nl = MUX_s_1_2_2(or_150_nl, or_149_nl, fsm_output[2]);
  assign nor_265_nl = ~((~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[4]) |
      mux_107_nl);
  assign nor_266_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00)
      | mux_106_cse);
  assign mux_108_nl = MUX_s_1_2_2(nor_265_nl, nor_266_nl, fsm_output[0]);
  assign mux_110_nl = MUX_s_1_2_2(and_252_nl, mux_108_nl, fsm_output[1]);
  assign or_140_nl = (fsm_output[5]) | (fsm_output[4]) | (~ (fsm_output[2])) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      | (COMP_LOOP_acc_psp_1_sva[0]) | not_tmp_92;
  assign or_138_nl = (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[2])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_105_nl = MUX_s_1_2_2(or_140_nl, or_138_nl, fsm_output[7]);
  assign nor_267_nl = ~((fsm_output[1:0]!=2'b10) | mux_105_nl);
  assign vec_rsc_0_0_i_wea_d_pff = MUX_s_1_2_2(mux_110_nl, nor_267_nl, fsm_output[3]);
  assign nor_256_nl = ~((fsm_output[6:5]!=2'b01) | (VEC_LOOP_j_1_12_0_sva_11_0[0])
      | (z_out_2[0]) | (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[4])) |
      (fsm_output[8]));
  assign nor_257_nl = ~((fsm_output[6:5]!=2'b11) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      | (z_out_2[0]) | (~ (fsm_output[2])) | (~ (fsm_output[7])) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign mux_118_nl = MUX_s_1_2_2(nor_256_nl, nor_257_nl, fsm_output[3]);
  assign and_250_nl = (fsm_output[0]) & mux_118_nl;
  assign nor_258_nl = ~((z_out_1[2:1]!=2'b00) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[4]) | (~ (fsm_output[8])));
  assign mux_113_nl = MUX_s_1_2_2(and_251_cse, nor_258_nl, fsm_output[5]);
  assign mux_114_nl = MUX_s_1_2_2(mux_113_nl, nor_259_cse, fsm_output[6]);
  assign nor_260_nl = ~((fsm_output[6:5]!=2'b01) | (z_out_1[2:1]!=2'b00) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[4]) | (~ (fsm_output[8])));
  assign or_160_nl = (~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00);
  assign mux_115_nl = MUX_s_1_2_2(mux_114_nl, nor_260_nl, or_160_nl);
  assign nor_261_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_1[2:1]!=2'b00) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_116_nl = MUX_s_1_2_2(mux_115_nl, nor_261_nl, fsm_output[3]);
  assign or_157_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[4]) | (~
      (fsm_output[8])) | (z_out_1[2:1]!=2'b00);
  assign or_156_nl = (z_out_1[2:1]!=2'b00) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_112_nl = MUX_s_1_2_2(or_157_nl, or_156_nl, fsm_output[5]);
  assign nor_262_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | mux_112_nl);
  assign mux_117_nl = MUX_s_1_2_2(mux_116_nl, nor_262_nl, fsm_output[0]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(and_250_nl,
      mux_117_nl, fsm_output[1]);
  assign nor_251_nl = ~((~ (fsm_output[5])) | (fsm_output[4]) | (fsm_output[2]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01) | not_tmp_92);
  assign nor_252_nl = ~((fsm_output[5]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01) | (fsm_output[8]) | (fsm_output[6]));
  assign mux_124_nl = MUX_s_1_2_2(nor_251_nl, nor_252_nl, fsm_output[7]);
  assign and_249_nl = (fsm_output[0]) & mux_124_nl;
  assign or_184_nl = (COMP_LOOP_acc_psp_1_sva[0]) | (~ (VEC_LOOP_j_1_12_0_sva_11_0[0]))
      | (fsm_output[8]) | (fsm_output[6]);
  assign or_183_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01) | not_tmp_92;
  assign mux_122_nl = MUX_s_1_2_2(or_184_nl, or_183_nl, fsm_output[2]);
  assign nor_253_nl = ~((~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[4]) |
      mux_122_nl);
  assign nor_254_nl = ~((~((fsm_output[7]) & (fsm_output[5]) & (COMP_LOOP_acc_1_cse_2_sva[1:0]==2'b01)))
      | mux_106_cse);
  assign mux_123_nl = MUX_s_1_2_2(nor_253_nl, nor_254_nl, fsm_output[0]);
  assign mux_125_nl = MUX_s_1_2_2(and_249_nl, mux_123_nl, fsm_output[1]);
  assign or_174_nl = (fsm_output[5]) | (fsm_output[4]) | (~ (fsm_output[2])) | (~
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])) | (COMP_LOOP_acc_psp_1_sva[0]) | not_tmp_92;
  assign or_172_nl = (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[2])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_120_nl = MUX_s_1_2_2(or_174_nl, or_172_nl, fsm_output[7]);
  assign nor_255_nl = ~((fsm_output[1:0]!=2'b10) | mux_120_nl);
  assign vec_rsc_0_1_i_wea_d_pff = MUX_s_1_2_2(mux_125_nl, nor_255_nl, fsm_output[3]);
  assign nor_245_nl = ~((fsm_output[6:5]!=2'b01) | (~ (VEC_LOOP_j_1_12_0_sva_11_0[0]))
      | (z_out_2[0]) | (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[4])) |
      (fsm_output[8]));
  assign and_247_nl = (fsm_output[6:5]==2'b11) & (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      & (~ (z_out_2[0])) & (fsm_output[2]) & (fsm_output[7]) & (fsm_output[4]) &
      (~ (fsm_output[8]));
  assign mux_133_nl = MUX_s_1_2_2(nor_245_nl, and_247_nl, fsm_output[3]);
  assign and_246_nl = (fsm_output[0]) & mux_133_nl;
  assign nor_246_nl = ~((z_out_1[2:1]!=2'b01) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[4]) | (~ (fsm_output[8])));
  assign mux_128_nl = MUX_s_1_2_2(and_251_cse, nor_246_nl, fsm_output[5]);
  assign mux_129_nl = MUX_s_1_2_2(mux_128_nl, nor_259_cse, fsm_output[6]);
  assign nor_248_nl = ~((fsm_output[6:5]!=2'b01) | (z_out_1[2:1]!=2'b01) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[4]) | (~ (fsm_output[8])));
  assign or_195_nl = (~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01);
  assign mux_130_nl = MUX_s_1_2_2(mux_129_nl, nor_248_nl, or_195_nl);
  assign nor_249_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_1[2:1]!=2'b01) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_131_nl = MUX_s_1_2_2(mux_130_nl, nor_249_nl, fsm_output[3]);
  assign or_192_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[4]) | (~
      (fsm_output[8])) | (z_out_1[2:1]!=2'b01);
  assign or_190_nl = (z_out_1[2:1]!=2'b01) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_127_nl = MUX_s_1_2_2(or_192_nl, or_190_nl, fsm_output[5]);
  assign nor_250_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | mux_127_nl);
  assign mux_132_nl = MUX_s_1_2_2(mux_131_nl, nor_250_nl, fsm_output[0]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(and_246_nl,
      mux_132_nl, fsm_output[1]);
  assign nor_239_nl = ~((~ (fsm_output[5])) | (fsm_output[4]) | (fsm_output[2]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[0]) | not_tmp_109);
  assign nor_240_nl = ~((fsm_output[5]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b10) | (fsm_output[8]) | (fsm_output[6]));
  assign mux_139_nl = MUX_s_1_2_2(nor_239_nl, nor_240_nl, fsm_output[7]);
  assign and_244_nl = (fsm_output[0]) & mux_139_nl;
  assign or_216_nl = (~ (COMP_LOOP_acc_psp_1_sva[0])) | (VEC_LOOP_j_1_12_0_sva_11_0[0])
      | (fsm_output[8]) | (fsm_output[6]);
  assign or_215_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[0]) | not_tmp_109;
  assign mux_137_nl = MUX_s_1_2_2(or_216_nl, or_215_nl, fsm_output[2]);
  assign nor_241_nl = ~((~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[4]) |
      mux_137_nl);
  assign and_245_nl = (fsm_output[7]) & (fsm_output[5]) & (COMP_LOOP_acc_1_cse_2_sva[1:0]==2'b10)
      & mux_136_cse;
  assign mux_138_nl = MUX_s_1_2_2(nor_241_nl, and_245_nl, fsm_output[0]);
  assign mux_140_nl = MUX_s_1_2_2(and_244_nl, mux_138_nl, fsm_output[1]);
  assign or_209_nl = (fsm_output[5]) | (fsm_output[4]) | (~ (fsm_output[2])) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      | (~((COMP_LOOP_acc_psp_1_sva[0]) & (fsm_output[8]) & (fsm_output[6])));
  assign or_207_nl = (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[2])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b10) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_135_nl = MUX_s_1_2_2(or_209_nl, or_207_nl, fsm_output[7]);
  assign nor_244_nl = ~((fsm_output[1:0]!=2'b10) | mux_135_nl);
  assign vec_rsc_0_2_i_wea_d_pff = MUX_s_1_2_2(mux_140_nl, nor_244_nl, fsm_output[3]);
  assign nor_233_nl = ~((fsm_output[6:5]!=2'b01) | (VEC_LOOP_j_1_12_0_sva_11_0[0])
      | (~ (z_out_2[0])) | (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign and_242_nl = (fsm_output[6:5]==2'b11) & (~ (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]))
      & (z_out_2[0]) & (fsm_output[2]) & (fsm_output[7]) & (fsm_output[4]) & (~ (fsm_output[8]));
  assign mux_148_nl = MUX_s_1_2_2(nor_233_nl, and_242_nl, fsm_output[3]);
  assign and_241_nl = (fsm_output[0]) & mux_148_nl;
  assign nor_234_nl = ~((fsm_output[6:5]!=2'b01) | (z_out_1[2:1]!=2'b10) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[4]) | (~ (fsm_output[8])));
  assign nor_235_nl = ~((z_out_1[2:1]!=2'b10) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[4]) | (~ (fsm_output[8])));
  assign mux_143_nl = MUX_s_1_2_2(and_251_cse, nor_235_nl, fsm_output[5]);
  assign mux_144_nl = MUX_s_1_2_2(mux_143_nl, nor_259_cse, fsm_output[6]);
  assign nor_45_nl = ~((~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10));
  assign mux_145_nl = MUX_s_1_2_2(nor_234_nl, mux_144_nl, nor_45_nl);
  assign nor_237_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_1[2:1]!=2'b10) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_146_nl = MUX_s_1_2_2(mux_145_nl, nor_237_nl, fsm_output[3]);
  assign or_223_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[4]) | (~
      (fsm_output[8])) | (z_out_1[2:1]!=2'b10);
  assign or_222_nl = (z_out_1[2:1]!=2'b10) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_142_nl = MUX_s_1_2_2(or_223_nl, or_222_nl, fsm_output[5]);
  assign nor_238_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | mux_142_nl);
  assign mux_147_nl = MUX_s_1_2_2(mux_146_nl, nor_238_nl, fsm_output[0]);
  assign vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(and_241_nl,
      mux_147_nl, fsm_output[1]);
  assign nor_226_nl = ~((~ (fsm_output[5])) | (fsm_output[4]) | (fsm_output[2]) |
      (~ nor_tmp_48));
  assign nor_227_nl = ~((fsm_output[5]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b11) | (fsm_output[8]) | (fsm_output[6]));
  assign mux_154_nl = MUX_s_1_2_2(nor_226_nl, nor_227_nl, fsm_output[7]);
  assign and_238_nl = (fsm_output[0]) & mux_154_nl;
  assign nor_229_nl = ~((~ (COMP_LOOP_acc_psp_1_sva[0])) | (~ (VEC_LOOP_j_1_12_0_sva_11_0[0]))
      | (fsm_output[8]) | (fsm_output[6]));
  assign mux_152_nl = MUX_s_1_2_2(nor_229_nl, nor_tmp_48, fsm_output[2]);
  assign nor_228_nl = ~((~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[4]) |
      (~ mux_152_nl));
  assign and_239_nl = (fsm_output[7]) & (fsm_output[5]) & (COMP_LOOP_acc_1_cse_2_sva[1:0]==2'b11)
      & mux_136_cse;
  assign mux_153_nl = MUX_s_1_2_2(nor_228_nl, and_239_nl, fsm_output[0]);
  assign mux_155_nl = MUX_s_1_2_2(and_238_nl, mux_153_nl, fsm_output[1]);
  assign or_239_nl = (fsm_output[5:4]!=2'b00) | (~((fsm_output[2]) & (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      & (COMP_LOOP_acc_psp_1_sva[0]) & (fsm_output[8]) & (fsm_output[6])));
  assign nand_90_nl = ~((fsm_output[5]) & (fsm_output[4]) & (~ (fsm_output[2])) &
      (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b11) & (~ (fsm_output[8])) & (fsm_output[6]));
  assign mux_150_nl = MUX_s_1_2_2(or_239_nl, nand_90_nl, fsm_output[7]);
  assign nor_232_nl = ~((fsm_output[1:0]!=2'b10) | mux_150_nl);
  assign vec_rsc_0_3_i_wea_d_pff = MUX_s_1_2_2(mux_155_nl, nor_232_nl, fsm_output[3]);
  assign nor_220_nl = ~((fsm_output[6:5]!=2'b01) | (~ (VEC_LOOP_j_1_12_0_sva_11_0[0]))
      | (~ (z_out_2[0])) | (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[4]))
      | (fsm_output[8]));
  assign and_235_nl = (fsm_output[6:5]==2'b11) & (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      & (z_out_2[0]) & (fsm_output[2]) & (fsm_output[7]) & (fsm_output[4]) & (~ (fsm_output[8]));
  assign mux_163_nl = MUX_s_1_2_2(nor_220_nl, and_235_nl, fsm_output[3]);
  assign and_234_nl = (fsm_output[0]) & mux_163_nl;
  assign nor_221_nl = ~((fsm_output[6:5]!=2'b01) | (z_out_1[2:1]!=2'b11) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[4]) | (~ (fsm_output[8])));
  assign nor_222_nl = ~((z_out_1[2:1]!=2'b11) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[4]) | (~ (fsm_output[8])));
  assign mux_158_nl = MUX_s_1_2_2(and_251_cse, nor_222_nl, fsm_output[5]);
  assign mux_159_nl = MUX_s_1_2_2(mux_158_nl, nor_259_cse, fsm_output[6]);
  assign and_237_nl = VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm
      & (COMP_LOOP_acc_1_cse_2_sva[1:0]==2'b11);
  assign mux_160_nl = MUX_s_1_2_2(nor_221_nl, mux_159_nl, and_237_nl);
  assign nor_224_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_1[2:1]!=2'b11) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[4])) | (fsm_output[8]));
  assign mux_161_nl = MUX_s_1_2_2(mux_160_nl, nor_224_nl, fsm_output[3]);
  assign or_253_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[4]) | (~((fsm_output[8])
      & (z_out_1[2:1]==2'b11)));
  assign nand_64_nl = ~((z_out_1[2:1]==2'b11) & (fsm_output[2]) & (fsm_output[7])
      & (fsm_output[4]) & (~ (fsm_output[8])));
  assign mux_157_nl = MUX_s_1_2_2(or_253_nl, nand_64_nl, fsm_output[5]);
  assign nor_225_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | mux_157_nl);
  assign mux_162_nl = MUX_s_1_2_2(mux_161_nl, nor_225_nl, fsm_output[0]);
  assign vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(and_234_nl,
      mux_162_nl, fsm_output[1]);
  assign and_dcpl_150 = mux_462_cse & (fsm_output[3]) & (fsm_output[7]) & (~ (fsm_output[6]))
      & (fsm_output[1]) & (fsm_output[0]);
  assign or_tmp_550 = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (fsm_output[7])
      | nand_86_cse;
  assign or_642_nl = (~ (fsm_output[5])) | (fsm_output[1]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[0]);
  assign mux_500_nl = MUX_s_1_2_2(or_642_nl, or_tmp_550, fsm_output[4]);
  assign nor_343_nl = ~((~ (fsm_output[8])) | (fsm_output[6]) | mux_500_nl);
  assign or_638_nl = (fsm_output[5]) | (fsm_output[1]) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[0]);
  assign mux_499_nl = MUX_s_1_2_2(or_tmp_550, or_638_nl, fsm_output[4]);
  assign nor_344_nl = ~((fsm_output[8]) | (~ (fsm_output[6])) | mux_499_nl);
  assign not_tmp_321 = MUX_s_1_2_2(nor_343_nl, nor_344_nl, fsm_output[2]);
  assign nor_nl = ~((fsm_output[6]) | (fsm_output[7]) | (fsm_output[3]));
  assign mux_502_nl = MUX_s_1_2_2(nor_nl, and_220_cse, fsm_output[2]);
  assign and_dcpl_155 = mux_502_nl & (fsm_output[4]) & (~ (fsm_output[8])) & (fsm_output[5])
      & (~ (fsm_output[1])) & (fsm_output[0]);
  assign and_dcpl_156 = (~ (fsm_output[2])) & (fsm_output[0]);
  assign and_dcpl_159 = ~((fsm_output[7]) | (fsm_output[5]));
  assign and_dcpl_160 = ~((fsm_output[4]) | (fsm_output[8]));
  assign and_dcpl_163 = and_dcpl_160 & (~ (fsm_output[3])) & and_dcpl_159 & (~ (fsm_output[6]))
      & (~ (fsm_output[1])) & and_dcpl_156;
  assign and_dcpl_164 = ~((fsm_output[2]) | (fsm_output[0]));
  assign and_dcpl_165 = (~ (fsm_output[6])) & (fsm_output[1]);
  assign and_dcpl_169 = and_dcpl_160 & (fsm_output[3]) & and_dcpl_159 & and_dcpl_165
      & and_dcpl_164;
  assign and_dcpl_173 = (fsm_output[4]) & (~ (fsm_output[8])) & (fsm_output[3]);
  assign and_dcpl_175 = and_dcpl_173 & and_dcpl_159 & (fsm_output[6]) & (fsm_output[1])
      & and_dcpl_164;
  assign and_dcpl_179 = and_dcpl_173 & (fsm_output[7]) & (fsm_output[5]);
  assign and_dcpl_180 = and_dcpl_179 & and_dcpl_165 & (fsm_output[2]) & (fsm_output[0]);
  assign and_dcpl_181 = (fsm_output[2]) & (~ (fsm_output[0]));
  assign and_dcpl_184 = (~ (fsm_output[4])) & (fsm_output[8]);
  assign and_dcpl_187 = and_dcpl_184 & (~ (fsm_output[3])) & (~ (fsm_output[7]))
      & (fsm_output[5]) & and_dcpl_165 & and_dcpl_181;
  assign and_dcpl_191 = and_dcpl_184 & (fsm_output[3]) & (fsm_output[7]) & (~ (fsm_output[5]));
  assign and_dcpl_192 = and_dcpl_191 & and_dcpl_165 & and_dcpl_156;
  assign and_dcpl_193 = (fsm_output[6]) & (~ (fsm_output[1]));
  assign and_dcpl_195 = and_dcpl_179 & and_dcpl_193 & and_dcpl_181;
  assign and_dcpl_197 = and_dcpl_191 & and_dcpl_193 & and_dcpl_164;
  assign and_dcpl_199 = and_dcpl_191 & and_dcpl_193 & and_dcpl_156;
  assign nor_tmp_146 = (fsm_output[5]) & (fsm_output[2]);
  assign not_tmp_368 = ~((fsm_output[3]) & (fsm_output[0]) & (fsm_output[7]));
  assign nor_352_nl = ~((fsm_output[8:3]!=6'b010011));
  assign nor_353_nl = ~((fsm_output[8:3]!=6'b101100));
  assign mux_503_nl = MUX_s_1_2_2(nor_352_nl, nor_353_nl, fsm_output[2]);
  assign and_379_ssc = mux_503_nl & nor_161_cse;
  assign and_387_ssc = (fsm_output==9'b111001001);
  assign and_392_ssc = mux_462_cse & (fsm_output[3]) & (fsm_output[7]) & (~ (fsm_output[6]))
      & and_231_cse;
  assign nand_112_nl = ~((fsm_output[6]) & (fsm_output[7]) & (fsm_output[3]));
  assign mux_505_nl = MUX_s_1_2_2(or_303_cse, nand_112_nl, fsm_output[2]);
  assign and_396_ssc = (~(mux_505_nl | (fsm_output[8]))) & (fsm_output[5:4]==2'b11)
      & and_231_cse;
  assign nor_tmp = or_605_cse & (fsm_output[3]);
  assign or_tmp_586 = and_231_cse | (fsm_output[3]);
  assign or_708_nl = (fsm_output[0]) | (~ modExp_exp_1_0_1_sva) | (fsm_output[3])
      | (~ (fsm_output[1]));
  assign nand_127_nl = ~((fsm_output[0]) & (fsm_output[3]) & (fsm_output[1]));
  assign mux_536_nl = MUX_s_1_2_2(or_708_nl, nand_127_nl, fsm_output[5]);
  assign or_tmp_598 = (fsm_output[7]) | mux_536_nl;
  assign or_tmp_600 = (fsm_output[0]) | (~(modExp_exp_1_0_1_sva & (fsm_output[3])
      & (fsm_output[1])));
  assign and_420_nl = (fsm_output[2]) & (fsm_output[4]) & (fsm_output[5]);
  assign nor_388_nl = ~((fsm_output[2]) | (fsm_output[4]) | (fsm_output[5]));
  assign not_tmp_395 = MUX_s_1_2_2(and_420_nl, nor_388_nl, fsm_output[8]);
  assign COMP_LOOP_nor_3_itm = ~(and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199);
  assign COMP_LOOP_or_24_itm = and_dcpl_175 | and_dcpl_180;
  assign COMP_LOOP_or_25_itm = and_dcpl_187 | and_dcpl_192;
  always @(posedge clk) begin
    if ( mux_96_itm ) begin
      p_sva <= p_rsci_idat;
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_15 & and_dcpl_11) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, (z_out_4[3:0]), STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_3_obj_ld_cse <= 1'b0;
      modExp_exp_1_0_1_sva <= 1'b0;
      modExp_exp_1_1_1_sva <= 1'b0;
      modExp_exp_1_7_1_sva <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_3_obj_ld_cse <= and_dcpl_21 & and_266_cse & (fsm_output[3])
          & (fsm_output[0]) & (~ (z_out_1[2]));
      modExp_exp_1_0_1_sva <= (COMP_LOOP_mux1h_11_nl & (~ and_dcpl_124)) | and_dcpl_127;
      modExp_exp_1_1_1_sva <= COMP_LOOP_mux1h_20_nl & (~((~ mux_tmp_315) & and_dcpl_84
          & (fsm_output[0])));
      modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_37_nl & (~(and_dcpl_76 & and_dcpl_42
          & and_dcpl_29));
    end
  end
  always @(posedge clk) begin
    modulo_result_rem_cmp_a <= MUX1HOT_v_64_5_2(z_out_5, operator_64_false_acc_mut_63_0,
        VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_mul_itm, COMP_LOOP_mux1h_1_itm, VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w5,
        {modulo_result_or_nl , (~ mux_206_nl) , (~ mux_221_nl) , (~ mux_245_nl) ,
        not_tmp_156});
    modulo_result_rem_cmp_b <= p_sva;
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_1, ({operator_64_false_acc_mut_64
        , operator_64_false_acc_mut_63_0}), and_dcpl_68);
    operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_68);
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_tmp_95, mux_252_nl, fsm_output[0]) ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_534_nl ) begin
      operator_64_false_acc_mut_64 <= operator_64_false_mux1h_2_rgt[64];
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_548_nl, mux_539_nl, fsm_output[8]) ) begin
      operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_2_rgt[63:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_1_12_0_sva_11_0 <= 12'b000000000000;
    end
    else if ( and_dcpl_72 | VEC_LOOP_j_1_12_0_sva_11_0_mx0c1 ) begin
      VEC_LOOP_j_1_12_0_sva_11_0 <= MUX_v_12_2_2(12'b000000000000, (z_out_1[11:0]),
          VEC_LOOP_j_1_12_0_sva_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_k_9_1_1_sva_7_0 <= 8'b00000000;
    end
    else if ( MUX_s_1_2_2(mux_552_nl, and_419_nl, fsm_output[6]) ) begin
      COMP_LOOP_k_9_1_1_sva_7_0 <= MUX_v_8_2_2(8'b00000000, (z_out_4[7:0]), or_nl);
    end
  end
  always @(posedge clk) begin
    if ( (modExp_while_and_3 | modExp_while_and_5 | modExp_result_sva_mx0c0 | (~
        mux_314_nl)) & (modExp_result_sva_mx0c0 | modExp_result_and_rgt | modExp_result_and_1_rgt)
        ) begin
      modExp_result_sva <= MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w11, {modExp_result_sva_mx0c0
          , modExp_result_and_rgt , modExp_result_and_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_363_nl, mux_346_nl, fsm_output[8]) ) begin
      COMP_LOOP_mux1h_1_itm <= MUX1HOT_v_64_10_2(r_sva, modulo_result_rem_cmp_z,
          modulo_qr_sva_1_mx0w11, modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
          vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, z_out_5, VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w5,
          {and_100_nl , r_or_nl , r_or_1_nl , and_dcpl_86 , and_105_nl , and_107_nl
          , and_109_nl , and_111_nl , nor_301_nl , not_tmp_156});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_2_lpi_4_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( MUX_s_1_2_2(mux_379_nl, mux_372_nl, fsm_output[8]) ) begin
      tmp_2_lpi_4_dfm <= MUX1HOT_v_64_5_2(({1'b0 , operator_64_false_slc_modExp_exp_63_1_3}),
          vec_rsc_0_0_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_3_i_qa_d,
          {and_dcpl_72 , COMP_LOOP_or_3_nl , COMP_LOOP_or_4_nl , COMP_LOOP_or_5_nl
          , COMP_LOOP_or_6_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva <= 1'b0;
    end
    else if ( and_dcpl_62 | and_dcpl_132 | and_dcpl_77 ) begin
      exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva <= MUX1HOT_s_1_3_2((~ (z_out_1[63])),
          (~ (z_out_4[8])), (~ (readslicef_10_1_9(VEC_LOOP_1_COMP_LOOP_1_acc_11_nl))),
          {and_dcpl_62 , and_dcpl_132 , and_dcpl_77});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_330_nl, nor_331_nl, fsm_output[2]) ) begin
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_mul_itm <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_psp_1_sva <= 11'b00000000000;
    end
    else if ( COMP_LOOP_or_cse ) begin
      COMP_LOOP_acc_psp_1_sva <= z_out_2;
    end
  end
  always @(posedge clk) begin
    if ( VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c0
        | VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c1
        | and_dcpl_64 ) begin
      VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm
          <= MUX1HOT_s_1_3_2((z_out_1[9]), (z_out[9]), (z_out_4[8]), {VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c0
          , VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c1
          , and_dcpl_64});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_449_nl, mux_446_nl, fsm_output[6]) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= nl_COMP_LOOP_acc_1_cse_2_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_0_1_sva_1 <= 1'b0;
    end
    else if ( ~ mux_460_nl ) begin
      modExp_exp_1_0_1_sva_1 <= MUX_s_1_2_2((COMP_LOOP_k_9_1_1_sva_7_0[0]), modExp_exp_1_1_1_sva,
          mux_463_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_2_1_sva <= 1'b0;
    end
    else if ( ~ not_tmp_310 ) begin
      modExp_exp_1_2_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[1]), modExp_exp_1_3_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[2]), {and_dcpl_124 , and_dcpl_139 , and_dcpl_127});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_3_1_sva <= 1'b0;
    end
    else if ( ~ not_tmp_310 ) begin
      modExp_exp_1_3_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[2]), modExp_exp_1_4_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[3]), {and_dcpl_124 , and_dcpl_139 , and_dcpl_127});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_4_1_sva <= 1'b0;
    end
    else if ( ~ not_tmp_310 ) begin
      modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[3]), modExp_exp_1_5_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[4]), {and_dcpl_124 , and_dcpl_139 , and_dcpl_127});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_5_1_sva <= 1'b0;
    end
    else if ( ~ not_tmp_310 ) begin
      modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[4]), modExp_exp_1_6_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[5]), {and_dcpl_124 , and_dcpl_139 , and_dcpl_127});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_6_1_sva <= 1'b0;
    end
    else if ( ~ not_tmp_310 ) begin
      modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[5]), modExp_exp_1_7_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[6]), {and_dcpl_124 , and_dcpl_139 , and_dcpl_127});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= 12'b000000000000;
    end
    else if ( COMP_LOOP_or_1_cse ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_1[12:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_VEC_LOOP_1_acc_1_psp_ftd_1 <= 12'b000000000000;
    end
    else if ( ~((~ and_dcpl_44) | (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[6]))
        | (~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[0])) ) begin
      reg_VEC_LOOP_1_acc_1_psp_ftd_1 <= z_out_1[11:0];
    end
  end
  assign nand_89_nl = ~((fsm_output[2]) & (fsm_output[6]) & (~ (fsm_output[8])) &
      (fsm_output[4]));
  assign or_294_nl = (fsm_output[2]) | (fsm_output[6]) | (~ (fsm_output[8])) | (fsm_output[4]);
  assign mux_225_nl = MUX_s_1_2_2(nand_89_nl, or_294_nl, fsm_output[5]);
  assign nor_212_nl = ~((~ (fsm_output[3])) | (fsm_output[7]) | (fsm_output[1]) |
      mux_225_nl);
  assign nor_213_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[5])) | (fsm_output[2])
      | (fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[4])));
  assign nor_214_nl = ~((fsm_output[1]) | (fsm_output[5]) | (fsm_output[2]) | (~
      (fsm_output[6])) | (fsm_output[8]) | (fsm_output[4]));
  assign mux_223_nl = MUX_s_1_2_2(nor_213_nl, nor_214_nl, fsm_output[7]);
  assign nor_215_nl = ~((fsm_output[5]) | (~ (fsm_output[2])) | (fsm_output[6]) |
      (~ (fsm_output[8])) | (fsm_output[4]));
  assign and_284_nl = (fsm_output[5]) & (fsm_output[2]) & (fsm_output[6]) & (~ (fsm_output[8]))
      & (fsm_output[4]);
  assign mux_222_nl = MUX_s_1_2_2(nor_215_nl, and_284_nl, fsm_output[1]);
  assign and_228_nl = (fsm_output[7]) & mux_222_nl;
  assign mux_224_nl = MUX_s_1_2_2(mux_223_nl, and_228_nl, fsm_output[3]);
  assign mux_226_nl = MUX_s_1_2_2(nor_212_nl, mux_224_nl, fsm_output[0]);
  assign modulo_result_or_nl = and_dcpl_62 | mux_226_nl | and_dcpl_64;
  assign mux_201_nl = MUX_s_1_2_2(nor_tmp_51, or_tmp_242, fsm_output[7]);
  assign mux_202_nl = MUX_s_1_2_2(or_tmp_251, (~ mux_201_nl), fsm_output[4]);
  assign mux_203_nl = MUX_s_1_2_2(mux_202_nl, and_tmp_10, fsm_output[5]);
  assign mux_197_nl = MUX_s_1_2_2(or_tmp_249, or_tmp_247, fsm_output[7]);
  assign mux_198_nl = MUX_s_1_2_2(mux_197_nl, mux_tmp_195, fsm_output[4]);
  assign mux_196_nl = MUX_s_1_2_2(or_tmp_244, mux_tmp_195, fsm_output[4]);
  assign mux_199_nl = MUX_s_1_2_2(mux_198_nl, mux_196_nl, fsm_output[0]);
  assign mux_200_nl = MUX_s_1_2_2(mux_tmp_179, mux_199_nl, fsm_output[5]);
  assign mux_204_nl = MUX_s_1_2_2((~ mux_203_nl), mux_200_nl, fsm_output[6]);
  assign mux_192_nl = MUX_s_1_2_2(mux_tmp_184, mux_tmp_175, fsm_output[0]);
  assign mux_191_nl = MUX_s_1_2_2(or_tmp_244, (~ or_tmp_245), fsm_output[4]);
  assign mux_193_nl = MUX_s_1_2_2(mux_192_nl, mux_191_nl, fsm_output[5]);
  assign mux_194_nl = MUX_s_1_2_2(mux_193_nl, mux_tmp_180, fsm_output[6]);
  assign mux_205_nl = MUX_s_1_2_2(mux_204_nl, mux_194_nl, fsm_output[2]);
  assign mux_185_nl = MUX_s_1_2_2((~ (fsm_output[8])), nor_tmp_51, fsm_output[7]);
  assign mux_186_nl = MUX_s_1_2_2(mux_185_nl, or_tmp_251, fsm_output[4]);
  assign mux_187_nl = MUX_s_1_2_2(mux_186_nl, mux_tmp_184, fsm_output[0]);
  assign nor_219_nl = ~((fsm_output[7]) | (~ or_tmp_247));
  assign mux_181_nl = MUX_s_1_2_2(or_tmp_244, nor_219_nl, fsm_output[4]);
  assign mux_183_nl = MUX_s_1_2_2((~ and_tmp_10), mux_181_nl, fsm_output[0]);
  assign mux_188_nl = MUX_s_1_2_2(mux_187_nl, mux_183_nl, fsm_output[5]);
  assign mux_189_nl = MUX_s_1_2_2(mux_188_nl, mux_tmp_180, fsm_output[6]);
  assign mux_172_nl = MUX_s_1_2_2((fsm_output[8]), (~ or_tmp_247), fsm_output[7]);
  assign mux_173_nl = MUX_s_1_2_2(or_tmp_244, mux_172_nl, fsm_output[4]);
  assign mux_176_nl = MUX_s_1_2_2(mux_tmp_175, mux_173_nl, fsm_output[5]);
  assign or_269_nl = (fsm_output[7]) | (~ nor_tmp_51);
  assign mux_170_nl = MUX_s_1_2_2(or_269_nl, or_tmp_245, fsm_output[4]);
  assign or_266_nl = (fsm_output[8:7]!=2'b01);
  assign mux_165_nl = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_242, fsm_output[7]);
  assign mux_166_nl = MUX_s_1_2_2(or_266_nl, mux_165_nl, fsm_output[4]);
  assign mux_169_nl = MUX_s_1_2_2(mux_tmp_168, mux_166_nl, fsm_output[0]);
  assign mux_171_nl = MUX_s_1_2_2(mux_170_nl, mux_169_nl, fsm_output[5]);
  assign mux_177_nl = MUX_s_1_2_2(mux_176_nl, mux_171_nl, fsm_output[6]);
  assign mux_190_nl = MUX_s_1_2_2(mux_189_nl, mux_177_nl, fsm_output[2]);
  assign mux_206_nl = MUX_s_1_2_2(mux_205_nl, mux_190_nl, fsm_output[1]);
  assign or_286_nl = (fsm_output[8]) | (~ (fsm_output[1])) | (~ (fsm_output[2]))
      | (~ (fsm_output[6])) | (fsm_output[7]);
  assign and_229_nl = or_605_cse & (fsm_output[2]);
  assign mux_217_nl = MUX_s_1_2_2(or_298_cse, or_tmp_255, and_229_nl);
  assign mux_218_nl = MUX_s_1_2_2((fsm_output[6]), mux_217_nl, fsm_output[8]);
  assign mux_219_nl = MUX_s_1_2_2(or_286_nl, mux_218_nl, fsm_output[5]);
  assign or_284_nl = nor_217_cse | (fsm_output[7:6]!=2'b00);
  assign mux_215_nl = MUX_s_1_2_2(or_tmp_255, or_284_nl, fsm_output[8]);
  assign nand_17_nl = ~((fsm_output[8]) & (~(and_230_cse | (fsm_output[7:6]!=2'b01))));
  assign mux_216_nl = MUX_s_1_2_2(mux_215_nl, nand_17_nl, fsm_output[5]);
  assign mux_220_nl = MUX_s_1_2_2(mux_219_nl, mux_216_nl, fsm_output[4]);
  assign or_281_nl = (fsm_output[8:6]!=3'b001);
  assign mux_211_nl = MUX_s_1_2_2((fsm_output[6]), or_298_cse, or_280_cse);
  assign mux_212_nl = MUX_s_1_2_2(mux_211_nl, or_tmp_255, fsm_output[8]);
  assign mux_213_nl = MUX_s_1_2_2(or_281_nl, mux_212_nl, fsm_output[5]);
  assign mux_208_nl = MUX_s_1_2_2(or_tmp_255, or_tmp_254, fsm_output[2]);
  assign mux_207_nl = MUX_s_1_2_2(or_tmp_254, (fsm_output[6]), fsm_output[2]);
  assign mux_209_nl = MUX_s_1_2_2(mux_208_nl, mux_207_nl, or_605_cse);
  assign mux_210_nl = MUX_s_1_2_2(mux_209_nl, or_298_cse, fsm_output[8]);
  assign or_279_nl = (fsm_output[5]) | mux_210_nl;
  assign mux_214_nl = MUX_s_1_2_2(mux_213_nl, or_279_nl, fsm_output[4]);
  assign mux_221_nl = MUX_s_1_2_2(mux_220_nl, mux_214_nl, fsm_output[3]);
  assign or_314_nl = (fsm_output[4]) | (fsm_output[1]) | (fsm_output[3]);
  assign mux_242_nl = MUX_s_1_2_2(or_tmp_254, (~ and_266_cse), or_314_nl);
  assign nand_99_nl = ~((~(or_603_cse & (fsm_output[7]))) & (fsm_output[6]));
  assign mux_243_nl = MUX_s_1_2_2(mux_242_nl, nand_99_nl, fsm_output[5]);
  assign and_221_nl = or_604_cse & (fsm_output[6]);
  assign mux_239_nl = MUX_s_1_2_2(and_220_cse, and_221_nl, or_605_cse);
  assign mux_240_nl = MUX_s_1_2_2(and_266_cse, mux_239_nl, fsm_output[4]);
  assign nand_101_nl = ~((~((fsm_output[3]) & (fsm_output[7]))) & (fsm_output[6]));
  assign or_308_nl = (fsm_output[3]) | (fsm_output[7]) | (~ (fsm_output[6]));
  assign mux_237_nl = MUX_s_1_2_2(nand_101_nl, or_308_nl, and_231_cse);
  assign mux_238_nl = MUX_s_1_2_2(mux_237_nl, or_tmp_255, fsm_output[4]);
  assign mux_241_nl = MUX_s_1_2_2((~ mux_240_nl), mux_238_nl, fsm_output[5]);
  assign mux_244_nl = MUX_s_1_2_2(mux_243_nl, mux_241_nl, fsm_output[2]);
  assign mux_234_nl = MUX_s_1_2_2(or_tmp_255, or_tmp_254, fsm_output[4]);
  assign or_306_nl = (~ (fsm_output[3])) | (~ (fsm_output[7])) | (fsm_output[6]);
  assign mux_232_nl = MUX_s_1_2_2(or_306_nl, or_tmp_277, or_605_cse);
  assign or_304_nl = and_224_cse | (fsm_output[6]);
  assign mux_231_nl = MUX_s_1_2_2(or_304_nl, or_303_cse, and_231_cse);
  assign mux_233_nl = MUX_s_1_2_2(mux_232_nl, mux_231_nl, fsm_output[4]);
  assign mux_235_nl = MUX_s_1_2_2(mux_234_nl, mux_233_nl, fsm_output[5]);
  assign mux_228_nl = MUX_s_1_2_2(or_tmp_255, or_tmp_254, and_226_cse);
  assign mux_229_nl = MUX_s_1_2_2(mux_228_nl, or_tmp_254, fsm_output[4]);
  assign mux_227_nl = MUX_s_1_2_2(or_tmp_277, or_298_cse, fsm_output[4]);
  assign mux_230_nl = MUX_s_1_2_2(mux_229_nl, mux_227_nl, fsm_output[5]);
  assign mux_236_nl = MUX_s_1_2_2(mux_235_nl, mux_230_nl, fsm_output[2]);
  assign mux_245_nl = MUX_s_1_2_2(mux_244_nl, mux_236_nl, fsm_output[8]);
  assign COMP_LOOP_and_11_nl = (~ and_dcpl_82) & and_dcpl_72;
  assign and_288_nl = (~((fsm_output[5]) & (fsm_output[1]) & (fsm_output[2]))) &
      (fsm_output[8]);
  assign or_592_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[2]) | (~
      (fsm_output[8]));
  assign nor_165_nl = ~((~(and_231_cse | (fsm_output[2]))) | (fsm_output[8]));
  assign mux_397_nl = MUX_s_1_2_2(or_592_nl, nor_165_nl, fsm_output[5]);
  assign mux_398_nl = MUX_s_1_2_2(and_288_nl, mux_397_nl, fsm_output[4]);
  assign nor_167_nl = ~((~((fsm_output[2:0]!=3'b110))) | (fsm_output[8]));
  assign and_186_nl = (fsm_output[2]) & (fsm_output[8]);
  assign mux_395_nl = MUX_s_1_2_2(nor_167_nl, and_186_nl, fsm_output[5]);
  assign mux_396_nl = MUX_s_1_2_2(mux_395_nl, mux_tmp_387, fsm_output[4]);
  assign mux_399_nl = MUX_s_1_2_2(mux_398_nl, mux_396_nl, fsm_output[6]);
  assign or_463_nl = (fsm_output[5]) | not_tmp_252;
  assign nor_168_nl = ~(nor_161_cse | (~ (fsm_output[2])) | (fsm_output[8]));
  assign mux_392_nl = MUX_s_1_2_2(nor_168_nl, (fsm_output[8]), fsm_output[5]);
  assign mux_393_nl = MUX_s_1_2_2(or_463_nl, mux_392_nl, fsm_output[4]);
  assign mux_390_nl = MUX_s_1_2_2(not_tmp_252, (fsm_output[8]), fsm_output[5]);
  assign mux_391_nl = MUX_s_1_2_2(mux_tmp_387, mux_390_nl, fsm_output[4]);
  assign mux_394_nl = MUX_s_1_2_2((~ mux_393_nl), mux_391_nl, fsm_output[6]);
  assign mux_400_nl = MUX_s_1_2_2(mux_399_nl, mux_394_nl, fsm_output[3]);
  assign or_458_nl = (~ (fsm_output[5])) | (fsm_output[8]);
  assign mux_388_nl = MUX_s_1_2_2(mux_tmp_387, or_458_nl, fsm_output[4]);
  assign or_459_nl = (fsm_output[6]) | mux_388_nl;
  assign or_457_nl = (fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[8]));
  assign mux_384_nl = MUX_s_1_2_2(or_457_nl, (fsm_output[8]), fsm_output[5]);
  assign or_455_nl = and_187_cse | (fsm_output[8]);
  assign mux_385_nl = MUX_s_1_2_2(mux_384_nl, or_455_nl, fsm_output[4]);
  assign nand_49_nl = ~((fsm_output[4]) & (fsm_output[5]) & (fsm_output[0]) & (fsm_output[1])
      & (fsm_output[2]) & (~ (fsm_output[8])));
  assign mux_386_nl = MUX_s_1_2_2(mux_385_nl, nand_49_nl, fsm_output[6]);
  assign mux_389_nl = MUX_s_1_2_2(or_459_nl, mux_386_nl, fsm_output[3]);
  assign mux_401_nl = MUX_s_1_2_2(mux_400_nl, (~ mux_389_nl), fsm_output[7]);
  assign COMP_LOOP_mux1h_11_nl = MUX1HOT_s_1_4_2((operator_66_true_div_cmp_z[0]),
      (tmp_2_lpi_4_dfm[0]), modExp_exp_1_0_1_sva_1, modExp_exp_1_0_1_sva, {COMP_LOOP_and_11_nl
      , and_dcpl_82 , and_dcpl_125 , mux_401_nl});
  assign nand_38_nl = ~(((fsm_output[7]) | (fsm_output[2])) & (fsm_output[5]));
  assign mux_478_nl = MUX_s_1_2_2(nand_38_nl, or_tmp_524, fsm_output[6]);
  assign mux_479_nl = MUX_s_1_2_2(mux_tmp_476, mux_478_nl, fsm_output[4]);
  assign mux_474_nl = MUX_s_1_2_2((~ (fsm_output[5])), and_187_cse, fsm_output[7]);
  assign or_558_nl = (fsm_output[7]) | (fsm_output[2]) | (fsm_output[0]) | (fsm_output[1])
      | (fsm_output[5]);
  assign mux_475_nl = MUX_s_1_2_2(mux_474_nl, or_558_nl, fsm_output[6]);
  assign mux_477_nl = MUX_s_1_2_2(mux_tmp_476, mux_475_nl, fsm_output[4]);
  assign mux_480_nl = MUX_s_1_2_2(mux_479_nl, mux_477_nl, fsm_output[3]);
  assign and_162_nl = (fsm_output[2]) & or_605_cse & (fsm_output[5]);
  assign mux_470_nl = MUX_s_1_2_2(and_162_nl, (fsm_output[5]), fsm_output[7]);
  assign or_556_nl = (fsm_output[7]) | (~((fsm_output[2]) & (fsm_output[5])));
  assign mux_471_nl = MUX_s_1_2_2(mux_470_nl, or_556_nl, fsm_output[6]);
  assign mux_472_nl = MUX_s_1_2_2(mux_471_nl, mux_tmp_466, fsm_output[4]);
  assign or_555_nl = (fsm_output[2]) | (fsm_output[1]) | (fsm_output[5]);
  assign mux_467_nl = MUX_s_1_2_2((fsm_output[5]), or_555_nl, fsm_output[7]);
  assign mux_468_nl = MUX_s_1_2_2(mux_467_nl, or_tmp_523, fsm_output[6]);
  assign mux_469_nl = MUX_s_1_2_2(mux_468_nl, mux_tmp_466, fsm_output[4]);
  assign mux_473_nl = MUX_s_1_2_2(mux_472_nl, mux_469_nl, fsm_output[3]);
  assign mux_481_nl = MUX_s_1_2_2(mux_480_nl, mux_473_nl, fsm_output[8]);
  assign COMP_LOOP_mux1h_20_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_1_1_sva_7_0[7]),
      modExp_exp_1_2_1_sva, modExp_exp_1_1_1_sva, (COMP_LOOP_k_9_1_1_sva_7_0[1]),
      {and_dcpl_124 , and_dcpl_139 , (~ mux_481_nl) , and_dcpl_127});
  assign COMP_LOOP_mux1h_37_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_1_1_sva_7_0[6]),
      modExp_exp_1_1_1_sva, modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_1_1_sva_7_0[7]),
      {and_dcpl_124 , and_dcpl_132 , not_tmp_310 , and_dcpl_127});
  assign mux_252_nl = MUX_s_1_2_2(mux_tmp_94, and_215_cse, fsm_output[3]);
  assign or_684_nl = (~ (fsm_output[1])) | (fsm_output[3]);
  assign mux_529_nl = MUX_s_1_2_2(and_226_cse, or_684_nl, fsm_output[0]);
  assign mux_530_nl = MUX_s_1_2_2(mux_529_nl, (fsm_output[3]), fsm_output[2]);
  assign nor_394_nl = ~((fsm_output[6]) | mux_530_nl);
  assign and_425_nl = (fsm_output[3:2]==2'b11);
  assign mux_531_nl = MUX_s_1_2_2(nor_394_nl, and_425_nl, fsm_output[4]);
  assign nand_128_nl = ~((fsm_output[6]) & (fsm_output[2]) & (fsm_output[0]) & (fsm_output[1])
      & (fsm_output[3]));
  assign nor_395_nl = ~((fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[0])) |
      (fsm_output[1]) | (fsm_output[3]));
  assign mux_528_nl = MUX_s_1_2_2(nand_128_nl, nor_395_nl, fsm_output[4]);
  assign mux_532_nl = MUX_s_1_2_2(mux_531_nl, mux_528_nl, fsm_output[5]);
  assign nor_398_nl = ~((fsm_output[2]) | or_tmp_586);
  assign mux_526_nl = MUX_s_1_2_2((fsm_output[3]), nor_398_nl, fsm_output[6]);
  assign and_427_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[3]);
  assign mux_525_nl = MUX_s_1_2_2(and_427_nl, (fsm_output[3]), fsm_output[2]);
  assign nor_399_nl = ~((fsm_output[6]) | mux_525_nl);
  assign mux_527_nl = MUX_s_1_2_2(mux_526_nl, nor_399_nl, fsm_output[4]);
  assign and_426_nl = (fsm_output[5]) & mux_527_nl;
  assign mux_533_nl = MUX_s_1_2_2(mux_532_nl, and_426_nl, fsm_output[8]);
  assign and_428_nl = (fsm_output[6]) & ((fsm_output[3:0]!=4'b0000));
  assign and_429_nl = (fsm_output[2]) & (~ or_tmp_586);
  assign nor_396_nl = ~((fsm_output[3:2]!=2'b00));
  assign mux_521_nl = MUX_s_1_2_2(and_429_nl, nor_396_nl, fsm_output[6]);
  assign mux_522_nl = MUX_s_1_2_2(and_428_nl, mux_521_nl, fsm_output[4]);
  assign nor_397_nl = ~((fsm_output[1]) | (~ (fsm_output[3])));
  assign mux_520_nl = MUX_s_1_2_2(nor_tmp, nor_397_nl, fsm_output[2]);
  assign and_430_nl = (fsm_output[4]) & (fsm_output[6]) & mux_520_nl;
  assign mux_523_nl = MUX_s_1_2_2(mux_522_nl, and_430_nl, fsm_output[5]);
  assign and_431_nl = (fsm_output[2]) & nor_tmp;
  assign mux_nl = MUX_s_1_2_2((fsm_output[3]), or_674_cse, fsm_output[2]);
  assign mux_518_nl = MUX_s_1_2_2(and_431_nl, mux_nl, fsm_output[6]);
  assign or_676_nl = (fsm_output[4]) | mux_518_nl;
  assign mux_519_nl = MUX_s_1_2_2(or_676_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_524_nl = MUX_s_1_2_2(mux_523_nl, mux_519_nl, fsm_output[8]);
  assign mux_534_nl = MUX_s_1_2_2(mux_533_nl, mux_524_nl, fsm_output[7]);
  assign nand_125_nl = ~((fsm_output[3]) & (fsm_output[1]));
  assign mux_545_nl = MUX_s_1_2_2(nand_125_nl, (fsm_output[1]), fsm_output[0]);
  assign nor_389_nl = ~((fsm_output[7]) | (fsm_output[5]) | mux_545_nl);
  assign or_700_nl = (~ modExp_exp_1_0_1_sva) | (fsm_output[3]) | (~ (fsm_output[1]));
  assign mux_543_nl = MUX_s_1_2_2((fsm_output[3]), or_700_nl, fsm_output[0]);
  assign and_421_nl = (fsm_output[5]) & (~ mux_543_nl);
  assign nor_390_nl = ~((fsm_output[5]) | (~ (fsm_output[0])) | (~ modExp_exp_1_0_1_sva)
      | (~ (fsm_output[3])) | (fsm_output[1]));
  assign mux_544_nl = MUX_s_1_2_2(and_421_nl, nor_390_nl, fsm_output[7]);
  assign mux_546_nl = MUX_s_1_2_2(nor_389_nl, mux_544_nl, fsm_output[4]);
  assign or_697_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[1]));
  assign mux_542_nl = MUX_s_1_2_2(or_697_nl, or_tmp_600, fsm_output[5]);
  assign and_422_nl = (fsm_output[4]) & (fsm_output[7]) & (~ mux_542_nl);
  assign mux_547_nl = MUX_s_1_2_2(mux_546_nl, and_422_nl, fsm_output[2]);
  assign and_424_nl = ((~ (fsm_output[0])) | modExp_exp_1_0_1_sva) & (fsm_output[3])
      & (fsm_output[1]);
  assign mux_540_nl = MUX_s_1_2_2((~ or_674_cse), and_424_nl, fsm_output[5]);
  assign and_415_nl = (fsm_output[7]) & mux_540_nl;
  assign mux_541_nl = MUX_s_1_2_2((~ or_tmp_598), and_415_nl, fsm_output[4]);
  assign and_423_nl = (fsm_output[2]) & mux_541_nl;
  assign mux_548_nl = MUX_s_1_2_2(mux_547_nl, and_423_nl, fsm_output[6]);
  assign mux_537_nl = MUX_s_1_2_2(or_tmp_600, or_674_cse, fsm_output[5]);
  assign nand_118_nl = ~((fsm_output[7]) & (~ mux_537_nl));
  assign mux_538_nl = MUX_s_1_2_2(nand_118_nl, or_tmp_598, fsm_output[4]);
  assign nor_391_nl = ~((fsm_output[2]) | mux_538_nl);
  assign nor_392_nl = ~((fsm_output[4]) | (fsm_output[7]) | (~ (fsm_output[5])) |
      (~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[1])));
  assign nor_393_nl = ~((fsm_output[4]) | (fsm_output[7]) | (~ (fsm_output[5])) |
      (~ (fsm_output[0])) | (~ modExp_exp_1_0_1_sva) | (fsm_output[3]) | (fsm_output[1]));
  assign mux_535_nl = MUX_s_1_2_2(nor_392_nl, nor_393_nl, fsm_output[2]);
  assign mux_539_nl = MUX_s_1_2_2(nor_391_nl, mux_535_nl, fsm_output[6]);
  assign nand_25_nl = ~((fsm_output[7:6]==2'b11) & (~ mux_tmp_296));
  assign mux_297_nl = MUX_s_1_2_2(or_tmp_351, nand_25_nl, fsm_output[3]);
  assign or_372_nl = (fsm_output[8:2]!=7'b0000010);
  assign mux_298_nl = MUX_s_1_2_2(mux_297_nl, or_372_nl, fsm_output[0]);
  assign or_nl = mux_298_nl | (fsm_output[1]);
  assign nor_386_nl = ~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[7]) | (fsm_output[8])
      | (fsm_output[2]) | (~((fsm_output[5:4]==2'b11))));
  assign nor_387_nl = ~((fsm_output[7]) | (fsm_output[8]) | (fsm_output[2]) | (fsm_output[4])
      | (fsm_output[5]));
  assign and_418_nl = (fsm_output[7]) & not_tmp_395;
  assign mux_551_nl = MUX_s_1_2_2(nor_387_nl, and_418_nl, fsm_output[1]);
  assign and_417_nl = (fsm_output[0]) & mux_551_nl;
  assign mux_552_nl = MUX_s_1_2_2(nor_386_nl, and_417_nl, fsm_output[3]);
  assign and_419_nl = (~((~ (fsm_output[3])) | (fsm_output[0]) | (fsm_output[1])
      | (~ (fsm_output[7])))) & not_tmp_395;
  assign mux_312_nl = MUX_s_1_2_2(not_tmp_197, and_215_cse, fsm_output[4]);
  assign mux_309_nl = MUX_s_1_2_2(not_tmp_197, and_215_cse, or_581_cse);
  assign mux_307_nl = MUX_s_1_2_2(mux_tmp_40, and_215_cse, fsm_output[4]);
  assign mux_306_nl = MUX_s_1_2_2(and_215_cse, mux_tmp_40, fsm_output[4]);
  assign mux_308_nl = MUX_s_1_2_2(mux_307_nl, mux_306_nl, fsm_output[2]);
  assign mux_310_nl = MUX_s_1_2_2(mux_309_nl, mux_308_nl, fsm_output[0]);
  assign mux_311_nl = MUX_s_1_2_2(mux_310_nl, and_215_cse, fsm_output[1]);
  assign mux_313_nl = MUX_s_1_2_2(mux_312_nl, mux_311_nl, fsm_output[3]);
  assign mux_314_nl = MUX_s_1_2_2(mux_313_nl, and_215_cse, fsm_output[5]);
  assign and_100_nl = and_dcpl_15 & and_dcpl_78;
  assign r_or_nl = ((~ (modulo_result_rem_cmp_z[63])) & and_102_m1c) | (not_tmp_236
      & and_dcpl_97 & (fsm_output[0]) & (~ (modulo_result_rem_cmp_z[63])));
  assign r_or_1_nl = ((modulo_result_rem_cmp_z[63]) & and_102_m1c) | (not_tmp_236
      & and_dcpl_97 & (fsm_output[0]) & (modulo_result_rem_cmp_z[63]));
  assign and_105_nl = not_tmp_208 & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b00);
  assign and_107_nl = not_tmp_208 & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b01);
  assign and_109_nl = not_tmp_208 & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b10);
  assign and_111_nl = not_tmp_208 & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b11);
  assign nor_302_nl = ~((fsm_output[4:2]!=3'b011) | not_tmp_20);
  assign nor_303_nl = ~((fsm_output[2]) | (~ (fsm_output[3])) | (fsm_output[4]) |
      (fsm_output[0]) | (fsm_output[7]));
  assign mux_17_nl = MUX_s_1_2_2(nor_302_nl, nor_303_nl, fsm_output[5]);
  assign nand_nl = ~((fsm_output[8]) & mux_17_nl);
  assign or_32_nl = (fsm_output[4:3]!=2'b00) | not_tmp_20;
  assign or_30_nl = (~ (fsm_output[3])) | (~ (fsm_output[4])) | (fsm_output[0]) |
      (fsm_output[7]);
  assign mux_16_nl = MUX_s_1_2_2(or_32_nl, or_30_nl, fsm_output[2]);
  assign or_620_nl = (fsm_output[8]) | (fsm_output[5]) | mux_16_nl;
  assign mux_18_nl = MUX_s_1_2_2(nand_nl, or_620_nl, fsm_output[6]);
  assign nor_301_nl = ~(mux_18_nl | (fsm_output[1]));
  assign or_593_nl = (fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[7]));
  assign or_594_nl = (fsm_output[0]) | (~ and_224_cse);
  assign mux_359_nl = MUX_s_1_2_2(or_593_nl, or_594_nl, fsm_output[4]);
  assign nand_51_nl = ~((fsm_output[4]) & (fsm_output[7]));
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, nand_51_nl, fsm_output[5]);
  assign mux_358_nl = MUX_s_1_2_2((~ nor_tmp_97), nor_tmp_97, fsm_output[5]);
  assign mux_361_nl = MUX_s_1_2_2(mux_360_nl, mux_358_nl, fsm_output[6]);
  assign nand_52_nl = ~((fsm_output[5]) & nor_tmp_97);
  assign mux_355_nl = MUX_s_1_2_2((fsm_output[7]), mux_tmp_341, fsm_output[4]);
  assign mux_356_nl = MUX_s_1_2_2((~ mux_355_nl), nor_tmp_97, fsm_output[5]);
  assign mux_357_nl = MUX_s_1_2_2(nand_52_nl, mux_356_nl, fsm_output[6]);
  assign mux_362_nl = MUX_s_1_2_2(mux_361_nl, mux_357_nl, fsm_output[2]);
  assign or_595_nl = (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign nand_53_nl = ~((fsm_output[4]) & ((~((~ (fsm_output[0])) | (fsm_output[3])))
      | (fsm_output[7])));
  assign mux_352_nl = MUX_s_1_2_2(or_595_nl, nand_53_nl, fsm_output[5]);
  assign nand_54_nl = ~(((~ (fsm_output[4])) | (~ (fsm_output[0])) | (fsm_output[3]))
      & (fsm_output[7]));
  assign mux_351_nl = MUX_s_1_2_2(nand_54_nl, nor_tmp_97, fsm_output[5]);
  assign mux_353_nl = MUX_s_1_2_2(mux_352_nl, mux_351_nl, fsm_output[6]);
  assign mux_349_nl = MUX_s_1_2_2(and_224_cse, (~ or_tmp_398), fsm_output[4]);
  assign nand_55_nl = ~((fsm_output[5]) & mux_349_nl);
  assign nor_181_nl = ~(((fsm_output[4:3]==2'b11)) | (fsm_output[7]));
  assign mux_347_nl = MUX_s_1_2_2(or_604_cse, (~ or_tmp_398), fsm_output[4]);
  assign mux_348_nl = MUX_s_1_2_2(nor_181_nl, mux_347_nl, fsm_output[5]);
  assign mux_350_nl = MUX_s_1_2_2(nand_55_nl, mux_348_nl, fsm_output[6]);
  assign mux_354_nl = MUX_s_1_2_2(mux_353_nl, mux_350_nl, fsm_output[2]);
  assign mux_363_nl = MUX_s_1_2_2(mux_362_nl, mux_354_nl, fsm_output[1]);
  assign mux_342_nl = MUX_s_1_2_2((~ mux_tmp_341), and_224_cse, fsm_output[4]);
  assign mux_343_nl = MUX_s_1_2_2((~ (fsm_output[7])), mux_342_nl, fsm_output[5]);
  assign mux_344_nl = MUX_s_1_2_2(mux_343_nl, mux_68_cse, fsm_output[6]);
  assign nor_182_nl = ~((fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_338_nl = MUX_s_1_2_2(nor_182_nl, (fsm_output[7]), fsm_output[4]);
  assign mux_339_nl = MUX_s_1_2_2((~ mux_338_nl), mux_63_cse, fsm_output[5]);
  assign or_426_nl = (fsm_output[4]) | and_196_cse | (fsm_output[7]);
  assign or_424_nl = (fsm_output[0]) | (fsm_output[3]) | (fsm_output[7]);
  assign or_104_nl = (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_336_nl = MUX_s_1_2_2(or_424_nl, or_104_nl, fsm_output[4]);
  assign mux_337_nl = MUX_s_1_2_2(or_426_nl, mux_336_nl, fsm_output[5]);
  assign mux_340_nl = MUX_s_1_2_2(mux_339_nl, mux_337_nl, fsm_output[6]);
  assign mux_345_nl = MUX_s_1_2_2(mux_344_nl, mux_340_nl, fsm_output[2]);
  assign mux_332_nl = MUX_s_1_2_2(or_tmp_398, (~ (fsm_output[7])), fsm_output[4]);
  assign mux_331_nl = MUX_s_1_2_2((~ or_604_cse), or_604_cse, fsm_output[4]);
  assign mux_333_nl = MUX_s_1_2_2(mux_332_nl, mux_331_nl, fsm_output[5]);
  assign mux_334_nl = MUX_s_1_2_2(mux_333_nl, mux_68_cse, fsm_output[6]);
  assign nand_87_nl = ~((~((fsm_output[4]) & (fsm_output[0]) & (fsm_output[3])))
      & (fsm_output[7]));
  assign mux_328_nl = MUX_s_1_2_2(nand_87_nl, mux_63_cse, fsm_output[5]);
  assign or_418_nl = (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7]);
  assign mux_326_nl = MUX_s_1_2_2(or_418_nl, or_tmp_69, fsm_output[5]);
  assign mux_329_nl = MUX_s_1_2_2(mux_328_nl, mux_326_nl, fsm_output[6]);
  assign mux_335_nl = MUX_s_1_2_2(mux_334_nl, mux_329_nl, fsm_output[2]);
  assign mux_346_nl = MUX_s_1_2_2(mux_345_nl, mux_335_nl, fsm_output[1]);
  assign COMP_LOOP_or_3_nl = ((~((VEC_LOOP_j_1_12_0_sva_11_0[0]) | (COMP_LOOP_acc_psp_1_sva[0])))
      & and_123_m1c) | ((~ mux_tmp_103) & and_dcpl_105 & (~ (COMP_LOOP_acc_1_cse_2_sva[0]))
      & and_dcpl_23) | ((~((reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) | (COMP_LOOP_acc_psp_1_sva[0])))
      & and_138_m1c);
  assign COMP_LOOP_or_4_nl = ((COMP_LOOP_acc_psp_1_sva[0]) & (~ (VEC_LOOP_j_1_12_0_sva_11_0[0]))
      & and_123_m1c) | ((~ mux_tmp_103) & and_dcpl_112 & (~ (COMP_LOOP_acc_1_cse_2_sva[0]))
      & and_dcpl_23) | ((COMP_LOOP_acc_psp_1_sva[0]) & (~ (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]))
      & and_138_m1c);
  assign COMP_LOOP_or_5_nl = ((VEC_LOOP_j_1_12_0_sva_11_0[0]) & (~ (COMP_LOOP_acc_psp_1_sva[0]))
      & and_123_m1c) | ((~ mux_tmp_103) & and_dcpl_105 & (COMP_LOOP_acc_1_cse_2_sva[0])
      & and_dcpl_23) | ((reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) & (~ (COMP_LOOP_acc_psp_1_sva[0]))
      & and_138_m1c);
  assign COMP_LOOP_or_6_nl = ((VEC_LOOP_j_1_12_0_sva_11_0[0]) & (COMP_LOOP_acc_psp_1_sva[0])
      & and_123_m1c) | ((~ mux_tmp_103) & and_dcpl_112 & (COMP_LOOP_acc_1_cse_2_sva[0])
      & and_dcpl_23) | ((reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) & (COMP_LOOP_acc_psp_1_sva[0])
      & and_138_m1c);
  assign and_189_nl = (fsm_output[2]) & (fsm_output[7]) & (fsm_output[4]);
  assign mux_377_nl = MUX_s_1_2_2(or_tmp_417, and_189_nl, fsm_output[6]);
  assign nor_174_nl = ~((fsm_output[2]) | and_231_cse | (fsm_output[7]) | (~ (fsm_output[4])));
  assign mux_376_nl = MUX_s_1_2_2(nor_174_nl, or_95_cse, fsm_output[6]);
  assign mux_378_nl = MUX_s_1_2_2(mux_377_nl, mux_376_nl, fsm_output[5]);
  assign nor_175_nl = ~((~(nor_217_cse | (fsm_output[7]))) | (fsm_output[4]));
  assign mux_374_nl = MUX_s_1_2_2(nor_175_nl, nor_tmp_103, fsm_output[6]);
  assign mux_373_nl = MUX_s_1_2_2(or_95_cse, (~ nor_tmp_103), and_230_cse);
  assign and_191_nl = (fsm_output[6]) & mux_373_nl;
  assign mux_375_nl = MUX_s_1_2_2(mux_374_nl, and_191_nl, fsm_output[5]);
  assign mux_379_nl = MUX_s_1_2_2(mux_378_nl, mux_375_nl, fsm_output[3]);
  assign or_440_nl = (~ (fsm_output[6])) | (fsm_output[2]);
  assign mux_370_nl = MUX_s_1_2_2(or_tmp_417, (fsm_output[7]), or_440_nl);
  assign mux_371_nl = MUX_s_1_2_2((fsm_output[6]), mux_370_nl, fsm_output[5]);
  assign mux_366_nl = MUX_s_1_2_2((fsm_output[7]), or_95_cse, and_231_cse);
  assign mux_367_nl = MUX_s_1_2_2(mux_366_nl, or_95_cse, fsm_output[2]);
  assign mux_368_nl = MUX_s_1_2_2(mux_367_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_369_nl = MUX_s_1_2_2((fsm_output[6]), mux_368_nl, fsm_output[5]);
  assign mux_372_nl = MUX_s_1_2_2(mux_371_nl, mux_369_nl, fsm_output[3]);
  assign nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl = ({z_out_4 , 1'b0}) + ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))})
      + 10'b0000000001;
  assign VEC_LOOP_1_COMP_LOOP_1_acc_11_nl = nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl[9:0];
  assign or_506_nl = (fsm_output[6]) | (~ (fsm_output[8])) | (fsm_output[0]) | (fsm_output[1])
      | (fsm_output[4]);
  assign or_505_nl = (fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[0])) | (~
      (fsm_output[1])) | (fsm_output[4]);
  assign mux_436_nl = MUX_s_1_2_2(or_506_nl, or_505_nl, fsm_output[3]);
  assign or_504_nl = (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[0])
      | (fsm_output[1]) | (~ (fsm_output[4]));
  assign mux_437_nl = MUX_s_1_2_2(mux_436_nl, or_504_nl, fsm_output[7]);
  assign nor_330_nl = ~((fsm_output[5]) | mux_437_nl);
  assign or_501_nl = (fsm_output[8]) | (fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[4]));
  assign or_499_nl = (~ (fsm_output[8])) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[4]);
  assign mux_435_nl = MUX_s_1_2_2(or_501_nl, or_499_nl, fsm_output[6]);
  assign nor_331_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[3]) |
      mux_435_nl);
  assign COMP_LOOP_mux_88_nl = MUX_v_12_2_2(VEC_LOOP_j_1_12_0_sva_11_0, reg_VEC_LOOP_1_acc_1_psp_ftd_1,
      and_434_cse);
  assign nl_COMP_LOOP_acc_1_cse_2_sva  = COMP_LOOP_mux_88_nl + conv_u2u_9_12({COMP_LOOP_k_9_1_1_sva_7_0
      , 1'b1});
  assign and_175_nl = (fsm_output[0]) & (fsm_output[8]) & (fsm_output[7]);
  assign mux_447_nl = MUX_s_1_2_2(not_tmp_38, and_175_nl, fsm_output[1]);
  assign mux_448_nl = MUX_s_1_2_2(mux_447_nl, and_182_cse, or_621_cse);
  assign mux_449_nl = MUX_s_1_2_2(not_tmp_38, mux_448_nl, and_206_cse);
  assign and_177_nl = (and_230_cse | (fsm_output[8])) & (fsm_output[7]);
  assign mux_444_nl = MUX_s_1_2_2(and_177_nl, (fsm_output[7]), fsm_output[3]);
  assign and_179_nl = (~((fsm_output[3]) & (fsm_output[2]) & (fsm_output[1]) & (~
      (fsm_output[8])))) & (fsm_output[7]);
  assign mux_445_nl = MUX_s_1_2_2(mux_444_nl, and_179_nl, fsm_output[4]);
  assign mux_446_nl = MUX_s_1_2_2(and_182_cse, mux_445_nl, fsm_output[5]);
  assign and_172_nl = (fsm_output[1]) & (fsm_output[7]) & (~ (fsm_output[6])) & (fsm_output[3])
      & mux_462_cse;
  assign or_544_nl = (fsm_output[3]) | (~ (fsm_output[2])) | (~ (fsm_output[5]))
      | (fsm_output[4]) | (~ (fsm_output[8]));
  assign or_542_nl = (~ (fsm_output[3])) | (fsm_output[2]) | (fsm_output[5]) | (~
      (fsm_output[4])) | (fsm_output[8]);
  assign mux_461_nl = MUX_s_1_2_2(or_544_nl, or_542_nl, fsm_output[6]);
  assign nor_148_nl = ~((fsm_output[1]) | (fsm_output[7]) | mux_461_nl);
  assign mux_463_nl = MUX_s_1_2_2(and_172_nl, nor_148_nl, fsm_output[0]);
  assign nor_326_nl = ~((fsm_output[3]) | (fsm_output[2]) | (fsm_output[1]) | (~
      (fsm_output[8])));
  assign mux_457_nl = MUX_s_1_2_2((fsm_output[8]), nor_326_nl, fsm_output[4]);
  assign or_538_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[8]);
  assign mux_456_nl = MUX_s_1_2_2(or_538_nl, (fsm_output[8]), or_621_cse);
  assign and_286_nl = (fsm_output[4]) & (~ mux_456_nl);
  assign mux_458_nl = MUX_s_1_2_2(mux_457_nl, and_286_nl, fsm_output[5]);
  assign nor_327_nl = ~((fsm_output[4:3]!=2'b00) | and_273_cse | (fsm_output[8]));
  assign and_287_nl = ((fsm_output[4:2]!=3'b000)) & (fsm_output[8]);
  assign mux_455_nl = MUX_s_1_2_2(nor_327_nl, and_287_nl, fsm_output[5]);
  assign mux_459_nl = MUX_s_1_2_2(mux_458_nl, mux_455_nl, fsm_output[6]);
  assign nor_316_nl = ~((fsm_output[2]) | (fsm_output[1]) | (~ (fsm_output[8])));
  assign mux_451_nl = MUX_s_1_2_2((fsm_output[8]), nor_316_nl, fsm_output[3]);
  assign nor_317_nl = ~((~ (fsm_output[3])) | (fsm_output[8]));
  assign mux_452_nl = MUX_s_1_2_2(mux_451_nl, nor_317_nl, fsm_output[4]);
  assign nor_318_nl = ~(((fsm_output[4:1]==4'b1111)) | (fsm_output[8]));
  assign mux_453_nl = MUX_s_1_2_2(mux_452_nl, nor_318_nl, fsm_output[5]);
  assign and_283_nl = (fsm_output[5]) & (fsm_output[4]) & (fsm_output[3]) & (fsm_output[2])
      & (fsm_output[0]) & (fsm_output[1]) & (~ (fsm_output[8]));
  assign mux_454_nl = MUX_s_1_2_2(mux_453_nl, and_283_nl, fsm_output[6]);
  assign mux_460_nl = MUX_s_1_2_2(mux_459_nl, mux_454_nl, fsm_output[7]);
  assign COMP_LOOP_mux_85_nl = MUX_v_10_2_2(({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))}),
      STAGE_LOOP_lshift_psp_sva, and_dcpl_150);
  assign nor_400_nl = ~((~ (fsm_output[6])) | (fsm_output[5]) | (~ (fsm_output[4]))
      | (fsm_output[8]) | (~ (fsm_output[3])));
  assign nor_401_nl = ~((fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[4]) |
      (~ (fsm_output[8])) | (fsm_output[3]));
  assign mux_555_nl = MUX_s_1_2_2(nor_400_nl, nor_401_nl, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_nand_1_nl = ~(and_dcpl_150 & (~(mux_555_nl & (~ (fsm_output[7]))
      & (fsm_output[1]) & (~ (fsm_output[0])))));
  assign nl_acc_nl = ({COMP_LOOP_mux_85_nl , COMP_LOOP_COMP_LOOP_nand_1_nl}) + conv_u2u_10_11({COMP_LOOP_k_9_1_1_sva_7_0
      , 2'b11});
  assign acc_nl = nl_acc_nl[10:0];
  assign z_out = readslicef_11_10_1(acc_nl);
  assign COMP_LOOP_mux_86_nl = MUX_s_1_2_2((tmp_2_lpi_4_dfm[63]), (p_sva[63]), and_dcpl_163);
  assign COMP_LOOP_COMP_LOOP_or_53_nl = (COMP_LOOP_mux_86_nl & COMP_LOOP_nor_3_itm)
      | and_dcpl_155 | and_dcpl_169;
  assign COMP_LOOP_mux1h_67_nl = MUX1HOT_v_51_3_2((tmp_2_lpi_4_dfm[62:12]), (p_sva[62:12]),
      (~ (operator_64_false_acc_mut_63_0[62:12])), {not_tmp_321 , and_dcpl_163 ,
      and_dcpl_169});
  assign COMP_LOOP_and_70_nl = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      COMP_LOOP_mux1h_67_nl, COMP_LOOP_nor_3_itm);
  assign COMP_LOOP_or_32_nl = MUX_v_51_2_2(COMP_LOOP_and_70_nl, 51'b111111111111111111111111111111111111111111111111111,
      and_dcpl_155);
  assign COMP_LOOP_mux1h_68_nl = MUX1HOT_v_2_5_2((tmp_2_lpi_4_dfm[11:10]), (p_sva[11:10]),
      (~ (operator_64_false_acc_mut_63_0[11:10])), (VEC_LOOP_j_1_12_0_sva_11_0[11:10]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:10]), {not_tmp_321 , and_dcpl_163 , and_dcpl_169
      , and_dcpl_195 , and_dcpl_197});
  assign COMP_LOOP_nor_59_nl = ~(and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_199);
  assign COMP_LOOP_and_71_nl = MUX_v_2_2_2(2'b00, COMP_LOOP_mux1h_68_nl, COMP_LOOP_nor_59_nl);
  assign COMP_LOOP_or_33_nl = MUX_v_2_2_2(COMP_LOOP_and_71_nl, 2'b11, and_dcpl_155);
  assign nl_COMP_LOOP_acc_33_nl = (STAGE_LOOP_lshift_psp_sva[9:1]) + conv_u2u_8_9(COMP_LOOP_k_9_1_1_sva_7_0);
  assign COMP_LOOP_acc_33_nl = nl_COMP_LOOP_acc_33_nl[8:0];
  assign COMP_LOOP_or_34_nl = and_dcpl_175 | and_dcpl_187;
  assign COMP_LOOP_or_35_nl = and_dcpl_180 | and_dcpl_192;
  assign COMP_LOOP_mux1h_69_nl = MUX1HOT_v_10_9_2((tmp_2_lpi_4_dfm[9:0]), ({1'b1
      , (~ COMP_LOOP_k_9_1_1_sva_7_0) , 1'b1}), (p_sva[9:0]), (~ (operator_64_false_acc_mut_63_0[9:0])),
      ({COMP_LOOP_acc_33_nl , (STAGE_LOOP_lshift_psp_sva[0])}), z_out, (VEC_LOOP_j_1_12_0_sva_11_0[9:0]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[9:0]), ({7'b0000000 , (z_out_4[3:1])}), {not_tmp_321
      , and_dcpl_155 , and_dcpl_163 , and_dcpl_169 , COMP_LOOP_or_34_nl , COMP_LOOP_or_35_nl
      , and_dcpl_195 , and_dcpl_197 , and_dcpl_199});
  assign COMP_LOOP_or_36_nl = (~(and_dcpl_155 | and_dcpl_163 | and_dcpl_169 | and_dcpl_175
      | and_dcpl_180 | and_dcpl_187 | and_dcpl_192 | and_dcpl_195 | and_dcpl_197
      | and_dcpl_199)) | not_tmp_321;
  assign COMP_LOOP_COMP_LOOP_or_54_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[63]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_55_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[62]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_56_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[61]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_57_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[60]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_58_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[59]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_59_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[58]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_60_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[57]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_61_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[56]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_62_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[55]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_63_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[54]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_64_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[53]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_65_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[52]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_66_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[51]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_67_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[50]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_68_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[49]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_69_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[48]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_70_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[47]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_71_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[46]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_72_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[45]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_73_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[44]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_74_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[43]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_75_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[42]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_76_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[41]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_77_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[40]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_78_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[39]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_79_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[38]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_80_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[37]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_81_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[36]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_82_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[35]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_83_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[34]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_84_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[33]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_85_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[32]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_86_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[31]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_87_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[30]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_88_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[29]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_89_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[28]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_90_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[27]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_91_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[26]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_92_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[25]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_93_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[24]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_94_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[23]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_95_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[22]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_96_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[21]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_97_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[20]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_98_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[19]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_99_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[18]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_100_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[17]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_101_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[16]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_102_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[15]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_103_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[14]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_104_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[13]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_COMP_LOOP_or_105_nl = (~((COMP_LOOP_mux1h_1_itm_mx1[12]) | and_dcpl_155
      | and_dcpl_169 | and_dcpl_175 | and_dcpl_180 | and_dcpl_187 | and_dcpl_192
      | and_dcpl_195 | and_dcpl_197 | and_dcpl_199)) | and_dcpl_163;
  assign COMP_LOOP_mux1h_70_nl = MUX1HOT_v_2_3_2((~ (COMP_LOOP_mux1h_1_itm_mx1[11:10])),
      (VEC_LOOP_j_1_12_0_sva_11_0[11:10]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:10]),
      {not_tmp_321 , COMP_LOOP_or_24_itm , COMP_LOOP_or_25_itm});
  assign COMP_LOOP_nor_61_nl = ~(and_dcpl_155 | and_dcpl_169 | and_dcpl_195 | and_dcpl_197
      | and_dcpl_199);
  assign COMP_LOOP_and_72_nl = MUX_v_2_2_2(2'b00, COMP_LOOP_mux1h_70_nl, COMP_LOOP_nor_61_nl);
  assign COMP_LOOP_or_37_nl = MUX_v_2_2_2(COMP_LOOP_and_72_nl, 2'b11, and_dcpl_163);
  assign COMP_LOOP_or_39_nl = and_dcpl_155 | and_dcpl_169;
  assign COMP_LOOP_or_40_nl = and_dcpl_195 | and_dcpl_197;
  assign COMP_LOOP_mux1h_71_nl = MUX1HOT_v_10_6_2((~ (COMP_LOOP_mux1h_1_itm_mx1[9:0])),
      10'b0000000001, (VEC_LOOP_j_1_12_0_sva_11_0[9:0]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[9:0]),
      STAGE_LOOP_lshift_psp_sva, 10'b0000000011, {not_tmp_321 , COMP_LOOP_or_39_nl
      , COMP_LOOP_or_24_itm , COMP_LOOP_or_25_itm , COMP_LOOP_or_40_nl , and_dcpl_199});
  assign COMP_LOOP_or_38_nl = MUX_v_10_2_2(COMP_LOOP_mux1h_71_nl, 10'b1111111111,
      and_dcpl_163);
  assign nl_acc_1_nl = conv_u2u_65_66({COMP_LOOP_COMP_LOOP_or_53_nl , COMP_LOOP_or_32_nl
      , COMP_LOOP_or_33_nl , COMP_LOOP_mux1h_69_nl , COMP_LOOP_or_36_nl}) + conv_s2u_65_66({COMP_LOOP_COMP_LOOP_or_54_nl
      , COMP_LOOP_COMP_LOOP_or_55_nl , COMP_LOOP_COMP_LOOP_or_56_nl , COMP_LOOP_COMP_LOOP_or_57_nl
      , COMP_LOOP_COMP_LOOP_or_58_nl , COMP_LOOP_COMP_LOOP_or_59_nl , COMP_LOOP_COMP_LOOP_or_60_nl
      , COMP_LOOP_COMP_LOOP_or_61_nl , COMP_LOOP_COMP_LOOP_or_62_nl , COMP_LOOP_COMP_LOOP_or_63_nl
      , COMP_LOOP_COMP_LOOP_or_64_nl , COMP_LOOP_COMP_LOOP_or_65_nl , COMP_LOOP_COMP_LOOP_or_66_nl
      , COMP_LOOP_COMP_LOOP_or_67_nl , COMP_LOOP_COMP_LOOP_or_68_nl , COMP_LOOP_COMP_LOOP_or_69_nl
      , COMP_LOOP_COMP_LOOP_or_70_nl , COMP_LOOP_COMP_LOOP_or_71_nl , COMP_LOOP_COMP_LOOP_or_72_nl
      , COMP_LOOP_COMP_LOOP_or_73_nl , COMP_LOOP_COMP_LOOP_or_74_nl , COMP_LOOP_COMP_LOOP_or_75_nl
      , COMP_LOOP_COMP_LOOP_or_76_nl , COMP_LOOP_COMP_LOOP_or_77_nl , COMP_LOOP_COMP_LOOP_or_78_nl
      , COMP_LOOP_COMP_LOOP_or_79_nl , COMP_LOOP_COMP_LOOP_or_80_nl , COMP_LOOP_COMP_LOOP_or_81_nl
      , COMP_LOOP_COMP_LOOP_or_82_nl , COMP_LOOP_COMP_LOOP_or_83_nl , COMP_LOOP_COMP_LOOP_or_84_nl
      , COMP_LOOP_COMP_LOOP_or_85_nl , COMP_LOOP_COMP_LOOP_or_86_nl , COMP_LOOP_COMP_LOOP_or_87_nl
      , COMP_LOOP_COMP_LOOP_or_88_nl , COMP_LOOP_COMP_LOOP_or_89_nl , COMP_LOOP_COMP_LOOP_or_90_nl
      , COMP_LOOP_COMP_LOOP_or_91_nl , COMP_LOOP_COMP_LOOP_or_92_nl , COMP_LOOP_COMP_LOOP_or_93_nl
      , COMP_LOOP_COMP_LOOP_or_94_nl , COMP_LOOP_COMP_LOOP_or_95_nl , COMP_LOOP_COMP_LOOP_or_96_nl
      , COMP_LOOP_COMP_LOOP_or_97_nl , COMP_LOOP_COMP_LOOP_or_98_nl , COMP_LOOP_COMP_LOOP_or_99_nl
      , COMP_LOOP_COMP_LOOP_or_100_nl , COMP_LOOP_COMP_LOOP_or_101_nl , COMP_LOOP_COMP_LOOP_or_102_nl
      , COMP_LOOP_COMP_LOOP_or_103_nl , COMP_LOOP_COMP_LOOP_or_104_nl , COMP_LOOP_COMP_LOOP_or_105_nl
      , COMP_LOOP_or_37_nl , COMP_LOOP_or_38_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[65:0];
  assign z_out_1 = readslicef_66_65_1(acc_1_nl);
  assign and_434_cse = (fsm_output==9'b011111101);
  assign COMP_LOOP_mux_87_nl = MUX_v_11_2_2((VEC_LOOP_j_1_12_0_sva_11_0[11:1]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:1]),
      and_434_cse);
  assign nl_z_out_2 = COMP_LOOP_mux_87_nl + conv_u2u_8_11(COMP_LOOP_k_9_1_1_sva_7_0);
  assign z_out_2 = nl_z_out_2[10:0];
  assign operator_64_false_1_operator_64_false_1_or_1_nl = (~(and_387_ssc | and_392_ssc))
      | and_379_ssc | and_396_ssc;
  assign operator_64_false_1_mux1h_9_nl = MUX1HOT_s_1_3_2(modExp_exp_1_7_1_sva, (~
      (COMP_LOOP_k_9_1_1_sva_7_0[7])), modExp_exp_1_1_1_sva, {and_379_ssc , and_392_ssc
      , and_396_ssc});
  assign operator_64_false_1_operator_64_false_1_nor_4_nl = ~(operator_64_false_1_mux1h_9_nl
      | and_387_ssc);
  assign operator_64_false_1_mux1h_10_nl = MUX1HOT_s_1_3_2(modExp_exp_1_6_1_sva,
      (~ (COMP_LOOP_k_9_1_1_sva_7_0[6])), modExp_exp_1_7_1_sva, {and_379_ssc , and_392_ssc
      , and_396_ssc});
  assign operator_64_false_1_operator_64_false_1_nor_5_nl = ~(operator_64_false_1_mux1h_10_nl
      | and_387_ssc);
  assign operator_64_false_1_mux1h_11_nl = MUX1HOT_s_1_3_2(modExp_exp_1_5_1_sva,
      (~ (COMP_LOOP_k_9_1_1_sva_7_0[5])), modExp_exp_1_6_1_sva, {and_379_ssc , and_392_ssc
      , and_396_ssc});
  assign operator_64_false_1_operator_64_false_1_nor_6_nl = ~(operator_64_false_1_mux1h_11_nl
      | and_387_ssc);
  assign operator_64_false_1_mux1h_12_nl = MUX1HOT_s_1_3_2(modExp_exp_1_4_1_sva,
      (~ (COMP_LOOP_k_9_1_1_sva_7_0[4])), modExp_exp_1_5_1_sva, {and_379_ssc , and_392_ssc
      , and_396_ssc});
  assign operator_64_false_1_operator_64_false_1_nor_7_nl = ~(operator_64_false_1_mux1h_12_nl
      | and_387_ssc);
  assign operator_64_false_1_mux1h_13_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_3_1_sva),
      (STAGE_LOOP_i_3_0_sva[3]), (COMP_LOOP_k_9_1_1_sva_7_0[3]), (~ modExp_exp_1_4_1_sva),
      {and_379_ssc , and_387_ssc , and_392_ssc , and_396_ssc});
  assign operator_64_false_1_mux1h_14_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_2_1_sva),
      (STAGE_LOOP_i_3_0_sva[2]), (COMP_LOOP_k_9_1_1_sva_7_0[2]), (~ modExp_exp_1_3_1_sva),
      {and_379_ssc , and_387_ssc , and_392_ssc , and_396_ssc});
  assign operator_64_false_1_mux1h_15_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_1_1_sva),
      (STAGE_LOOP_i_3_0_sva[1]), (COMP_LOOP_k_9_1_1_sva_7_0[1]), (~ modExp_exp_1_2_1_sva),
      {and_379_ssc , and_387_ssc , and_392_ssc , and_396_ssc});
  assign operator_64_false_1_or_2_nl = and_379_ssc | and_396_ssc;
  assign operator_64_false_1_mux1h_16_nl = MUX1HOT_s_1_3_2((~ modExp_exp_1_0_1_sva_1),
      (STAGE_LOOP_i_3_0_sva[0]), (COMP_LOOP_k_9_1_1_sva_7_0[0]), {operator_64_false_1_or_2_nl
      , and_387_ssc , and_392_ssc});
  assign nl_z_out_4 = ({operator_64_false_1_operator_64_false_1_or_1_nl , operator_64_false_1_operator_64_false_1_nor_4_nl
      , operator_64_false_1_operator_64_false_1_nor_5_nl , operator_64_false_1_operator_64_false_1_nor_6_nl
      , operator_64_false_1_operator_64_false_1_nor_7_nl , operator_64_false_1_mux1h_13_nl
      , operator_64_false_1_mux1h_14_nl , operator_64_false_1_mux1h_15_nl , operator_64_false_1_mux1h_16_nl})
      + 9'b000000001;
  assign z_out_4 = nl_z_out_4[8:0];
  assign and_436_nl = (fsm_output[3]) & (~ (fsm_output[8])) & (~ (fsm_output[4]))
      & and_dcpl_159 & (~ (fsm_output[6])) & (fsm_output[1]) & and_dcpl_164;
  assign nor_405_nl = ~((fsm_output[3]) | (fsm_output[6]) | (~ nor_tmp_146));
  assign nor_406_nl = ~((~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[5]) |
      (fsm_output[2]));
  assign mux_558_nl = MUX_s_1_2_2(nor_405_nl, nor_406_nl, fsm_output[7]);
  assign nand_129_nl = ~((fsm_output[4]) & mux_558_nl);
  assign nor_407_nl = ~((fsm_output[5]) | (fsm_output[2]));
  assign mux_559_nl = MUX_s_1_2_2(nor_407_nl, nor_tmp_146, fsm_output[6]);
  assign or_713_nl = (fsm_output[4]) | (fsm_output[7]) | (fsm_output[3]) | (~ mux_559_nl);
  assign mux_557_nl = MUX_s_1_2_2(nand_129_nl, or_713_nl, fsm_output[8]);
  assign nor_404_nl = ~((fsm_output[0]) | mux_557_nl);
  assign nor_408_nl = ~((~ (fsm_output[0])) | (fsm_output[8]) | (fsm_output[4]) |
      (fsm_output[7]) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[5]) |
      (fsm_output[2]));
  assign mux_556_nl = MUX_s_1_2_2(nor_404_nl, nor_408_nl, fsm_output[1]);
  assign nor_409_nl = ~((fsm_output[5]) | (fsm_output[2]) | (~ (fsm_output[6])) |
      (fsm_output[3]) | not_tmp_20);
  assign or_714_nl = (fsm_output[6]) | not_tmp_368;
  assign or_715_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[0])
      | (fsm_output[7]);
  assign mux_563_nl = MUX_s_1_2_2(or_714_nl, or_715_nl, fsm_output[2]);
  assign nor_410_nl = ~((fsm_output[5]) | mux_563_nl);
  assign mux_562_nl = MUX_s_1_2_2(nor_409_nl, nor_410_nl, fsm_output[4]);
  assign or_716_nl = (~ (fsm_output[2])) | (fsm_output[6]) | not_tmp_368;
  assign or_717_nl = (fsm_output[6]) | (~ (fsm_output[3])) | (fsm_output[0]) | (fsm_output[7]);
  assign or_718_nl = (~ (fsm_output[6])) | (fsm_output[3]) | (~ (fsm_output[0]))
      | (fsm_output[7]);
  assign mux_565_nl = MUX_s_1_2_2(or_717_nl, or_718_nl, fsm_output[2]);
  assign mux_564_nl = MUX_s_1_2_2(or_716_nl, mux_565_nl, fsm_output[5]);
  assign nor_411_nl = ~((fsm_output[4]) | mux_564_nl);
  assign mux_561_nl = MUX_s_1_2_2(mux_562_nl, nor_411_nl, fsm_output[8]);
  assign nor_413_nl = ~((fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[0])) |
      (fsm_output[7]));
  assign and_437_nl = (fsm_output[6]) & (fsm_output[3]) & (fsm_output[0]) & (fsm_output[7]);
  assign mux_566_nl = MUX_s_1_2_2(nor_413_nl, and_437_nl, fsm_output[2]);
  assign nor_412_nl = ~((fsm_output[8]) | (~((fsm_output[5:4]==2'b11) & mux_566_nl)));
  assign mux_560_nl = MUX_s_1_2_2(mux_561_nl, nor_412_nl, fsm_output[1]);
  assign modExp_while_if_mux1h_2_nl = MUX1HOT_v_64_3_2(modExp_result_sva, COMP_LOOP_mux1h_1_itm,
      operator_64_false_acc_mut_63_0, {and_436_nl , mux_556_nl , mux_560_nl});
  assign nl_z_out_5 = modExp_while_if_mux1h_2_nl * COMP_LOOP_mux1h_1_itm;
  assign z_out_5 = nl_z_out_5[63:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_6_2;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [5:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    MUX1HOT_v_10_6_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_9_2;
    input [9:0] input_8;
    input [9:0] input_7;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [8:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    result = result | ( input_6 & {10{sel[6]}});
    result = result | ( input_7 & {10{sel[7]}});
    result = result | ( input_8 & {10{sel[8]}});
    MUX1HOT_v_10_9_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_5_2;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [4:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    result = result | ( input_4 & {2{sel[4]}});
    MUX1HOT_v_2_5_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_3_2;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [2:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | ( input_1 & {51{sel[1]}});
    result = result | ( input_2 & {51{sel[2]}});
    MUX1HOT_v_51_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_10_2;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [9:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    MUX1HOT_v_64_10_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_5_2;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [4:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    MUX1HOT_v_64_5_2 = result;
  end
  endfunction


  function automatic [64:0] MUX1HOT_v_65_3_2;
    input [64:0] input_2;
    input [64:0] input_1;
    input [64:0] input_0;
    input [2:0] sel;
    reg [64:0] result;
  begin
    result = input_0 & {65{sel[0]}};
    result = result | ( input_1 & {65{sel[1]}});
    result = result | ( input_2 & {65{sel[2]}});
    MUX1HOT_v_65_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [50:0] MUX_v_51_2_2;
    input [50:0] input_0;
    input [50:0] input_1;
    input [0:0] sel;
    reg [50:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_51_2_2 = result;
  end
  endfunction


  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [0:0] readslicef_65_1_64;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 64;
    readslicef_65_1_64 = tmp[0:0];
  end
  endfunction


  function automatic [64:0] readslicef_66_65_1;
    input [65:0] vector;
    reg [65:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_66_65_1 = tmp[64:0];
  end
  endfunction


  function automatic [65:0] conv_s2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_s2u_65_66 = {vector[64], vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_11 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [65:0] conv_u2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_u2u_65_66 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      vec_rsc_0_2_adra, vec_rsc_0_2_da, vec_rsc_0_2_wea, vec_rsc_0_2_qa, vec_rsc_triosy_0_2_lz,
      vec_rsc_0_3_adra, vec_rsc_0_3_da, vec_rsc_0_3_wea, vec_rsc_0_3_qa, vec_rsc_triosy_0_3_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [9:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [9:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  output [9:0] vec_rsc_0_2_adra;
  output [63:0] vec_rsc_0_2_da;
  output vec_rsc_0_2_wea;
  input [63:0] vec_rsc_0_2_qa;
  output vec_rsc_triosy_0_2_lz;
  output [9:0] vec_rsc_0_3_adra;
  output [63:0] vec_rsc_0_3_da;
  output vec_rsc_0_3_wea;
  input [63:0] vec_rsc_0_3_qa;
  output vec_rsc_triosy_0_3_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_qa_d;
  wire vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_qa_d;
  wire vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;
  wire vec_rsc_0_2_i_wea_d_iff;
  wire vec_rsc_0_3_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
      vec_rsc_0_0_i (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
      vec_rsc_0_1_i (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
      vec_rsc_0_2_i (
      .qa(vec_rsc_0_2_qa),
      .wea(vec_rsc_0_2_wea),
      .da(vec_rsc_0_2_da),
      .adra(vec_rsc_0_2_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_2_i_qa_d),
      .wea_d(vec_rsc_0_2_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
      vec_rsc_0_3_i (
      .qa(vec_rsc_0_3_qa),
      .wea(vec_rsc_0_3_wea),
      .da(vec_rsc_0_3_da),
      .adra(vec_rsc_0_3_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_3_i_qa_d),
      .wea_d(vec_rsc_0_3_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_wea_d_iff)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_qa_d(vec_rsc_0_2_i_qa_d),
      .vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_qa_d(vec_rsc_0_3_i_qa_d),
      .vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff),
      .vec_rsc_0_2_i_wea_d_pff(vec_rsc_0_2_i_wea_d_iff),
      .vec_rsc_0_3_i_wea_d_pff(vec_rsc_0_3_i_wea_d_iff)
    );
endmodule



