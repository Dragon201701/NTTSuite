
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ../td_ccore_solutions/modulo_dev_0dc217f8ce5f309b848fa994f59fa3f66234_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Wed Aug 18 22:11:42 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    modulo_dev_core
// ------------------------------------------------------------------


module modulo_dev_core (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [63:0] base_rsci_idat;
  wire [63:0] m_rsci_idat;
  reg [63:0] return_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire [64:0] rem_2_cmp_z;
  wire [64:0] rem_2_cmp_1_z;
  reg [63:0] rem_2_cmp_b_63_0;
  reg [63:0] rem_2_cmp_1_b_63_0;
  reg [63:0] rem_2_cmp_a_63_0;
  reg [63:0] rem_2_cmp_1_a_63_0;
  wire and_dcpl;
  reg rem_2cyc;
  reg rem_2cyc_st_2;
  reg [63:0] result_sva_1;
  wire and_3_cse;
  wire and_5_cse;
  reg main_stage_0_2;
  reg main_stage_0_3;
  reg [63:0] m_buf_sva_1;
  reg [63:0] m_buf_sva_2;
  reg [63:0] m_buf_sva_3;
  reg asn_itm_1;
  reg asn_itm_2;
  wire and_8_cse;
  wire and_7_cse;

  wire[63:0] qelse_acc_nl;
  wire[64:0] nl_qelse_acc_nl;
  wire[0:0] mux_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [64:0] nl_rem_2_cmp_a;
  assign nl_rem_2_cmp_a = {{1{rem_2_cmp_a_63_0[63]}}, rem_2_cmp_a_63_0};
  wire [64:0] nl_rem_2_cmp_b;
  assign nl_rem_2_cmp_b = {1'b0 , rem_2_cmp_b_63_0};
  wire [64:0] nl_rem_2_cmp_1_a;
  assign nl_rem_2_cmp_1_a = {{1{rem_2_cmp_1_a_63_0[63]}}, rem_2_cmp_1_a_63_0};
  wire [64:0] nl_rem_2_cmp_1_b;
  assign nl_rem_2_cmp_1_b = {1'b0 , rem_2_cmp_1_b_63_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) base_rsci (
      .dat(base_rsc_dat),
      .idat(base_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .d(return_rsci_d),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_2_cmp (
      .a(nl_rem_2_cmp_a[64:0]),
      .b(nl_rem_2_cmp_b[64:0]),
      .z(rem_2_cmp_z)
    );
  mgc_rem #(.width_a(32'sd65),
  .width_b(32'sd65),
  .signd(32'sd1)) rem_2_cmp_1 (
      .a(nl_rem_2_cmp_1_a[64:0]),
      .b(nl_rem_2_cmp_1_b[64:0]),
      .z(rem_2_cmp_1_z)
    );
  assign and_8_cse = ccs_ccore_en & main_stage_0_2 & asn_itm_1;
  assign and_3_cse = ccs_ccore_en & rem_2cyc;
  assign and_5_cse = ccs_ccore_en & (~ rem_2cyc);
  assign and_7_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  assign and_dcpl = main_stage_0_3 & asn_itm_2;
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      return_rsci_d <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      asn_itm_2 <= 1'b0;
      asn_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
    end
    else if ( ccs_ccore_en ) begin
      return_rsci_d <= MUX_v_64_2_2(result_sva_1, qelse_acc_nl, result_sva_1[63]);
      asn_itm_2 <= asn_itm_1;
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_sva_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ccs_ccore_en & and_dcpl ) begin
      result_sva_1 <= MUX_v_64_2_2((rem_2_cmp_1_z[63:0]), (rem_2_cmp_z[63:0]), rem_2cyc_st_2);
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      m_buf_sva_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ccs_ccore_en & mux_2_nl & and_dcpl ) begin
      m_buf_sva_3 <= m_buf_sva_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_2cyc_st_2 <= 1'b0;
      m_buf_sva_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_8_cse ) begin
      rem_2cyc_st_2 <= rem_2cyc;
      m_buf_sva_2 <= m_buf_sva_1;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_2_cmp_1_b_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rem_2_cmp_1_a_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_3_cse ) begin
      rem_2_cmp_1_b_63_0 <= m_rsci_idat;
      rem_2_cmp_1_a_63_0 <= base_rsci_idat;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_2_cmp_b_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rem_2_cmp_a_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_5_cse ) begin
      rem_2_cmp_b_63_0 <= m_rsci_idat;
      rem_2_cmp_a_63_0 <= base_rsci_idat;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      rem_2cyc <= 1'b0;
      m_buf_sva_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_7_cse ) begin
      rem_2cyc <= ~ rem_2cyc;
      m_buf_sva_1 <= m_rsci_idat;
    end
  end
  assign nl_qelse_acc_nl = result_sva_1 + m_buf_sva_3;
  assign qelse_acc_nl = nl_qelse_acc_nl[63:0];
  assign mux_2_nl = MUX_s_1_2_2((rem_2_cmp_1_z[63]), (rem_2_cmp_z[63]), rem_2cyc_st_2);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    modulo_dev
// ------------------------------------------------------------------


module modulo_dev (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  modulo_dev_core modulo_dev_core_inst (
      .base_rsc_dat(base_rsc_dat),
      .m_rsc_dat(m_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v5.v 
module mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Thu Aug 19 00:32:38 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_24_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_24_64_7_128_128_64_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_23_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_23_64_7_128_128_64_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_22_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_22_64_7_128_128_64_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_21_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_21_64_7_128_128_64_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_20_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_20_64_7_128_128_64_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_19_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_19_64_7_128_128_64_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_18_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_18_64_7_128_128_64_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_17_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_17_64_7_128_128_64_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_16_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_16_64_7_128_128_64_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [63:0] d;
  output [6:0] wadr;
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [63:0] d_d;
  input we_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_15_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_15_64_7_128_128_64_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [63:0] d;
  output [6:0] wadr;
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [63:0] d_d;
  input we_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_14_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_14_64_7_128_128_64_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [63:0] d;
  output [6:0] wadr;
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [63:0] d_d;
  input we_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_13_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_13_64_7_128_128_64_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [63:0] d;
  output [6:0] wadr;
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [63:0] d_d;
  input we_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_12_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_12_64_7_128_128_64_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [63:0] d;
  output [6:0] wadr;
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [63:0] d_d;
  input we_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_11_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_11_64_7_128_128_64_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [63:0] d;
  output [6:0] wadr;
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [63:0] d_d;
  input we_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_10_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_10_64_7_128_128_64_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [63:0] d;
  output [6:0] wadr;
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [63:0] d_d;
  input we_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_9_64_7_128_128_64_5_gen
// ------------------------------------------------------------------


module DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_9_64_7_128_128_64_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [63:0] d;
  output [6:0] wadr;
  input [63:0] q;
  output re;
  output [6:0] radr;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input [63:0] d_d;
  input we_d;
  input re_d;
  output [63:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module DIT_RELOOP_core_core_fsm (
  clk, rst, fsm_output, IDX_LOOP_C_33_tr0, IDX_LOOP_C_65_tr0, IDX_LOOP_C_97_tr0,
      IDX_LOOP_C_129_tr0, IDX_LOOP_C_161_tr0, IDX_LOOP_C_193_tr0, IDX_LOOP_C_225_tr0,
      IDX_LOOP_C_257_tr0, GROUP_LOOP_C_0_tr0, STAGE_LOOP_C_1_tr0
);
  input clk;
  input rst;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input IDX_LOOP_C_33_tr0;
  input IDX_LOOP_C_65_tr0;
  input IDX_LOOP_C_97_tr0;
  input IDX_LOOP_C_129_tr0;
  input IDX_LOOP_C_161_tr0;
  input IDX_LOOP_C_193_tr0;
  input IDX_LOOP_C_225_tr0;
  input IDX_LOOP_C_257_tr0;
  input GROUP_LOOP_C_0_tr0;
  input STAGE_LOOP_C_1_tr0;


  // FSM State Type Declaration for DIT_RELOOP_core_core_fsm_1
  parameter
    main_C_0 = 9'd0,
    STAGE_LOOP_C_0 = 9'd1,
    IDX_LOOP_C_0 = 9'd2,
    IDX_LOOP_C_1 = 9'd3,
    IDX_LOOP_C_2 = 9'd4,
    IDX_LOOP_C_3 = 9'd5,
    IDX_LOOP_C_4 = 9'd6,
    IDX_LOOP_C_5 = 9'd7,
    IDX_LOOP_C_6 = 9'd8,
    IDX_LOOP_C_7 = 9'd9,
    IDX_LOOP_C_8 = 9'd10,
    IDX_LOOP_C_9 = 9'd11,
    IDX_LOOP_C_10 = 9'd12,
    IDX_LOOP_C_11 = 9'd13,
    IDX_LOOP_C_12 = 9'd14,
    IDX_LOOP_C_13 = 9'd15,
    IDX_LOOP_C_14 = 9'd16,
    IDX_LOOP_C_15 = 9'd17,
    IDX_LOOP_C_16 = 9'd18,
    IDX_LOOP_C_17 = 9'd19,
    IDX_LOOP_C_18 = 9'd20,
    IDX_LOOP_C_19 = 9'd21,
    IDX_LOOP_C_20 = 9'd22,
    IDX_LOOP_C_21 = 9'd23,
    IDX_LOOP_C_22 = 9'd24,
    IDX_LOOP_C_23 = 9'd25,
    IDX_LOOP_C_24 = 9'd26,
    IDX_LOOP_C_25 = 9'd27,
    IDX_LOOP_C_26 = 9'd28,
    IDX_LOOP_C_27 = 9'd29,
    IDX_LOOP_C_28 = 9'd30,
    IDX_LOOP_C_29 = 9'd31,
    IDX_LOOP_C_30 = 9'd32,
    IDX_LOOP_C_31 = 9'd33,
    IDX_LOOP_C_32 = 9'd34,
    IDX_LOOP_C_33 = 9'd35,
    IDX_LOOP_C_34 = 9'd36,
    IDX_LOOP_C_35 = 9'd37,
    IDX_LOOP_C_36 = 9'd38,
    IDX_LOOP_C_37 = 9'd39,
    IDX_LOOP_C_38 = 9'd40,
    IDX_LOOP_C_39 = 9'd41,
    IDX_LOOP_C_40 = 9'd42,
    IDX_LOOP_C_41 = 9'd43,
    IDX_LOOP_C_42 = 9'd44,
    IDX_LOOP_C_43 = 9'd45,
    IDX_LOOP_C_44 = 9'd46,
    IDX_LOOP_C_45 = 9'd47,
    IDX_LOOP_C_46 = 9'd48,
    IDX_LOOP_C_47 = 9'd49,
    IDX_LOOP_C_48 = 9'd50,
    IDX_LOOP_C_49 = 9'd51,
    IDX_LOOP_C_50 = 9'd52,
    IDX_LOOP_C_51 = 9'd53,
    IDX_LOOP_C_52 = 9'd54,
    IDX_LOOP_C_53 = 9'd55,
    IDX_LOOP_C_54 = 9'd56,
    IDX_LOOP_C_55 = 9'd57,
    IDX_LOOP_C_56 = 9'd58,
    IDX_LOOP_C_57 = 9'd59,
    IDX_LOOP_C_58 = 9'd60,
    IDX_LOOP_C_59 = 9'd61,
    IDX_LOOP_C_60 = 9'd62,
    IDX_LOOP_C_61 = 9'd63,
    IDX_LOOP_C_62 = 9'd64,
    IDX_LOOP_C_63 = 9'd65,
    IDX_LOOP_C_64 = 9'd66,
    IDX_LOOP_C_65 = 9'd67,
    IDX_LOOP_C_66 = 9'd68,
    IDX_LOOP_C_67 = 9'd69,
    IDX_LOOP_C_68 = 9'd70,
    IDX_LOOP_C_69 = 9'd71,
    IDX_LOOP_C_70 = 9'd72,
    IDX_LOOP_C_71 = 9'd73,
    IDX_LOOP_C_72 = 9'd74,
    IDX_LOOP_C_73 = 9'd75,
    IDX_LOOP_C_74 = 9'd76,
    IDX_LOOP_C_75 = 9'd77,
    IDX_LOOP_C_76 = 9'd78,
    IDX_LOOP_C_77 = 9'd79,
    IDX_LOOP_C_78 = 9'd80,
    IDX_LOOP_C_79 = 9'd81,
    IDX_LOOP_C_80 = 9'd82,
    IDX_LOOP_C_81 = 9'd83,
    IDX_LOOP_C_82 = 9'd84,
    IDX_LOOP_C_83 = 9'd85,
    IDX_LOOP_C_84 = 9'd86,
    IDX_LOOP_C_85 = 9'd87,
    IDX_LOOP_C_86 = 9'd88,
    IDX_LOOP_C_87 = 9'd89,
    IDX_LOOP_C_88 = 9'd90,
    IDX_LOOP_C_89 = 9'd91,
    IDX_LOOP_C_90 = 9'd92,
    IDX_LOOP_C_91 = 9'd93,
    IDX_LOOP_C_92 = 9'd94,
    IDX_LOOP_C_93 = 9'd95,
    IDX_LOOP_C_94 = 9'd96,
    IDX_LOOP_C_95 = 9'd97,
    IDX_LOOP_C_96 = 9'd98,
    IDX_LOOP_C_97 = 9'd99,
    IDX_LOOP_C_98 = 9'd100,
    IDX_LOOP_C_99 = 9'd101,
    IDX_LOOP_C_100 = 9'd102,
    IDX_LOOP_C_101 = 9'd103,
    IDX_LOOP_C_102 = 9'd104,
    IDX_LOOP_C_103 = 9'd105,
    IDX_LOOP_C_104 = 9'd106,
    IDX_LOOP_C_105 = 9'd107,
    IDX_LOOP_C_106 = 9'd108,
    IDX_LOOP_C_107 = 9'd109,
    IDX_LOOP_C_108 = 9'd110,
    IDX_LOOP_C_109 = 9'd111,
    IDX_LOOP_C_110 = 9'd112,
    IDX_LOOP_C_111 = 9'd113,
    IDX_LOOP_C_112 = 9'd114,
    IDX_LOOP_C_113 = 9'd115,
    IDX_LOOP_C_114 = 9'd116,
    IDX_LOOP_C_115 = 9'd117,
    IDX_LOOP_C_116 = 9'd118,
    IDX_LOOP_C_117 = 9'd119,
    IDX_LOOP_C_118 = 9'd120,
    IDX_LOOP_C_119 = 9'd121,
    IDX_LOOP_C_120 = 9'd122,
    IDX_LOOP_C_121 = 9'd123,
    IDX_LOOP_C_122 = 9'd124,
    IDX_LOOP_C_123 = 9'd125,
    IDX_LOOP_C_124 = 9'd126,
    IDX_LOOP_C_125 = 9'd127,
    IDX_LOOP_C_126 = 9'd128,
    IDX_LOOP_C_127 = 9'd129,
    IDX_LOOP_C_128 = 9'd130,
    IDX_LOOP_C_129 = 9'd131,
    IDX_LOOP_C_130 = 9'd132,
    IDX_LOOP_C_131 = 9'd133,
    IDX_LOOP_C_132 = 9'd134,
    IDX_LOOP_C_133 = 9'd135,
    IDX_LOOP_C_134 = 9'd136,
    IDX_LOOP_C_135 = 9'd137,
    IDX_LOOP_C_136 = 9'd138,
    IDX_LOOP_C_137 = 9'd139,
    IDX_LOOP_C_138 = 9'd140,
    IDX_LOOP_C_139 = 9'd141,
    IDX_LOOP_C_140 = 9'd142,
    IDX_LOOP_C_141 = 9'd143,
    IDX_LOOP_C_142 = 9'd144,
    IDX_LOOP_C_143 = 9'd145,
    IDX_LOOP_C_144 = 9'd146,
    IDX_LOOP_C_145 = 9'd147,
    IDX_LOOP_C_146 = 9'd148,
    IDX_LOOP_C_147 = 9'd149,
    IDX_LOOP_C_148 = 9'd150,
    IDX_LOOP_C_149 = 9'd151,
    IDX_LOOP_C_150 = 9'd152,
    IDX_LOOP_C_151 = 9'd153,
    IDX_LOOP_C_152 = 9'd154,
    IDX_LOOP_C_153 = 9'd155,
    IDX_LOOP_C_154 = 9'd156,
    IDX_LOOP_C_155 = 9'd157,
    IDX_LOOP_C_156 = 9'd158,
    IDX_LOOP_C_157 = 9'd159,
    IDX_LOOP_C_158 = 9'd160,
    IDX_LOOP_C_159 = 9'd161,
    IDX_LOOP_C_160 = 9'd162,
    IDX_LOOP_C_161 = 9'd163,
    IDX_LOOP_C_162 = 9'd164,
    IDX_LOOP_C_163 = 9'd165,
    IDX_LOOP_C_164 = 9'd166,
    IDX_LOOP_C_165 = 9'd167,
    IDX_LOOP_C_166 = 9'd168,
    IDX_LOOP_C_167 = 9'd169,
    IDX_LOOP_C_168 = 9'd170,
    IDX_LOOP_C_169 = 9'd171,
    IDX_LOOP_C_170 = 9'd172,
    IDX_LOOP_C_171 = 9'd173,
    IDX_LOOP_C_172 = 9'd174,
    IDX_LOOP_C_173 = 9'd175,
    IDX_LOOP_C_174 = 9'd176,
    IDX_LOOP_C_175 = 9'd177,
    IDX_LOOP_C_176 = 9'd178,
    IDX_LOOP_C_177 = 9'd179,
    IDX_LOOP_C_178 = 9'd180,
    IDX_LOOP_C_179 = 9'd181,
    IDX_LOOP_C_180 = 9'd182,
    IDX_LOOP_C_181 = 9'd183,
    IDX_LOOP_C_182 = 9'd184,
    IDX_LOOP_C_183 = 9'd185,
    IDX_LOOP_C_184 = 9'd186,
    IDX_LOOP_C_185 = 9'd187,
    IDX_LOOP_C_186 = 9'd188,
    IDX_LOOP_C_187 = 9'd189,
    IDX_LOOP_C_188 = 9'd190,
    IDX_LOOP_C_189 = 9'd191,
    IDX_LOOP_C_190 = 9'd192,
    IDX_LOOP_C_191 = 9'd193,
    IDX_LOOP_C_192 = 9'd194,
    IDX_LOOP_C_193 = 9'd195,
    IDX_LOOP_C_194 = 9'd196,
    IDX_LOOP_C_195 = 9'd197,
    IDX_LOOP_C_196 = 9'd198,
    IDX_LOOP_C_197 = 9'd199,
    IDX_LOOP_C_198 = 9'd200,
    IDX_LOOP_C_199 = 9'd201,
    IDX_LOOP_C_200 = 9'd202,
    IDX_LOOP_C_201 = 9'd203,
    IDX_LOOP_C_202 = 9'd204,
    IDX_LOOP_C_203 = 9'd205,
    IDX_LOOP_C_204 = 9'd206,
    IDX_LOOP_C_205 = 9'd207,
    IDX_LOOP_C_206 = 9'd208,
    IDX_LOOP_C_207 = 9'd209,
    IDX_LOOP_C_208 = 9'd210,
    IDX_LOOP_C_209 = 9'd211,
    IDX_LOOP_C_210 = 9'd212,
    IDX_LOOP_C_211 = 9'd213,
    IDX_LOOP_C_212 = 9'd214,
    IDX_LOOP_C_213 = 9'd215,
    IDX_LOOP_C_214 = 9'd216,
    IDX_LOOP_C_215 = 9'd217,
    IDX_LOOP_C_216 = 9'd218,
    IDX_LOOP_C_217 = 9'd219,
    IDX_LOOP_C_218 = 9'd220,
    IDX_LOOP_C_219 = 9'd221,
    IDX_LOOP_C_220 = 9'd222,
    IDX_LOOP_C_221 = 9'd223,
    IDX_LOOP_C_222 = 9'd224,
    IDX_LOOP_C_223 = 9'd225,
    IDX_LOOP_C_224 = 9'd226,
    IDX_LOOP_C_225 = 9'd227,
    IDX_LOOP_C_226 = 9'd228,
    IDX_LOOP_C_227 = 9'd229,
    IDX_LOOP_C_228 = 9'd230,
    IDX_LOOP_C_229 = 9'd231,
    IDX_LOOP_C_230 = 9'd232,
    IDX_LOOP_C_231 = 9'd233,
    IDX_LOOP_C_232 = 9'd234,
    IDX_LOOP_C_233 = 9'd235,
    IDX_LOOP_C_234 = 9'd236,
    IDX_LOOP_C_235 = 9'd237,
    IDX_LOOP_C_236 = 9'd238,
    IDX_LOOP_C_237 = 9'd239,
    IDX_LOOP_C_238 = 9'd240,
    IDX_LOOP_C_239 = 9'd241,
    IDX_LOOP_C_240 = 9'd242,
    IDX_LOOP_C_241 = 9'd243,
    IDX_LOOP_C_242 = 9'd244,
    IDX_LOOP_C_243 = 9'd245,
    IDX_LOOP_C_244 = 9'd246,
    IDX_LOOP_C_245 = 9'd247,
    IDX_LOOP_C_246 = 9'd248,
    IDX_LOOP_C_247 = 9'd249,
    IDX_LOOP_C_248 = 9'd250,
    IDX_LOOP_C_249 = 9'd251,
    IDX_LOOP_C_250 = 9'd252,
    IDX_LOOP_C_251 = 9'd253,
    IDX_LOOP_C_252 = 9'd254,
    IDX_LOOP_C_253 = 9'd255,
    IDX_LOOP_C_254 = 9'd256,
    IDX_LOOP_C_255 = 9'd257,
    IDX_LOOP_C_256 = 9'd258,
    IDX_LOOP_C_257 = 9'd259,
    GROUP_LOOP_C_0 = 9'd260,
    STAGE_LOOP_C_1 = 9'd261,
    main_C_1 = 9'd262;

  reg [8:0] state_var;
  reg [8:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : DIT_RELOOP_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 9'b000000001;
        state_var_NS = IDX_LOOP_C_0;
      end
      IDX_LOOP_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = IDX_LOOP_C_1;
      end
      IDX_LOOP_C_1 : begin
        fsm_output = 9'b000000011;
        state_var_NS = IDX_LOOP_C_2;
      end
      IDX_LOOP_C_2 : begin
        fsm_output = 9'b000000100;
        state_var_NS = IDX_LOOP_C_3;
      end
      IDX_LOOP_C_3 : begin
        fsm_output = 9'b000000101;
        state_var_NS = IDX_LOOP_C_4;
      end
      IDX_LOOP_C_4 : begin
        fsm_output = 9'b000000110;
        state_var_NS = IDX_LOOP_C_5;
      end
      IDX_LOOP_C_5 : begin
        fsm_output = 9'b000000111;
        state_var_NS = IDX_LOOP_C_6;
      end
      IDX_LOOP_C_6 : begin
        fsm_output = 9'b000001000;
        state_var_NS = IDX_LOOP_C_7;
      end
      IDX_LOOP_C_7 : begin
        fsm_output = 9'b000001001;
        state_var_NS = IDX_LOOP_C_8;
      end
      IDX_LOOP_C_8 : begin
        fsm_output = 9'b000001010;
        state_var_NS = IDX_LOOP_C_9;
      end
      IDX_LOOP_C_9 : begin
        fsm_output = 9'b000001011;
        state_var_NS = IDX_LOOP_C_10;
      end
      IDX_LOOP_C_10 : begin
        fsm_output = 9'b000001100;
        state_var_NS = IDX_LOOP_C_11;
      end
      IDX_LOOP_C_11 : begin
        fsm_output = 9'b000001101;
        state_var_NS = IDX_LOOP_C_12;
      end
      IDX_LOOP_C_12 : begin
        fsm_output = 9'b000001110;
        state_var_NS = IDX_LOOP_C_13;
      end
      IDX_LOOP_C_13 : begin
        fsm_output = 9'b000001111;
        state_var_NS = IDX_LOOP_C_14;
      end
      IDX_LOOP_C_14 : begin
        fsm_output = 9'b000010000;
        state_var_NS = IDX_LOOP_C_15;
      end
      IDX_LOOP_C_15 : begin
        fsm_output = 9'b000010001;
        state_var_NS = IDX_LOOP_C_16;
      end
      IDX_LOOP_C_16 : begin
        fsm_output = 9'b000010010;
        state_var_NS = IDX_LOOP_C_17;
      end
      IDX_LOOP_C_17 : begin
        fsm_output = 9'b000010011;
        state_var_NS = IDX_LOOP_C_18;
      end
      IDX_LOOP_C_18 : begin
        fsm_output = 9'b000010100;
        state_var_NS = IDX_LOOP_C_19;
      end
      IDX_LOOP_C_19 : begin
        fsm_output = 9'b000010101;
        state_var_NS = IDX_LOOP_C_20;
      end
      IDX_LOOP_C_20 : begin
        fsm_output = 9'b000010110;
        state_var_NS = IDX_LOOP_C_21;
      end
      IDX_LOOP_C_21 : begin
        fsm_output = 9'b000010111;
        state_var_NS = IDX_LOOP_C_22;
      end
      IDX_LOOP_C_22 : begin
        fsm_output = 9'b000011000;
        state_var_NS = IDX_LOOP_C_23;
      end
      IDX_LOOP_C_23 : begin
        fsm_output = 9'b000011001;
        state_var_NS = IDX_LOOP_C_24;
      end
      IDX_LOOP_C_24 : begin
        fsm_output = 9'b000011010;
        state_var_NS = IDX_LOOP_C_25;
      end
      IDX_LOOP_C_25 : begin
        fsm_output = 9'b000011011;
        state_var_NS = IDX_LOOP_C_26;
      end
      IDX_LOOP_C_26 : begin
        fsm_output = 9'b000011100;
        state_var_NS = IDX_LOOP_C_27;
      end
      IDX_LOOP_C_27 : begin
        fsm_output = 9'b000011101;
        state_var_NS = IDX_LOOP_C_28;
      end
      IDX_LOOP_C_28 : begin
        fsm_output = 9'b000011110;
        state_var_NS = IDX_LOOP_C_29;
      end
      IDX_LOOP_C_29 : begin
        fsm_output = 9'b000011111;
        state_var_NS = IDX_LOOP_C_30;
      end
      IDX_LOOP_C_30 : begin
        fsm_output = 9'b000100000;
        state_var_NS = IDX_LOOP_C_31;
      end
      IDX_LOOP_C_31 : begin
        fsm_output = 9'b000100001;
        state_var_NS = IDX_LOOP_C_32;
      end
      IDX_LOOP_C_32 : begin
        fsm_output = 9'b000100010;
        state_var_NS = IDX_LOOP_C_33;
      end
      IDX_LOOP_C_33 : begin
        fsm_output = 9'b000100011;
        if ( IDX_LOOP_C_33_tr0 ) begin
          state_var_NS = GROUP_LOOP_C_0;
        end
        else begin
          state_var_NS = IDX_LOOP_C_34;
        end
      end
      IDX_LOOP_C_34 : begin
        fsm_output = 9'b000100100;
        state_var_NS = IDX_LOOP_C_35;
      end
      IDX_LOOP_C_35 : begin
        fsm_output = 9'b000100101;
        state_var_NS = IDX_LOOP_C_36;
      end
      IDX_LOOP_C_36 : begin
        fsm_output = 9'b000100110;
        state_var_NS = IDX_LOOP_C_37;
      end
      IDX_LOOP_C_37 : begin
        fsm_output = 9'b000100111;
        state_var_NS = IDX_LOOP_C_38;
      end
      IDX_LOOP_C_38 : begin
        fsm_output = 9'b000101000;
        state_var_NS = IDX_LOOP_C_39;
      end
      IDX_LOOP_C_39 : begin
        fsm_output = 9'b000101001;
        state_var_NS = IDX_LOOP_C_40;
      end
      IDX_LOOP_C_40 : begin
        fsm_output = 9'b000101010;
        state_var_NS = IDX_LOOP_C_41;
      end
      IDX_LOOP_C_41 : begin
        fsm_output = 9'b000101011;
        state_var_NS = IDX_LOOP_C_42;
      end
      IDX_LOOP_C_42 : begin
        fsm_output = 9'b000101100;
        state_var_NS = IDX_LOOP_C_43;
      end
      IDX_LOOP_C_43 : begin
        fsm_output = 9'b000101101;
        state_var_NS = IDX_LOOP_C_44;
      end
      IDX_LOOP_C_44 : begin
        fsm_output = 9'b000101110;
        state_var_NS = IDX_LOOP_C_45;
      end
      IDX_LOOP_C_45 : begin
        fsm_output = 9'b000101111;
        state_var_NS = IDX_LOOP_C_46;
      end
      IDX_LOOP_C_46 : begin
        fsm_output = 9'b000110000;
        state_var_NS = IDX_LOOP_C_47;
      end
      IDX_LOOP_C_47 : begin
        fsm_output = 9'b000110001;
        state_var_NS = IDX_LOOP_C_48;
      end
      IDX_LOOP_C_48 : begin
        fsm_output = 9'b000110010;
        state_var_NS = IDX_LOOP_C_49;
      end
      IDX_LOOP_C_49 : begin
        fsm_output = 9'b000110011;
        state_var_NS = IDX_LOOP_C_50;
      end
      IDX_LOOP_C_50 : begin
        fsm_output = 9'b000110100;
        state_var_NS = IDX_LOOP_C_51;
      end
      IDX_LOOP_C_51 : begin
        fsm_output = 9'b000110101;
        state_var_NS = IDX_LOOP_C_52;
      end
      IDX_LOOP_C_52 : begin
        fsm_output = 9'b000110110;
        state_var_NS = IDX_LOOP_C_53;
      end
      IDX_LOOP_C_53 : begin
        fsm_output = 9'b000110111;
        state_var_NS = IDX_LOOP_C_54;
      end
      IDX_LOOP_C_54 : begin
        fsm_output = 9'b000111000;
        state_var_NS = IDX_LOOP_C_55;
      end
      IDX_LOOP_C_55 : begin
        fsm_output = 9'b000111001;
        state_var_NS = IDX_LOOP_C_56;
      end
      IDX_LOOP_C_56 : begin
        fsm_output = 9'b000111010;
        state_var_NS = IDX_LOOP_C_57;
      end
      IDX_LOOP_C_57 : begin
        fsm_output = 9'b000111011;
        state_var_NS = IDX_LOOP_C_58;
      end
      IDX_LOOP_C_58 : begin
        fsm_output = 9'b000111100;
        state_var_NS = IDX_LOOP_C_59;
      end
      IDX_LOOP_C_59 : begin
        fsm_output = 9'b000111101;
        state_var_NS = IDX_LOOP_C_60;
      end
      IDX_LOOP_C_60 : begin
        fsm_output = 9'b000111110;
        state_var_NS = IDX_LOOP_C_61;
      end
      IDX_LOOP_C_61 : begin
        fsm_output = 9'b000111111;
        state_var_NS = IDX_LOOP_C_62;
      end
      IDX_LOOP_C_62 : begin
        fsm_output = 9'b001000000;
        state_var_NS = IDX_LOOP_C_63;
      end
      IDX_LOOP_C_63 : begin
        fsm_output = 9'b001000001;
        state_var_NS = IDX_LOOP_C_64;
      end
      IDX_LOOP_C_64 : begin
        fsm_output = 9'b001000010;
        state_var_NS = IDX_LOOP_C_65;
      end
      IDX_LOOP_C_65 : begin
        fsm_output = 9'b001000011;
        if ( IDX_LOOP_C_65_tr0 ) begin
          state_var_NS = GROUP_LOOP_C_0;
        end
        else begin
          state_var_NS = IDX_LOOP_C_66;
        end
      end
      IDX_LOOP_C_66 : begin
        fsm_output = 9'b001000100;
        state_var_NS = IDX_LOOP_C_67;
      end
      IDX_LOOP_C_67 : begin
        fsm_output = 9'b001000101;
        state_var_NS = IDX_LOOP_C_68;
      end
      IDX_LOOP_C_68 : begin
        fsm_output = 9'b001000110;
        state_var_NS = IDX_LOOP_C_69;
      end
      IDX_LOOP_C_69 : begin
        fsm_output = 9'b001000111;
        state_var_NS = IDX_LOOP_C_70;
      end
      IDX_LOOP_C_70 : begin
        fsm_output = 9'b001001000;
        state_var_NS = IDX_LOOP_C_71;
      end
      IDX_LOOP_C_71 : begin
        fsm_output = 9'b001001001;
        state_var_NS = IDX_LOOP_C_72;
      end
      IDX_LOOP_C_72 : begin
        fsm_output = 9'b001001010;
        state_var_NS = IDX_LOOP_C_73;
      end
      IDX_LOOP_C_73 : begin
        fsm_output = 9'b001001011;
        state_var_NS = IDX_LOOP_C_74;
      end
      IDX_LOOP_C_74 : begin
        fsm_output = 9'b001001100;
        state_var_NS = IDX_LOOP_C_75;
      end
      IDX_LOOP_C_75 : begin
        fsm_output = 9'b001001101;
        state_var_NS = IDX_LOOP_C_76;
      end
      IDX_LOOP_C_76 : begin
        fsm_output = 9'b001001110;
        state_var_NS = IDX_LOOP_C_77;
      end
      IDX_LOOP_C_77 : begin
        fsm_output = 9'b001001111;
        state_var_NS = IDX_LOOP_C_78;
      end
      IDX_LOOP_C_78 : begin
        fsm_output = 9'b001010000;
        state_var_NS = IDX_LOOP_C_79;
      end
      IDX_LOOP_C_79 : begin
        fsm_output = 9'b001010001;
        state_var_NS = IDX_LOOP_C_80;
      end
      IDX_LOOP_C_80 : begin
        fsm_output = 9'b001010010;
        state_var_NS = IDX_LOOP_C_81;
      end
      IDX_LOOP_C_81 : begin
        fsm_output = 9'b001010011;
        state_var_NS = IDX_LOOP_C_82;
      end
      IDX_LOOP_C_82 : begin
        fsm_output = 9'b001010100;
        state_var_NS = IDX_LOOP_C_83;
      end
      IDX_LOOP_C_83 : begin
        fsm_output = 9'b001010101;
        state_var_NS = IDX_LOOP_C_84;
      end
      IDX_LOOP_C_84 : begin
        fsm_output = 9'b001010110;
        state_var_NS = IDX_LOOP_C_85;
      end
      IDX_LOOP_C_85 : begin
        fsm_output = 9'b001010111;
        state_var_NS = IDX_LOOP_C_86;
      end
      IDX_LOOP_C_86 : begin
        fsm_output = 9'b001011000;
        state_var_NS = IDX_LOOP_C_87;
      end
      IDX_LOOP_C_87 : begin
        fsm_output = 9'b001011001;
        state_var_NS = IDX_LOOP_C_88;
      end
      IDX_LOOP_C_88 : begin
        fsm_output = 9'b001011010;
        state_var_NS = IDX_LOOP_C_89;
      end
      IDX_LOOP_C_89 : begin
        fsm_output = 9'b001011011;
        state_var_NS = IDX_LOOP_C_90;
      end
      IDX_LOOP_C_90 : begin
        fsm_output = 9'b001011100;
        state_var_NS = IDX_LOOP_C_91;
      end
      IDX_LOOP_C_91 : begin
        fsm_output = 9'b001011101;
        state_var_NS = IDX_LOOP_C_92;
      end
      IDX_LOOP_C_92 : begin
        fsm_output = 9'b001011110;
        state_var_NS = IDX_LOOP_C_93;
      end
      IDX_LOOP_C_93 : begin
        fsm_output = 9'b001011111;
        state_var_NS = IDX_LOOP_C_94;
      end
      IDX_LOOP_C_94 : begin
        fsm_output = 9'b001100000;
        state_var_NS = IDX_LOOP_C_95;
      end
      IDX_LOOP_C_95 : begin
        fsm_output = 9'b001100001;
        state_var_NS = IDX_LOOP_C_96;
      end
      IDX_LOOP_C_96 : begin
        fsm_output = 9'b001100010;
        state_var_NS = IDX_LOOP_C_97;
      end
      IDX_LOOP_C_97 : begin
        fsm_output = 9'b001100011;
        if ( IDX_LOOP_C_97_tr0 ) begin
          state_var_NS = GROUP_LOOP_C_0;
        end
        else begin
          state_var_NS = IDX_LOOP_C_98;
        end
      end
      IDX_LOOP_C_98 : begin
        fsm_output = 9'b001100100;
        state_var_NS = IDX_LOOP_C_99;
      end
      IDX_LOOP_C_99 : begin
        fsm_output = 9'b001100101;
        state_var_NS = IDX_LOOP_C_100;
      end
      IDX_LOOP_C_100 : begin
        fsm_output = 9'b001100110;
        state_var_NS = IDX_LOOP_C_101;
      end
      IDX_LOOP_C_101 : begin
        fsm_output = 9'b001100111;
        state_var_NS = IDX_LOOP_C_102;
      end
      IDX_LOOP_C_102 : begin
        fsm_output = 9'b001101000;
        state_var_NS = IDX_LOOP_C_103;
      end
      IDX_LOOP_C_103 : begin
        fsm_output = 9'b001101001;
        state_var_NS = IDX_LOOP_C_104;
      end
      IDX_LOOP_C_104 : begin
        fsm_output = 9'b001101010;
        state_var_NS = IDX_LOOP_C_105;
      end
      IDX_LOOP_C_105 : begin
        fsm_output = 9'b001101011;
        state_var_NS = IDX_LOOP_C_106;
      end
      IDX_LOOP_C_106 : begin
        fsm_output = 9'b001101100;
        state_var_NS = IDX_LOOP_C_107;
      end
      IDX_LOOP_C_107 : begin
        fsm_output = 9'b001101101;
        state_var_NS = IDX_LOOP_C_108;
      end
      IDX_LOOP_C_108 : begin
        fsm_output = 9'b001101110;
        state_var_NS = IDX_LOOP_C_109;
      end
      IDX_LOOP_C_109 : begin
        fsm_output = 9'b001101111;
        state_var_NS = IDX_LOOP_C_110;
      end
      IDX_LOOP_C_110 : begin
        fsm_output = 9'b001110000;
        state_var_NS = IDX_LOOP_C_111;
      end
      IDX_LOOP_C_111 : begin
        fsm_output = 9'b001110001;
        state_var_NS = IDX_LOOP_C_112;
      end
      IDX_LOOP_C_112 : begin
        fsm_output = 9'b001110010;
        state_var_NS = IDX_LOOP_C_113;
      end
      IDX_LOOP_C_113 : begin
        fsm_output = 9'b001110011;
        state_var_NS = IDX_LOOP_C_114;
      end
      IDX_LOOP_C_114 : begin
        fsm_output = 9'b001110100;
        state_var_NS = IDX_LOOP_C_115;
      end
      IDX_LOOP_C_115 : begin
        fsm_output = 9'b001110101;
        state_var_NS = IDX_LOOP_C_116;
      end
      IDX_LOOP_C_116 : begin
        fsm_output = 9'b001110110;
        state_var_NS = IDX_LOOP_C_117;
      end
      IDX_LOOP_C_117 : begin
        fsm_output = 9'b001110111;
        state_var_NS = IDX_LOOP_C_118;
      end
      IDX_LOOP_C_118 : begin
        fsm_output = 9'b001111000;
        state_var_NS = IDX_LOOP_C_119;
      end
      IDX_LOOP_C_119 : begin
        fsm_output = 9'b001111001;
        state_var_NS = IDX_LOOP_C_120;
      end
      IDX_LOOP_C_120 : begin
        fsm_output = 9'b001111010;
        state_var_NS = IDX_LOOP_C_121;
      end
      IDX_LOOP_C_121 : begin
        fsm_output = 9'b001111011;
        state_var_NS = IDX_LOOP_C_122;
      end
      IDX_LOOP_C_122 : begin
        fsm_output = 9'b001111100;
        state_var_NS = IDX_LOOP_C_123;
      end
      IDX_LOOP_C_123 : begin
        fsm_output = 9'b001111101;
        state_var_NS = IDX_LOOP_C_124;
      end
      IDX_LOOP_C_124 : begin
        fsm_output = 9'b001111110;
        state_var_NS = IDX_LOOP_C_125;
      end
      IDX_LOOP_C_125 : begin
        fsm_output = 9'b001111111;
        state_var_NS = IDX_LOOP_C_126;
      end
      IDX_LOOP_C_126 : begin
        fsm_output = 9'b010000000;
        state_var_NS = IDX_LOOP_C_127;
      end
      IDX_LOOP_C_127 : begin
        fsm_output = 9'b010000001;
        state_var_NS = IDX_LOOP_C_128;
      end
      IDX_LOOP_C_128 : begin
        fsm_output = 9'b010000010;
        state_var_NS = IDX_LOOP_C_129;
      end
      IDX_LOOP_C_129 : begin
        fsm_output = 9'b010000011;
        if ( IDX_LOOP_C_129_tr0 ) begin
          state_var_NS = GROUP_LOOP_C_0;
        end
        else begin
          state_var_NS = IDX_LOOP_C_130;
        end
      end
      IDX_LOOP_C_130 : begin
        fsm_output = 9'b010000100;
        state_var_NS = IDX_LOOP_C_131;
      end
      IDX_LOOP_C_131 : begin
        fsm_output = 9'b010000101;
        state_var_NS = IDX_LOOP_C_132;
      end
      IDX_LOOP_C_132 : begin
        fsm_output = 9'b010000110;
        state_var_NS = IDX_LOOP_C_133;
      end
      IDX_LOOP_C_133 : begin
        fsm_output = 9'b010000111;
        state_var_NS = IDX_LOOP_C_134;
      end
      IDX_LOOP_C_134 : begin
        fsm_output = 9'b010001000;
        state_var_NS = IDX_LOOP_C_135;
      end
      IDX_LOOP_C_135 : begin
        fsm_output = 9'b010001001;
        state_var_NS = IDX_LOOP_C_136;
      end
      IDX_LOOP_C_136 : begin
        fsm_output = 9'b010001010;
        state_var_NS = IDX_LOOP_C_137;
      end
      IDX_LOOP_C_137 : begin
        fsm_output = 9'b010001011;
        state_var_NS = IDX_LOOP_C_138;
      end
      IDX_LOOP_C_138 : begin
        fsm_output = 9'b010001100;
        state_var_NS = IDX_LOOP_C_139;
      end
      IDX_LOOP_C_139 : begin
        fsm_output = 9'b010001101;
        state_var_NS = IDX_LOOP_C_140;
      end
      IDX_LOOP_C_140 : begin
        fsm_output = 9'b010001110;
        state_var_NS = IDX_LOOP_C_141;
      end
      IDX_LOOP_C_141 : begin
        fsm_output = 9'b010001111;
        state_var_NS = IDX_LOOP_C_142;
      end
      IDX_LOOP_C_142 : begin
        fsm_output = 9'b010010000;
        state_var_NS = IDX_LOOP_C_143;
      end
      IDX_LOOP_C_143 : begin
        fsm_output = 9'b010010001;
        state_var_NS = IDX_LOOP_C_144;
      end
      IDX_LOOP_C_144 : begin
        fsm_output = 9'b010010010;
        state_var_NS = IDX_LOOP_C_145;
      end
      IDX_LOOP_C_145 : begin
        fsm_output = 9'b010010011;
        state_var_NS = IDX_LOOP_C_146;
      end
      IDX_LOOP_C_146 : begin
        fsm_output = 9'b010010100;
        state_var_NS = IDX_LOOP_C_147;
      end
      IDX_LOOP_C_147 : begin
        fsm_output = 9'b010010101;
        state_var_NS = IDX_LOOP_C_148;
      end
      IDX_LOOP_C_148 : begin
        fsm_output = 9'b010010110;
        state_var_NS = IDX_LOOP_C_149;
      end
      IDX_LOOP_C_149 : begin
        fsm_output = 9'b010010111;
        state_var_NS = IDX_LOOP_C_150;
      end
      IDX_LOOP_C_150 : begin
        fsm_output = 9'b010011000;
        state_var_NS = IDX_LOOP_C_151;
      end
      IDX_LOOP_C_151 : begin
        fsm_output = 9'b010011001;
        state_var_NS = IDX_LOOP_C_152;
      end
      IDX_LOOP_C_152 : begin
        fsm_output = 9'b010011010;
        state_var_NS = IDX_LOOP_C_153;
      end
      IDX_LOOP_C_153 : begin
        fsm_output = 9'b010011011;
        state_var_NS = IDX_LOOP_C_154;
      end
      IDX_LOOP_C_154 : begin
        fsm_output = 9'b010011100;
        state_var_NS = IDX_LOOP_C_155;
      end
      IDX_LOOP_C_155 : begin
        fsm_output = 9'b010011101;
        state_var_NS = IDX_LOOP_C_156;
      end
      IDX_LOOP_C_156 : begin
        fsm_output = 9'b010011110;
        state_var_NS = IDX_LOOP_C_157;
      end
      IDX_LOOP_C_157 : begin
        fsm_output = 9'b010011111;
        state_var_NS = IDX_LOOP_C_158;
      end
      IDX_LOOP_C_158 : begin
        fsm_output = 9'b010100000;
        state_var_NS = IDX_LOOP_C_159;
      end
      IDX_LOOP_C_159 : begin
        fsm_output = 9'b010100001;
        state_var_NS = IDX_LOOP_C_160;
      end
      IDX_LOOP_C_160 : begin
        fsm_output = 9'b010100010;
        state_var_NS = IDX_LOOP_C_161;
      end
      IDX_LOOP_C_161 : begin
        fsm_output = 9'b010100011;
        if ( IDX_LOOP_C_161_tr0 ) begin
          state_var_NS = GROUP_LOOP_C_0;
        end
        else begin
          state_var_NS = IDX_LOOP_C_162;
        end
      end
      IDX_LOOP_C_162 : begin
        fsm_output = 9'b010100100;
        state_var_NS = IDX_LOOP_C_163;
      end
      IDX_LOOP_C_163 : begin
        fsm_output = 9'b010100101;
        state_var_NS = IDX_LOOP_C_164;
      end
      IDX_LOOP_C_164 : begin
        fsm_output = 9'b010100110;
        state_var_NS = IDX_LOOP_C_165;
      end
      IDX_LOOP_C_165 : begin
        fsm_output = 9'b010100111;
        state_var_NS = IDX_LOOP_C_166;
      end
      IDX_LOOP_C_166 : begin
        fsm_output = 9'b010101000;
        state_var_NS = IDX_LOOP_C_167;
      end
      IDX_LOOP_C_167 : begin
        fsm_output = 9'b010101001;
        state_var_NS = IDX_LOOP_C_168;
      end
      IDX_LOOP_C_168 : begin
        fsm_output = 9'b010101010;
        state_var_NS = IDX_LOOP_C_169;
      end
      IDX_LOOP_C_169 : begin
        fsm_output = 9'b010101011;
        state_var_NS = IDX_LOOP_C_170;
      end
      IDX_LOOP_C_170 : begin
        fsm_output = 9'b010101100;
        state_var_NS = IDX_LOOP_C_171;
      end
      IDX_LOOP_C_171 : begin
        fsm_output = 9'b010101101;
        state_var_NS = IDX_LOOP_C_172;
      end
      IDX_LOOP_C_172 : begin
        fsm_output = 9'b010101110;
        state_var_NS = IDX_LOOP_C_173;
      end
      IDX_LOOP_C_173 : begin
        fsm_output = 9'b010101111;
        state_var_NS = IDX_LOOP_C_174;
      end
      IDX_LOOP_C_174 : begin
        fsm_output = 9'b010110000;
        state_var_NS = IDX_LOOP_C_175;
      end
      IDX_LOOP_C_175 : begin
        fsm_output = 9'b010110001;
        state_var_NS = IDX_LOOP_C_176;
      end
      IDX_LOOP_C_176 : begin
        fsm_output = 9'b010110010;
        state_var_NS = IDX_LOOP_C_177;
      end
      IDX_LOOP_C_177 : begin
        fsm_output = 9'b010110011;
        state_var_NS = IDX_LOOP_C_178;
      end
      IDX_LOOP_C_178 : begin
        fsm_output = 9'b010110100;
        state_var_NS = IDX_LOOP_C_179;
      end
      IDX_LOOP_C_179 : begin
        fsm_output = 9'b010110101;
        state_var_NS = IDX_LOOP_C_180;
      end
      IDX_LOOP_C_180 : begin
        fsm_output = 9'b010110110;
        state_var_NS = IDX_LOOP_C_181;
      end
      IDX_LOOP_C_181 : begin
        fsm_output = 9'b010110111;
        state_var_NS = IDX_LOOP_C_182;
      end
      IDX_LOOP_C_182 : begin
        fsm_output = 9'b010111000;
        state_var_NS = IDX_LOOP_C_183;
      end
      IDX_LOOP_C_183 : begin
        fsm_output = 9'b010111001;
        state_var_NS = IDX_LOOP_C_184;
      end
      IDX_LOOP_C_184 : begin
        fsm_output = 9'b010111010;
        state_var_NS = IDX_LOOP_C_185;
      end
      IDX_LOOP_C_185 : begin
        fsm_output = 9'b010111011;
        state_var_NS = IDX_LOOP_C_186;
      end
      IDX_LOOP_C_186 : begin
        fsm_output = 9'b010111100;
        state_var_NS = IDX_LOOP_C_187;
      end
      IDX_LOOP_C_187 : begin
        fsm_output = 9'b010111101;
        state_var_NS = IDX_LOOP_C_188;
      end
      IDX_LOOP_C_188 : begin
        fsm_output = 9'b010111110;
        state_var_NS = IDX_LOOP_C_189;
      end
      IDX_LOOP_C_189 : begin
        fsm_output = 9'b010111111;
        state_var_NS = IDX_LOOP_C_190;
      end
      IDX_LOOP_C_190 : begin
        fsm_output = 9'b011000000;
        state_var_NS = IDX_LOOP_C_191;
      end
      IDX_LOOP_C_191 : begin
        fsm_output = 9'b011000001;
        state_var_NS = IDX_LOOP_C_192;
      end
      IDX_LOOP_C_192 : begin
        fsm_output = 9'b011000010;
        state_var_NS = IDX_LOOP_C_193;
      end
      IDX_LOOP_C_193 : begin
        fsm_output = 9'b011000011;
        if ( IDX_LOOP_C_193_tr0 ) begin
          state_var_NS = GROUP_LOOP_C_0;
        end
        else begin
          state_var_NS = IDX_LOOP_C_194;
        end
      end
      IDX_LOOP_C_194 : begin
        fsm_output = 9'b011000100;
        state_var_NS = IDX_LOOP_C_195;
      end
      IDX_LOOP_C_195 : begin
        fsm_output = 9'b011000101;
        state_var_NS = IDX_LOOP_C_196;
      end
      IDX_LOOP_C_196 : begin
        fsm_output = 9'b011000110;
        state_var_NS = IDX_LOOP_C_197;
      end
      IDX_LOOP_C_197 : begin
        fsm_output = 9'b011000111;
        state_var_NS = IDX_LOOP_C_198;
      end
      IDX_LOOP_C_198 : begin
        fsm_output = 9'b011001000;
        state_var_NS = IDX_LOOP_C_199;
      end
      IDX_LOOP_C_199 : begin
        fsm_output = 9'b011001001;
        state_var_NS = IDX_LOOP_C_200;
      end
      IDX_LOOP_C_200 : begin
        fsm_output = 9'b011001010;
        state_var_NS = IDX_LOOP_C_201;
      end
      IDX_LOOP_C_201 : begin
        fsm_output = 9'b011001011;
        state_var_NS = IDX_LOOP_C_202;
      end
      IDX_LOOP_C_202 : begin
        fsm_output = 9'b011001100;
        state_var_NS = IDX_LOOP_C_203;
      end
      IDX_LOOP_C_203 : begin
        fsm_output = 9'b011001101;
        state_var_NS = IDX_LOOP_C_204;
      end
      IDX_LOOP_C_204 : begin
        fsm_output = 9'b011001110;
        state_var_NS = IDX_LOOP_C_205;
      end
      IDX_LOOP_C_205 : begin
        fsm_output = 9'b011001111;
        state_var_NS = IDX_LOOP_C_206;
      end
      IDX_LOOP_C_206 : begin
        fsm_output = 9'b011010000;
        state_var_NS = IDX_LOOP_C_207;
      end
      IDX_LOOP_C_207 : begin
        fsm_output = 9'b011010001;
        state_var_NS = IDX_LOOP_C_208;
      end
      IDX_LOOP_C_208 : begin
        fsm_output = 9'b011010010;
        state_var_NS = IDX_LOOP_C_209;
      end
      IDX_LOOP_C_209 : begin
        fsm_output = 9'b011010011;
        state_var_NS = IDX_LOOP_C_210;
      end
      IDX_LOOP_C_210 : begin
        fsm_output = 9'b011010100;
        state_var_NS = IDX_LOOP_C_211;
      end
      IDX_LOOP_C_211 : begin
        fsm_output = 9'b011010101;
        state_var_NS = IDX_LOOP_C_212;
      end
      IDX_LOOP_C_212 : begin
        fsm_output = 9'b011010110;
        state_var_NS = IDX_LOOP_C_213;
      end
      IDX_LOOP_C_213 : begin
        fsm_output = 9'b011010111;
        state_var_NS = IDX_LOOP_C_214;
      end
      IDX_LOOP_C_214 : begin
        fsm_output = 9'b011011000;
        state_var_NS = IDX_LOOP_C_215;
      end
      IDX_LOOP_C_215 : begin
        fsm_output = 9'b011011001;
        state_var_NS = IDX_LOOP_C_216;
      end
      IDX_LOOP_C_216 : begin
        fsm_output = 9'b011011010;
        state_var_NS = IDX_LOOP_C_217;
      end
      IDX_LOOP_C_217 : begin
        fsm_output = 9'b011011011;
        state_var_NS = IDX_LOOP_C_218;
      end
      IDX_LOOP_C_218 : begin
        fsm_output = 9'b011011100;
        state_var_NS = IDX_LOOP_C_219;
      end
      IDX_LOOP_C_219 : begin
        fsm_output = 9'b011011101;
        state_var_NS = IDX_LOOP_C_220;
      end
      IDX_LOOP_C_220 : begin
        fsm_output = 9'b011011110;
        state_var_NS = IDX_LOOP_C_221;
      end
      IDX_LOOP_C_221 : begin
        fsm_output = 9'b011011111;
        state_var_NS = IDX_LOOP_C_222;
      end
      IDX_LOOP_C_222 : begin
        fsm_output = 9'b011100000;
        state_var_NS = IDX_LOOP_C_223;
      end
      IDX_LOOP_C_223 : begin
        fsm_output = 9'b011100001;
        state_var_NS = IDX_LOOP_C_224;
      end
      IDX_LOOP_C_224 : begin
        fsm_output = 9'b011100010;
        state_var_NS = IDX_LOOP_C_225;
      end
      IDX_LOOP_C_225 : begin
        fsm_output = 9'b011100011;
        if ( IDX_LOOP_C_225_tr0 ) begin
          state_var_NS = GROUP_LOOP_C_0;
        end
        else begin
          state_var_NS = IDX_LOOP_C_226;
        end
      end
      IDX_LOOP_C_226 : begin
        fsm_output = 9'b011100100;
        state_var_NS = IDX_LOOP_C_227;
      end
      IDX_LOOP_C_227 : begin
        fsm_output = 9'b011100101;
        state_var_NS = IDX_LOOP_C_228;
      end
      IDX_LOOP_C_228 : begin
        fsm_output = 9'b011100110;
        state_var_NS = IDX_LOOP_C_229;
      end
      IDX_LOOP_C_229 : begin
        fsm_output = 9'b011100111;
        state_var_NS = IDX_LOOP_C_230;
      end
      IDX_LOOP_C_230 : begin
        fsm_output = 9'b011101000;
        state_var_NS = IDX_LOOP_C_231;
      end
      IDX_LOOP_C_231 : begin
        fsm_output = 9'b011101001;
        state_var_NS = IDX_LOOP_C_232;
      end
      IDX_LOOP_C_232 : begin
        fsm_output = 9'b011101010;
        state_var_NS = IDX_LOOP_C_233;
      end
      IDX_LOOP_C_233 : begin
        fsm_output = 9'b011101011;
        state_var_NS = IDX_LOOP_C_234;
      end
      IDX_LOOP_C_234 : begin
        fsm_output = 9'b011101100;
        state_var_NS = IDX_LOOP_C_235;
      end
      IDX_LOOP_C_235 : begin
        fsm_output = 9'b011101101;
        state_var_NS = IDX_LOOP_C_236;
      end
      IDX_LOOP_C_236 : begin
        fsm_output = 9'b011101110;
        state_var_NS = IDX_LOOP_C_237;
      end
      IDX_LOOP_C_237 : begin
        fsm_output = 9'b011101111;
        state_var_NS = IDX_LOOP_C_238;
      end
      IDX_LOOP_C_238 : begin
        fsm_output = 9'b011110000;
        state_var_NS = IDX_LOOP_C_239;
      end
      IDX_LOOP_C_239 : begin
        fsm_output = 9'b011110001;
        state_var_NS = IDX_LOOP_C_240;
      end
      IDX_LOOP_C_240 : begin
        fsm_output = 9'b011110010;
        state_var_NS = IDX_LOOP_C_241;
      end
      IDX_LOOP_C_241 : begin
        fsm_output = 9'b011110011;
        state_var_NS = IDX_LOOP_C_242;
      end
      IDX_LOOP_C_242 : begin
        fsm_output = 9'b011110100;
        state_var_NS = IDX_LOOP_C_243;
      end
      IDX_LOOP_C_243 : begin
        fsm_output = 9'b011110101;
        state_var_NS = IDX_LOOP_C_244;
      end
      IDX_LOOP_C_244 : begin
        fsm_output = 9'b011110110;
        state_var_NS = IDX_LOOP_C_245;
      end
      IDX_LOOP_C_245 : begin
        fsm_output = 9'b011110111;
        state_var_NS = IDX_LOOP_C_246;
      end
      IDX_LOOP_C_246 : begin
        fsm_output = 9'b011111000;
        state_var_NS = IDX_LOOP_C_247;
      end
      IDX_LOOP_C_247 : begin
        fsm_output = 9'b011111001;
        state_var_NS = IDX_LOOP_C_248;
      end
      IDX_LOOP_C_248 : begin
        fsm_output = 9'b011111010;
        state_var_NS = IDX_LOOP_C_249;
      end
      IDX_LOOP_C_249 : begin
        fsm_output = 9'b011111011;
        state_var_NS = IDX_LOOP_C_250;
      end
      IDX_LOOP_C_250 : begin
        fsm_output = 9'b011111100;
        state_var_NS = IDX_LOOP_C_251;
      end
      IDX_LOOP_C_251 : begin
        fsm_output = 9'b011111101;
        state_var_NS = IDX_LOOP_C_252;
      end
      IDX_LOOP_C_252 : begin
        fsm_output = 9'b011111110;
        state_var_NS = IDX_LOOP_C_253;
      end
      IDX_LOOP_C_253 : begin
        fsm_output = 9'b011111111;
        state_var_NS = IDX_LOOP_C_254;
      end
      IDX_LOOP_C_254 : begin
        fsm_output = 9'b100000000;
        state_var_NS = IDX_LOOP_C_255;
      end
      IDX_LOOP_C_255 : begin
        fsm_output = 9'b100000001;
        state_var_NS = IDX_LOOP_C_256;
      end
      IDX_LOOP_C_256 : begin
        fsm_output = 9'b100000010;
        state_var_NS = IDX_LOOP_C_257;
      end
      IDX_LOOP_C_257 : begin
        fsm_output = 9'b100000011;
        if ( IDX_LOOP_C_257_tr0 ) begin
          state_var_NS = GROUP_LOOP_C_0;
        end
        else begin
          state_var_NS = IDX_LOOP_C_0;
        end
      end
      GROUP_LOOP_C_0 : begin
        fsm_output = 9'b100000100;
        if ( GROUP_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_1;
        end
        else begin
          state_var_NS = IDX_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 9'b100000101;
        if ( STAGE_LOOP_C_1_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 9'b100000110;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 9'b000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_core_wait_dp
// ------------------------------------------------------------------


module DIT_RELOOP_core_wait_dp (
  ensig_cgo_iro, ensig_cgo, IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo;
  output IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_en = ensig_cgo | ensig_cgo_iro;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP_core
// ------------------------------------------------------------------


module DIT_RELOOP_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_triosy_lz, twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz, twiddle_rsc_triosy_0_2_lz, twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz, twiddle_rsc_triosy_0_5_lz, twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz, vec_rsc_0_0_i_radr_d, vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_radr_d,
      vec_rsc_0_1_i_q_d, vec_rsc_0_2_i_radr_d, vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_radr_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_radr_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_radr_d,
      vec_rsc_0_5_i_q_d, vec_rsc_0_6_i_radr_d, vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_radr_d,
      vec_rsc_0_7_i_q_d, twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d, twiddle_rsc_0_2_i_q_d,
      twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_5_i_q_d, twiddle_rsc_0_6_i_q_d,
      twiddle_rsc_0_7_i_q_d, vec_rsc_0_0_i_wadr_d_pff, vec_rsc_0_0_i_d_d_pff, vec_rsc_0_0_i_we_d_pff,
      vec_rsc_0_0_i_re_d_pff, vec_rsc_0_1_i_wadr_d_pff, vec_rsc_0_1_i_d_d_pff, vec_rsc_0_1_i_we_d_pff,
      vec_rsc_0_1_i_re_d_pff, vec_rsc_0_2_i_we_d_pff, vec_rsc_0_2_i_re_d_pff, vec_rsc_0_3_i_we_d_pff,
      vec_rsc_0_3_i_re_d_pff, vec_rsc_0_4_i_we_d_pff, vec_rsc_0_4_i_re_d_pff, vec_rsc_0_5_i_we_d_pff,
      vec_rsc_0_5_i_re_d_pff, vec_rsc_0_6_i_we_d_pff, vec_rsc_0_6_i_re_d_pff, vec_rsc_0_7_i_we_d_pff,
      vec_rsc_0_7_i_re_d_pff, twiddle_rsc_0_0_i_radr_d_pff, twiddle_rsc_0_0_i_re_d_pff,
      twiddle_rsc_0_1_i_re_d_pff, twiddle_rsc_0_2_i_re_d_pff, twiddle_rsc_0_3_i_re_d_pff,
      twiddle_rsc_0_4_i_re_d_pff, twiddle_rsc_0_5_i_re_d_pff, twiddle_rsc_0_6_i_re_d_pff,
      twiddle_rsc_0_7_i_re_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  output r_rsc_triosy_lz;
  output twiddle_rsc_triosy_0_0_lz;
  output twiddle_rsc_triosy_0_1_lz;
  output twiddle_rsc_triosy_0_2_lz;
  output twiddle_rsc_triosy_0_3_lz;
  output twiddle_rsc_triosy_0_4_lz;
  output twiddle_rsc_triosy_0_5_lz;
  output twiddle_rsc_triosy_0_6_lz;
  output twiddle_rsc_triosy_0_7_lz;
  output [6:0] vec_rsc_0_0_i_radr_d;
  input [63:0] vec_rsc_0_0_i_q_d;
  output [6:0] vec_rsc_0_1_i_radr_d;
  input [63:0] vec_rsc_0_1_i_q_d;
  output [6:0] vec_rsc_0_2_i_radr_d;
  input [63:0] vec_rsc_0_2_i_q_d;
  output [6:0] vec_rsc_0_3_i_radr_d;
  input [63:0] vec_rsc_0_3_i_q_d;
  output [6:0] vec_rsc_0_4_i_radr_d;
  input [63:0] vec_rsc_0_4_i_q_d;
  output [6:0] vec_rsc_0_5_i_radr_d;
  input [63:0] vec_rsc_0_5_i_q_d;
  output [6:0] vec_rsc_0_6_i_radr_d;
  input [63:0] vec_rsc_0_6_i_q_d;
  output [6:0] vec_rsc_0_7_i_radr_d;
  input [63:0] vec_rsc_0_7_i_q_d;
  input [63:0] twiddle_rsc_0_0_i_q_d;
  input [63:0] twiddle_rsc_0_1_i_q_d;
  input [63:0] twiddle_rsc_0_2_i_q_d;
  input [63:0] twiddle_rsc_0_3_i_q_d;
  input [63:0] twiddle_rsc_0_4_i_q_d;
  input [63:0] twiddle_rsc_0_5_i_q_d;
  input [63:0] twiddle_rsc_0_6_i_q_d;
  input [63:0] twiddle_rsc_0_7_i_q_d;
  output [6:0] vec_rsc_0_0_i_wadr_d_pff;
  output [63:0] vec_rsc_0_0_i_d_d_pff;
  output vec_rsc_0_0_i_we_d_pff;
  output vec_rsc_0_0_i_re_d_pff;
  output [6:0] vec_rsc_0_1_i_wadr_d_pff;
  output [63:0] vec_rsc_0_1_i_d_d_pff;
  output vec_rsc_0_1_i_we_d_pff;
  output vec_rsc_0_1_i_re_d_pff;
  output vec_rsc_0_2_i_we_d_pff;
  output vec_rsc_0_2_i_re_d_pff;
  output vec_rsc_0_3_i_we_d_pff;
  output vec_rsc_0_3_i_re_d_pff;
  output vec_rsc_0_4_i_we_d_pff;
  output vec_rsc_0_4_i_re_d_pff;
  output vec_rsc_0_5_i_we_d_pff;
  output vec_rsc_0_5_i_re_d_pff;
  output vec_rsc_0_6_i_we_d_pff;
  output vec_rsc_0_6_i_re_d_pff;
  output vec_rsc_0_7_i_we_d_pff;
  output vec_rsc_0_7_i_re_d_pff;
  output [6:0] twiddle_rsc_0_0_i_radr_d_pff;
  output twiddle_rsc_0_0_i_re_d_pff;
  output twiddle_rsc_0_1_i_re_d_pff;
  output twiddle_rsc_0_2_i_re_d_pff;
  output twiddle_rsc_0_3_i_re_d_pff;
  output twiddle_rsc_0_4_i_re_d_pff;
  output twiddle_rsc_0_5_i_re_d_pff;
  output twiddle_rsc_0_6_i_re_d_pff;
  output twiddle_rsc_0_7_i_re_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  reg [127:0] IDX_LOOP_1_IDX_LOOP_rem_1_cmp_a;
  wire [63:0] IDX_LOOP_1_IDX_LOOP_rem_1_cmp_z;
  wire [63:0] IDX_LOOP_1_modulo_dev_cmp_return_rsc_z;
  wire IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_en;
  wire [8:0] fsm_output;
  wire [8:0] IDX_LOOP_idx2_acc_tmp;
  wire [9:0] nl_IDX_LOOP_idx2_acc_tmp;
  wire and_dcpl;
  wire and_dcpl_1;
  wire or_tmp_2;
  wire or_tmp_3;
  wire or_tmp_4;
  wire and_dcpl_15;
  wire or_tmp_11;
  wire or_tmp_16;
  wire or_tmp_19;
  wire or_tmp_26;
  wire and_dcpl_55;
  wire and_dcpl_66;
  wire and_dcpl_93;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_113;
  wire and_dcpl_114;
  wire and_dcpl_116;
  wire and_dcpl_117;
  wire and_dcpl_119;
  wire and_dcpl_120;
  wire and_dcpl_122;
  wire and_dcpl_123;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire and_dcpl_134;
  wire and_dcpl_135;
  wire and_dcpl_138;
  wire and_dcpl_151;
  wire and_dcpl_153;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire not_tmp_162;
  wire not_tmp_164;
  wire and_dcpl_176;
  wire not_tmp_180;
  wire and_dcpl_179;
  wire and_dcpl_183;
  wire and_dcpl_184;
  wire and_dcpl_185;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_193;
  wire and_dcpl_194;
  wire and_dcpl_198;
  wire and_dcpl_200;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire or_dcpl_74;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire and_dcpl_210;
  wire and_dcpl_212;
  wire and_dcpl_214;
  wire and_dcpl_215;
  wire and_dcpl_216;
  wire or_dcpl_76;
  wire and_dcpl_217;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_222;
  wire and_dcpl_224;
  wire and_dcpl_225;
  wire and_dcpl_227;
  wire and_dcpl_228;
  wire and_dcpl_230;
  wire and_dcpl_232;
  wire and_dcpl_234;
  wire or_dcpl_79;
  wire and_dcpl_235;
  wire nor_tmp_55;
  wire or_tmp_248;
  wire and_dcpl_241;
  wire and_dcpl_247;
  wire and_dcpl_249;
  wire and_dcpl_251;
  wire and_dcpl_252;
  wire and_dcpl_254;
  wire and_dcpl_256;
  wire and_dcpl_259;
  wire and_dcpl_261;
  wire and_dcpl_263;
  wire and_dcpl_265;
  wire and_dcpl_267;
  wire and_dcpl_271;
  wire or_dcpl_81;
  wire and_dcpl_275;
  wire and_dcpl_277;
  wire or_dcpl_83;
  wire and_dcpl_279;
  wire or_dcpl_84;
  wire and_dcpl_282;
  wire and_dcpl_284;
  wire and_dcpl_286;
  wire or_dcpl_85;
  wire and_dcpl_288;
  wire and_dcpl_293;
  wire and_dcpl_299;
  wire and_dcpl_306;
  wire and_dcpl_311;
  wire or_dcpl_87;
  wire and_dcpl_313;
  wire and_dcpl_315;
  wire and_dcpl_317;
  wire and_dcpl_319;
  wire and_dcpl_322;
  wire or_dcpl_90;
  wire and_dcpl_324;
  wire or_tmp_395;
  wire and_dcpl_331;
  wire and_dcpl_342;
  wire and_dcpl_345;
  wire and_dcpl_348;
  wire and_tmp_7;
  wire or_dcpl_103;
  wire and_dcpl_367;
  wire and_dcpl_368;
  wire and_tmp_9;
  wire and_dcpl_374;
  wire and_tmp_10;
  wire and_dcpl_377;
  wire and_tmp_11;
  wire and_dcpl_380;
  wire or_tmp_502;
  wire and_dcpl_383;
  wire or_tmp_505;
  wire mux_tmp_457;
  wire and_dcpl_386;
  wire and_dcpl_387;
  wire mux_tmp_461;
  wire and_dcpl_388;
  wire not_tmp_290;
  wire and_dcpl_390;
  wire not_tmp_292;
  wire not_tmp_296;
  wire not_tmp_298;
  wire or_tmp_516;
  wire and_dcpl_404;
  wire and_dcpl_407;
  wire and_dcpl_408;
  wire and_dcpl_413;
  wire and_dcpl_416;
  wire and_dcpl_417;
  wire and_dcpl_419;
  wire and_tmp_14;
  wire and_dcpl_423;
  wire and_dcpl_430;
  reg IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm;
  wire [6:0] IDX_LOOP_idx1_acc_psp_8_sva_mx0w0;
  wire [7:0] nl_IDX_LOOP_idx1_acc_psp_8_sva_mx0w0;
  reg [9:0] STAGE_LOOP_op_rshift_psp_1_sva;
  wire IDX_LOOP_f1_equal_tmp_3_mx0w0;
  wire IDX_LOOP_f1_equal_tmp_2_mx0w0;
  wire IDX_LOOP_f1_equal_tmp_1_mx0w0;
  wire IDX_LOOP_f1_equal_tmp_mx0w0;
  reg [9:0] GROUP_LOOP_j_10_0_sva_9_0;
  reg IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm;
  wire [8:0] IDX_LOOP_idx1_acc_psp_3_sva_mx0w0;
  wire [9:0] nl_IDX_LOOP_idx1_acc_psp_3_sva_mx0w0;
  reg [6:0] IDX_LOOP_t_10_3_sva_6_0;
  reg IDX_LOOP_slc_IDX_LOOP_acc_8_itm;
  reg IDX_LOOP_f1_equal_tmp_2;
  reg IDX_LOOP_f1_equal_tmp;
  reg IDX_LOOP_f1_equal_tmp_1;
  reg IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm;
  reg IDX_LOOP_f1_equal_tmp_3;
  wire [7:0] IDX_LOOP_idx1_acc_2_psp_sva_mx0w0;
  wire [8:0] nl_IDX_LOOP_idx1_acc_2_psp_sva_mx0w0;
  reg IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm;
  reg IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm;
  wire [8:0] IDX_LOOP_idx1_acc_psp_7_sva_mx0w0;
  wire [9:0] nl_IDX_LOOP_idx1_acc_psp_7_sva_mx0w0;
  reg IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm;
  reg IDX_LOOP_1_slc_IDX_LOOP_acc_10_itm;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_90_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_97_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_104_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_34_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_41_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_48_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_160_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_153_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_146_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_216_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_209_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_202_itm;
  reg [9:0] IDX_LOOP_idx2_9_0_2_sva;
  reg [9:0] IDX_LOOP_idx2_9_0_4_sva;
  reg [9:0] IDX_LOOP_idx2_9_0_sva;
  reg [9:0] IDX_LOOP_idx2_9_0_6_sva;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_30_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_44_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_51_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_107_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_100_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_86_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_163_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_156_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_142_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_212_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_198_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_219_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_32_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_39_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_53_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_109_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_88_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_95_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_165_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_151_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_144_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_207_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_200_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_221_itm;
  reg IDX_LOOP_f1_and_94_itm;
  reg IDX_LOOP_f1_and_78_itm;
  reg IDX_LOOP_f1_and_86_itm;
  reg IDX_LOOP_f1_and_42_itm;
  reg IDX_LOOP_f1_and_50_itm;
  reg IDX_LOOP_f1_and_58_itm;
  reg IDX_LOOP_f1_and_114_itm;
  reg IDX_LOOP_f1_and_122_itm;
  reg IDX_LOOP_f1_and_130_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_nor_16_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_nor_24_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_nor_8_itm;
  reg [8:0] IDX_LOOP_idx2_acc_1_psp_sva;
  reg [8:0] IDX_LOOP_idx2_acc_2_psp_sva;
  reg [8:0] IDX_LOOP_idx2_acc_3_psp_sva;
  reg [8:0] IDX_LOOP_idx2_acc_psp_sva;
  reg [8:0] IDX_LOOP_idx1_acc_psp_7_sva;
  reg [7:0] IDX_LOOP_idx1_acc_2_psp_sva;
  reg [8:0] IDX_LOOP_idx1_acc_psp_3_sva;
  wire [9:0] IDX_LOOP_idx2_9_0_2_sva_mx0w0;
  wire [10:0] nl_IDX_LOOP_idx2_9_0_2_sva_mx0w0;
  wire [8:0] IDX_LOOP_idx2_acc_1_psp_sva_mx0w0;
  wire [9:0] nl_IDX_LOOP_idx2_acc_1_psp_sva_mx0w0;
  wire [9:0] IDX_LOOP_idx2_9_0_4_sva_mx0w0;
  wire [10:0] nl_IDX_LOOP_idx2_9_0_4_sva_mx0w0;
  wire [8:0] IDX_LOOP_idx2_acc_2_psp_sva_mx0w0;
  wire [9:0] nl_IDX_LOOP_idx2_acc_2_psp_sva_mx0w0;
  wire [9:0] IDX_LOOP_idx2_9_0_6_sva_mx0w0;
  wire [10:0] nl_IDX_LOOP_idx2_9_0_6_sva_mx0w0;
  wire [9:0] IDX_LOOP_idx2_9_0_sva_mx0w0;
  wire [10:0] nl_IDX_LOOP_idx2_9_0_sva_mx0w0;
  wire [8:0] IDX_LOOP_idx2_acc_3_psp_sva_mx0w0;
  wire [9:0] nl_IDX_LOOP_idx2_acc_3_psp_sva_mx0w0;
  reg [6:0] reg_IDX_LOOP_t_10_3_ftd_1;
  reg [1:0] reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7;
  reg [2:0] reg_IDX_LOOP_1_lshift_idiv_ftd_7;
  reg [63:0] reg_IDX_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse;
  reg reg_twiddle_rsc_triosy_0_0_obj_ld_cse;
  reg reg_ensig_cgo_cse;
  wire or_676_cse;
  wire or_680_cse;
  wire and_509_cse;
  reg [63:0] reg_cse;
  reg [63:0] reg_1_cse;
  reg [63:0] reg_2_cse;
  wire and_513_cse;
  wire or_200_cse;
  wire nand_44_cse;
  wire or_677_cse;
  wire and_481_cse;
  wire or_290_cse;
  wire or_288_cse;
  wire or_286_cse;
  wire mux_256_cse;
  wire nand_23_cse;
  wire or_362_cse;
  wire or_425_cse;
  wire or_439_cse;
  wire or_437_cse;
  wire or_435_cse;
  wire or_504_cse;
  wire IDX_LOOP_f2_IDX_LOOP_f2_nor_cse;
  wire or_520_cse;
  wire or_519_cse;
  wire or_517_cse;
  wire or_515_cse;
  wire or_44_cse;
  wire or_51_cse;
  wire or_40_cse;
  wire or_347_cse;
  wire mux_293_cse;
  wire mux_289_cse;
  wire mux_286_cse;
  wire and_448_cse;
  wire or_47_cse;
  wire or_90_cse;
  wire mux_180_cse;
  wire nor_302_rmff;
  reg [63:0] IDX_LOOP_modulo_dev_return_1_sva;
  reg [63:0] tmp_10_lpi_4_dfm;
  reg [6:0] IDX_LOOP_idx1_acc_psp_8_sva;
  reg [63:0] p_sva;
  wire [9:0] STAGE_LOOP_op_rshift_itm;
  wire and_dcpl_431;
  wire and_dcpl_436;
  wire and_dcpl_443;
  wire [10:0] z_out;
  wire and_dcpl_454;
  wire [7:0] z_out_1;
  wire [8:0] nl_z_out_1;
  wire and_dcpl_468;
  wire and_dcpl_469;
  wire and_dcpl_475;
  wire and_dcpl_476;
  wire and_dcpl_477;
  wire and_dcpl_479;
  wire and_dcpl_480;
  wire and_dcpl_482;
  wire and_dcpl_484;
  wire and_dcpl_491;
  wire and_dcpl_492;
  wire and_dcpl_493;
  wire and_dcpl_496;
  wire and_dcpl_498;
  wire and_dcpl_503;
  wire [63:0] z_out_4;
  wire and_dcpl_509;
  wire and_dcpl_533;
  wire [127:0] z_out_5;
  wire and_dcpl_536;
  wire and_dcpl_544;
  wire and_dcpl_547;
  wire and_dcpl_551;
  wire and_dcpl_553;
  wire and_dcpl_555;
  wire and_dcpl_557;
  wire and_dcpl_559;
  wire and_dcpl_561;
  wire and_dcpl_563;
  wire [9:0] z_out_6;
  wire and_dcpl_570;
  wire and_dcpl_571;
  wire and_dcpl_574;
  wire and_dcpl_577;
  wire and_dcpl_579;
  wire [63:0] z_out_7;
  wire and_dcpl_587;
  wire and_dcpl_591;
  wire and_dcpl_593;
  wire [63:0] z_out_8;
  wire and_dcpl_600;
  wire and_dcpl_601;
  wire and_dcpl_604;
  wire and_dcpl_607;
  wire and_dcpl_610;
  wire and_dcpl_612;
  wire and_dcpl_615;
  wire and_dcpl_618;
  wire and_dcpl_620;
  wire and_dcpl_622;
  reg [3:0] STAGE_LOOP_gp_acc_psp_sva;
  reg [9:0] STAGE_LOOP_gp_lshift_psp_sva;
  reg [63:0] tmp_11_sva_3;
  reg [63:0] tmp_11_sva_5;
  reg [63:0] tmp_11_sva_7;
  reg [63:0] tmp_11_sva_9;
  reg [63:0] tmp_11_sva_29;
  reg [127:0] IDX_LOOP_1_mul_mut;
  reg IDX_LOOP_f2_IDX_LOOP_f2_nor_4_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_33_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_37_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_40_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_46_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_47_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_54_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_55_itm;
  reg [63:0] IDX_LOOP_mux1h_1_itm;
  reg IDX_LOOP_f1_and_39_itm;
  reg IDX_LOOP_f1_and_41_itm;
  reg IDX_LOOP_f1_and_43_itm;
  reg IDX_LOOP_f1_and_47_itm;
  reg IDX_LOOP_f1_and_49_itm;
  reg IDX_LOOP_f1_and_51_itm;
  reg IDX_LOOP_f1_and_55_itm;
  reg IDX_LOOP_f1_and_57_itm;
  reg IDX_LOOP_f1_and_59_itm;
  reg IDX_LOOP_f1_and_63_itm;
  reg IDX_LOOP_f1_and_65_itm;
  reg IDX_LOOP_f1_and_66_itm;
  reg IDX_LOOP_f1_and_67_itm;
  reg [63:0] IDX_LOOP_mux1h_2_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_nor_12_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_89_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_93_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_96_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_102_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_103_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_110_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_111_itm;
  reg [63:0] IDX_LOOP_mux1h_3_itm;
  reg IDX_LOOP_f1_and_75_itm;
  reg IDX_LOOP_f1_and_77_itm;
  reg IDX_LOOP_f1_and_79_itm;
  reg IDX_LOOP_f1_and_83_itm;
  reg IDX_LOOP_f1_and_85_itm;
  reg IDX_LOOP_f1_and_87_itm;
  reg IDX_LOOP_f1_and_91_itm;
  reg IDX_LOOP_f1_and_93_itm;
  reg IDX_LOOP_f1_and_95_itm;
  reg IDX_LOOP_f1_and_99_itm;
  reg IDX_LOOP_f1_and_101_itm;
  reg IDX_LOOP_f1_and_102_itm;
  reg IDX_LOOP_f1_and_103_itm;
  reg IDX_LOOP_IDX_LOOP_nor_12_itm;
  reg [63:0] IDX_LOOP_mux1h_4_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_145_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_nor_21_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_149_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_152_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_158_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_159_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_166_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_167_itm;
  reg [63:0] IDX_LOOP_mux1h_5_itm;
  reg IDX_LOOP_f1_and_111_itm;
  reg IDX_LOOP_f1_and_113_itm;
  reg IDX_LOOP_f1_and_115_itm;
  reg IDX_LOOP_f1_and_119_itm;
  reg IDX_LOOP_f1_and_121_itm;
  reg IDX_LOOP_f1_and_123_itm;
  reg IDX_LOOP_f1_and_127_itm;
  reg IDX_LOOP_f1_and_129_itm;
  reg IDX_LOOP_f1_and_131_itm;
  reg IDX_LOOP_f1_and_135_itm;
  reg IDX_LOOP_f1_and_137_itm;
  reg IDX_LOOP_f1_and_138_itm;
  reg IDX_LOOP_f1_and_139_itm;
  reg IDX_LOOP_IDX_LOOP_and_104_itm;
  reg IDX_LOOP_IDX_LOOP_and_106_itm;
  reg IDX_LOOP_IDX_LOOP_and_107_itm;
  reg IDX_LOOP_IDX_LOOP_and_108_itm;
  reg [63:0] IDX_LOOP_mux1h_6_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_nor_28_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_201_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_205_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_208_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_214_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_222_itm;
  reg IDX_LOOP_f2_IDX_LOOP_f2_and_223_itm;
  reg [63:0] IDX_LOOP_mux1h_7_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [3:0] STAGE_LOOP_i_3_0_sva_2;
  wire [4:0] nl_STAGE_LOOP_i_3_0_sva_2;
  wire GROUP_LOOP_j_10_0_sva_9_0_mx0c0;
  wire IDX_LOOP_f2_nor_cse_1;
  wire IDX_LOOP_f2_nor_1_cse_1;
  wire IDX_LOOP_f2_nor_2_cse_1;
  wire [63:0] IDX_LOOP_mux1h_68_itm_mx0w0;
  wire IDX_LOOP_modulo_dev_return_1_sva_mx0c1;
  wire IDX_LOOP_f2_nor_12_cse_1;
  wire IDX_LOOP_f2_nor_13_cse_1;
  wire IDX_LOOP_f2_nor_14_cse_1;
  wire IDX_LOOP_f2_nor_24_cse_1;
  wire IDX_LOOP_f2_nor_25_cse_1;
  wire IDX_LOOP_f2_nor_26_cse_1;
  wire IDX_LOOP_f2_nor_36_cse_1;
  wire IDX_LOOP_f2_nor_37_cse_1;
  wire IDX_LOOP_f2_nor_38_cse_1;
  wire IDX_LOOP_f2_nor_48_cse_1;
  wire IDX_LOOP_f2_nor_49_cse_1;
  wire IDX_LOOP_f2_nor_50_cse_1;
  wire IDX_LOOP_f2_nor_60_cse_1;
  wire IDX_LOOP_f2_nor_61_cse_1;
  wire IDX_LOOP_f2_nor_62_cse_1;
  wire IDX_LOOP_f2_nor_72_cse_1;
  wire IDX_LOOP_f2_nor_73_cse_1;
  wire IDX_LOOP_f2_nor_74_cse_1;
  wire IDX_LOOP_f2_nor_84_cse_1;
  wire IDX_LOOP_f2_nor_85_cse_1;
  wire IDX_LOOP_f2_nor_86_cse_1;
  wire and_636_ssc;
  wire IDX_LOOP_f2_and_8_cse;
  wire IDX_LOOP_f2_and_10_cse;
  wire IDX_LOOP_f2_and_14_cse;
  wire IDX_LOOP_f2_and_9_cse;
  wire IDX_LOOP_f2_and_11_cse;
  wire IDX_LOOP_f2_and_15_cse;
  wire nor_175_cse;
  wire nor_183_cse;
  wire nor_191_cse;
  wire nor_199_cse;
  wire nor_207_cse;
  wire nor_215_cse;
  wire nor_223_cse;
  wire and_489_cse;
  wire nor_327_cse;
  wire nor_326_cse;
  wire IDX_LOOP_f1_or_69_cse;
  wire IDX_LOOP_f1_or_70_cse;
  wire or_tmp;
  wire or_tmp_545;
  wire STAGE_LOOP_acc_itm_4_1;
  wire z_out_2_10;
  wire xnor_cse;
  wire IDX_LOOP_f1_or_64_tmp;

  wire[0:0] mux_187_nl;
  wire[0:0] nor_230_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] or_199_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] or_203_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] or_202_nl;
  wire[0:0] or_201_nl;
  wire[0:0] GROUP_LOOP_j_not_1_nl;
  wire[0:0] or_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] or_690_nl;
  wire[0:0] or_691_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] or_697_nl;
  wire[0:0] mux_530_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] nor_300_nl;
  wire[10:0] IDX_LOOP_3_acc_nl;
  wire[11:0] nl_IDX_LOOP_3_acc_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] nor_251_nl;
  wire[8:0] IDX_LOOP_acc_nl;
  wire[9:0] nl_IDX_LOOP_acc_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] mux_473_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] or_35_nl;
  wire[10:0] IDX_LOOP_5_acc_nl;
  wire[11:0] nl_IDX_LOOP_5_acc_nl;
  wire[0:0] mux_476_nl;
  wire[0:0] mux_475_nl;
  wire[10:0] IDX_LOOP_6_acc_nl;
  wire[11:0] nl_IDX_LOOP_6_acc_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] nand_15_nl;
  wire[10:0] IDX_LOOP_7_acc_nl;
  wire[11:0] nl_IDX_LOOP_7_acc_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] mux_482_nl;
  wire[7:0] IDX_LOOP_acc_5_nl;
  wire[8:0] nl_IDX_LOOP_acc_5_nl;
  wire[0:0] IDX_LOOP_f1_and_11_nl;
  wire[0:0] IDX_LOOP_f1_and_101_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] IDX_LOOP_f1_and_13_nl;
  wire[0:0] IDX_LOOP_f1_and_102_nl;
  wire[0:0] IDX_LOOP_f1_and_14_nl;
  wire[0:0] IDX_LOOP_f1_and_103_nl;
  wire[0:0] IDX_LOOP_f1_and_15_nl;
  wire[0:0] IDX_LOOP_f1_and_111_nl;
  wire[0:0] and_169_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] IDX_LOOP_f1_and_19_nl;
  wire[0:0] IDX_LOOP_f1_and_113_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] IDX_LOOP_f1_and_21_nl;
  wire[0:0] IDX_LOOP_f1_and_114_nl;
  wire[0:0] IDX_LOOP_f1_and_22_nl;
  wire[0:0] IDX_LOOP_f1_and_115_nl;
  wire[0:0] IDX_LOOP_f1_and_23_nl;
  wire[0:0] IDX_LOOP_f1_and_119_nl;
  wire[0:0] IDX_LOOP_f1_and_27_nl;
  wire[0:0] IDX_LOOP_f1_and_122_nl;
  wire[0:0] and_164_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] IDX_LOOP_f1_and_29_nl;
  wire[0:0] IDX_LOOP_f1_and_127_nl;
  wire[0:0] IDX_LOOP_f1_and_3_nl;
  wire[0:0] IDX_LOOP_f1_and_129_nl;
  wire[0:0] and_166_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] IDX_LOOP_f1_and_30_nl;
  wire[0:0] IDX_LOOP_f1_and_130_nl;
  wire[0:0] mux_497_nl;
  wire[0:0] IDX_LOOP_f1_and_31_nl;
  wire[0:0] IDX_LOOP_f1_and_135_nl;
  wire[0:0] IDX_LOOP_f1_and_5_nl;
  wire[0:0] IDX_LOOP_f1_and_137_nl;
  wire[0:0] and_412_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] nor_117_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] IDX_LOOP_f1_and_6_nl;
  wire[0:0] IDX_LOOP_f1_and_138_nl;
  wire[0:0] IDX_LOOP_f1_and_7_nl;
  wire[0:0] IDX_LOOP_f1_and_139_nl;
  wire[0:0] IDX_LOOP_IDX_LOOP_and_2_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_215_nl;
  wire[0:0] and_416_nl;
  wire[0:0] mux_501_nl;
  wire[0:0] nor_116_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] IDX_LOOP_f1_and_51_nl;
  wire[0:0] mux_504_nl;
  wire[0:0] mux_509_nl;
  wire[0:0] nor_115_nl;
  wire[0:0] mux_508_nl;
  wire[0:0] or_633_nl;
  wire[0:0] mux_507_nl;
  wire[0:0] or_630_nl;
  wire[0:0] IDX_LOOP_f2_and_nl;
  wire[0:0] IDX_LOOP_f2_and_1_nl;
  wire[0:0] IDX_LOOP_f2_or_nl;
  wire[0:0] IDX_LOOP_f2_and_3_nl;
  wire[0:0] IDX_LOOP_f2_or_1_nl;
  wire[0:0] IDX_LOOP_f2_or_4_nl;
  wire[0:0] IDX_LOOP_f2_and_6_nl;
  wire[0:0] IDX_LOOP_f2_and_7_nl;
  wire[0:0] IDX_LOOP_f2_or_2_nl;
  wire[0:0] IDX_LOOP_f2_or_3_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] nor_114_nl;
  wire[0:0] IDX_LOOP_f1_and_208_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_201_nl;
  wire[0:0] IDX_LOOP_f1_and_209_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_202_nl;
  wire[0:0] IDX_LOOP_f1_and_210_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_203_nl;
  wire[0:0] IDX_LOOP_f1_and_211_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_204_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] nor_113_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] nor_260_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] or_657_nl;
  wire[0:0] and_521_nl;
  wire[0:0] IDX_LOOP_f2_or_5_nl;
  wire[0:0] IDX_LOOP_f2_or_6_nl;
  wire[0:0] IDX_LOOP_IDX_LOOP_and_126_nl;
  wire[0:0] IDX_LOOP_IDX_LOOP_and_128_nl;
  wire[0:0] IDX_LOOP_IDX_LOOP_and_130_nl;
  wire[4:0] STAGE_LOOP_acc_nl;
  wire[5:0] nl_STAGE_LOOP_acc_nl;
  wire[0:0] nor_236_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] and_375_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] mux_485_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] nand_14_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] mux_491_nl;
  wire[0:0] or_587_nl;
  wire[0:0] mux_503_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] mux_506_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] nor_112_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] and_359_nl;
  wire[0:0] and_360_nl;
  wire[0:0] and_361_nl;
  wire[0:0] and_362_nl;
  wire[0:0] and_363_nl;
  wire[0:0] and_364_nl;
  wire[0:0] and_247_nl;
  wire[0:0] and_248_nl;
  wire[0:0] and_249_nl;
  wire[0:0] and_250_nl;
  wire[0:0] and_246_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] and_453_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] nor_130_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] or_549_nl;
  wire[0:0] or_548_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] nor_131_nl;
  wire[0:0] nor_132_nl;
  wire[0:0] nor_133_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] or_544_nl;
  wire[0:0] or_542_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] or_541_nl;
  wire[0:0] or_540_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] or_539_nl;
  wire[0:0] or_538_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] or_537_nl;
  wire[0:0] or_536_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] nor_128_nl;
  wire[0:0] or_570_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] or_568_nl;
  wire[0:0] or_566_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] or_565_nl;
  wire[0:0] or_563_nl;
  wire[0:0] mux_440_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] or_561_nl;
  wire[0:0] or_559_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] or_558_nl;
  wire[0:0] or_556_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] or_554_nl;
  wire[0:0] or_552_nl;
  wire[0:0] and_345_nl;
  wire[0:0] and_347_nl;
  wire[0:0] and_348_nl;
  wire[0:0] and_350_nl;
  wire[0:0] and_351_nl;
  wire[0:0] and_353_nl;
  wire[0:0] and_354_nl;
  wire[0:0] and_356_nl;
  wire[0:0] and_190_nl;
  wire[0:0] and_193_nl;
  wire[0:0] and_196_nl;
  wire[0:0] and_199_nl;
  wire[0:0] and_186_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] nor_138_nl;
  wire[0:0] mux_410_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] or_512_nl;
  wire[0:0] or_510_nl;
  wire[0:0] or_509_nl;
  wire[0:0] nor_139_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] or_506_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] or_502_nl;
  wire[0:0] or_500_nl;
  wire[0:0] or_498_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] or_497_nl;
  wire[0:0] or_495_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] or_493_nl;
  wire[0:0] or_491_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] nand_10_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] nor_134_nl;
  wire[0:0] nor_135_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] nor_136_nl;
  wire[0:0] nor_137_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] and_343_nl;
  wire[0:0] or_522_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] and_454_nl;
  wire[0:0] nor_99_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] and_455_nl;
  wire[0:0] nor_97_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] and_456_nl;
  wire[0:0] nor_95_nl;
  wire[0:0] and_334_nl;
  wire[0:0] and_335_nl;
  wire[0:0] and_338_nl;
  wire[0:0] and_339_nl;
  wire[0:0] and_340_nl;
  wire[0:0] and_341_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] and_458_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] and_459_nl;
  wire[0:0] mux_380_nl;
  wire[0:0] nor_142_nl;
  wire[0:0] nor_143_nl;
  wire[0:0] mux_379_nl;
  wire[0:0] nor_144_nl;
  wire[0:0] nor_145_nl;
  wire[0:0] nor_146_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] or_465_nl;
  wire[0:0] or_463_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] or_462_nl;
  wire[0:0] or_461_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] or_460_nl;
  wire[0:0] or_459_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] or_458_nl;
  wire[0:0] or_457_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] nor_140_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] nor_94_nl;
  wire[0:0] or_485_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] or_483_nl;
  wire[0:0] nor_93_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] or_481_nl;
  wire[0:0] or_479_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] or_478_nl;
  wire[0:0] or_476_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] or_474_nl;
  wire[0:0] or_472_nl;
  wire[0:0] and_313_nl;
  wire[0:0] and_315_nl;
  wire[0:0] and_318_nl;
  wire[0:0] and_320_nl;
  wire[0:0] and_324_nl;
  wire[0:0] and_326_nl;
  wire[0:0] and_329_nl;
  wire[0:0] and_331_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] nor_151_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] or_432_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] or_430_nl;
  wire[0:0] nor_152_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] nand_16_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] or_423_nl;
  wire[0:0] or_422_nl;
  wire[0:0] or_420_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] or_419_nl;
  wire[0:0] or_418_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] or_416_nl;
  wire[0:0] or_415_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] nor_147_nl;
  wire[0:0] and_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] and_525_nl;
  wire[0:0] and_526_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] or_443_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] and_308_nl;
  wire[0:0] nor_90_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] and_460_nl;
  wire[0:0] nor_88_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] and_461_nl;
  wire[0:0] nor_86_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] and_462_nl;
  wire[0:0] nor_84_nl;
  wire[0:0] and_299_nl;
  wire[0:0] and_300_nl;
  wire[0:0] and_301_nl;
  wire[0:0] and_302_nl;
  wire[0:0] and_305_nl;
  wire[0:0] and_306_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] and_466_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] nor_155_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] or_391_nl;
  wire[0:0] or_390_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] nor_156_nl;
  wire[0:0] nor_157_nl;
  wire[0:0] nor_158_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] or_386_nl;
  wire[0:0] or_384_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] or_383_nl;
  wire[0:0] or_382_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] or_381_nl;
  wire[0:0] or_380_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] or_379_nl;
  wire[0:0] or_378_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] or_413_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] nor_153_nl;
  wire[0:0] or_409_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] and_463_nl;
  wire[0:0] nor_79_nl;
  wire[0:0] or_406_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] or_405_nl;
  wire[0:0] or_403_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] and_464_nl;
  wire[0:0] or_399_nl;
  wire[0:0] nor_77_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] or_398_nl;
  wire[0:0] and_465_nl;
  wire[0:0] nor_75_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] or_396_nl;
  wire[0:0] or_394_nl;
  wire[0:0] and_277_nl;
  wire[0:0] and_279_nl;
  wire[0:0] and_283_nl;
  wire[0:0] and_285_nl;
  wire[0:0] and_286_nl;
  wire[0:0] and_288_nl;
  wire[0:0] and_292_nl;
  wire[0:0] and_294_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] nor_163_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] or_354_nl;
  wire[0:0] or_353_nl;
  wire[0:0] or_352_nl;
  wire[0:0] nor_164_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] or_349_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] or_346_nl;
  wire[0:0] or_344_nl;
  wire[0:0] or_342_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] or_341_nl;
  wire[0:0] or_339_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] or_338_nl;
  wire[0:0] or_336_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] nand_4_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] nor_159_nl;
  wire[0:0] and_522_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] and_523_nl;
  wire[0:0] and_524_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] mux_317_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] and_273_nl;
  wire[0:0] or_364_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] or_361_nl;
  wire[0:0] and_467_nl;
  wire[0:0] nor_71_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] or_359_nl;
  wire[0:0] and_468_nl;
  wire[0:0] nor_69_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] or_357_nl;
  wire[0:0] and_469_nl;
  wire[0:0] nor_67_nl;
  wire[0:0] and_254_nl;
  wire[0:0] and_257_nl;
  wire[0:0] and_261_nl;
  wire[0:0] and_264_nl;
  wire[0:0] and_268_nl;
  wire[0:0] and_270_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] and_478_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] and_479_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] nor_167_nl;
  wire[0:0] nor_168_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] nor_169_nl;
  wire[0:0] nor_170_nl;
  wire[0:0] nor_171_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] nand_31_nl;
  wire[0:0] or_313_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] or_312_nl;
  wire[0:0] or_311_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] or_310_nl;
  wire[0:0] or_309_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] or_308_nl;
  wire[0:0] or_307_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] or_674_nl;
  wire[0:0] nor_165_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] and_471_nl;
  wire[0:0] and_472_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] and_473_nl;
  wire[0:0] and_474_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] and_475_nl;
  wire[0:0] and_476_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] nand_68_nl;
  wire[0:0] nand_69_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] nand_67_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] and_205_nl;
  wire[0:0] and_210_nl;
  wire[0:0] and_217_nl;
  wire[0:0] and_222_nl;
  wire[0:0] and_227_nl;
  wire[0:0] and_230_nl;
  wire[0:0] and_237_nl;
  wire[0:0] and_240_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] nor_172_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] nand_42_nl;
  wire[0:0] or_283_nl;
  wire[0:0] nor_173_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] nand_43_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] nand_45_nl;
  wire[0:0] or_280_nl;
  wire[0:0] or_278_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] nand_48_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] nand_49_nl;
  wire[0:0] nand_50_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] or_297_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] or_295_nl;
  wire[0:0] or_293_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] or_291_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] and_480_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] and_482_nl;
  wire[0:0] and_483_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] and_484_nl;
  wire[0:0] and_485_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] and_486_nl;
  wire[0:0] and_487_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] nor_174_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] nor_182_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] nor_186_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] nor_190_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] nor_194_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] nor_198_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] nor_206_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] and_520_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] nor_218_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] nor_222_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] and_519_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] and_488_nl;
  wire[0:0] mux_nl;
  wire[0:0] or_698_nl;
  wire[0:0] nand_71_nl;
  wire[11:0] acc_nl;
  wire[12:0] nl_acc_nl;
  wire[9:0] IDX_LOOP_mux_25_nl;
  wire[0:0] IDX_LOOP_IDX_LOOP_nand_1_nl;
  wire[6:0] IDX_LOOP_IDX_LOOP_and_132_nl;
  wire[0:0] not_1293_nl;
  wire[6:0] STAGE_LOOP_gp_mux_5_nl;
  wire[11:0] acc_2_nl;
  wire[12:0] nl_acc_2_nl;
  wire[10:0] IDX_LOOP_mux_26_nl;
  wire[9:0] IDX_LOOP_mux_27_nl;
  wire[63:0] IDX_LOOP_mux1h_102_nl;
  wire[0:0] and_719_nl;
  wire[0:0] and_720_nl;
  wire[0:0] and_721_nl;
  wire[0:0] and_722_nl;
  wire[0:0] and_723_nl;
  wire[0:0] and_724_nl;
  wire[0:0] and_725_nl;
  wire[63:0] IDX_LOOP_mux_28_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_205_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_206_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_207_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_208_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_209_nl;
  wire[0:0] IDX_LOOP_f1_or_82_nl;
  wire[0:0] IDX_LOOP_f1_or_83_nl;
  wire[0:0] IDX_LOOP_f1_or_84_nl;
  wire[0:0] IDX_LOOP_f1_or_85_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_210_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_224_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_225_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_226_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_227_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_211_nl;
  wire[0:0] IDX_LOOP_f1_or_86_nl;
  wire[0:0] IDX_LOOP_f1_or_87_nl;
  wire[0:0] IDX_LOOP_f1_or_88_nl;
  wire[0:0] IDX_LOOP_f1_or_89_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_212_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_213_nl;
  wire[0:0] IDX_LOOP_f1_or_90_nl;
  wire[0:0] IDX_LOOP_f1_or_91_nl;
  wire[0:0] IDX_LOOP_f1_or_92_nl;
  wire[0:0] IDX_LOOP_f1_or_93_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_214_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_215_nl;
  wire[0:0] IDX_LOOP_f1_or_94_nl;
  wire[0:0] IDX_LOOP_f1_or_95_nl;
  wire[0:0] IDX_LOOP_f1_or_96_nl;
  wire[0:0] IDX_LOOP_f1_or_97_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_216_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_217_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_260_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_261_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_262_nl;
  wire[0:0] IDX_LOOP_f2_IDX_LOOP_f2_and_263_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_218_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_219_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_220_nl;
  wire[0:0] IDX_LOOP_f1_or_98_nl;
  wire[0:0] IDX_LOOP_f1_or_99_nl;
  wire[0:0] IDX_LOOP_f1_or_100_nl;
  wire[0:0] IDX_LOOP_f1_or_101_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_221_nl;
  wire[0:0] IDX_LOOP_f1_or_102_nl;
  wire[0:0] IDX_LOOP_f1_or_103_nl;
  wire[0:0] IDX_LOOP_f1_or_104_nl;
  wire[0:0] IDX_LOOP_f1_or_105_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_222_nl;
  wire[0:0] IDX_LOOP_f1_or_106_nl;
  wire[0:0] IDX_LOOP_f1_or_107_nl;
  wire[0:0] IDX_LOOP_f1_or_108_nl;
  wire[0:0] IDX_LOOP_f1_or_109_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_223_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_224_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_225_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_226_nl;
  wire[0:0] IDX_LOOP_f1_and_160_nl;
  wire[0:0] IDX_LOOP_f1_and_161_nl;
  wire[0:0] IDX_LOOP_f1_and_162_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_227_nl;
  wire[0:0] IDX_LOOP_f1_or_110_nl;
  wire[0:0] IDX_LOOP_f1_or_111_nl;
  wire[0:0] IDX_LOOP_f1_or_112_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_228_nl;
  wire[0:0] IDX_LOOP_f1_or_113_nl;
  wire[0:0] IDX_LOOP_f1_or_114_nl;
  wire[0:0] IDX_LOOP_f1_or_115_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_229_nl;
  wire[0:0] IDX_LOOP_f1_or_116_nl;
  wire[0:0] IDX_LOOP_f1_or_117_nl;
  wire[0:0] IDX_LOOP_f1_or_118_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_230_nl;
  wire[0:0] IDX_LOOP_f1_or_119_nl;
  wire[0:0] IDX_LOOP_f1_or_120_nl;
  wire[0:0] IDX_LOOP_f1_or_121_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_231_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_232_nl;
  wire[0:0] IDX_LOOP_f1_or_122_nl;
  wire[0:0] IDX_LOOP_f1_or_123_nl;
  wire[0:0] IDX_LOOP_f1_or_124_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_233_nl;
  wire[0:0] IDX_LOOP_f1_and_187_nl;
  wire[0:0] IDX_LOOP_f1_and_188_nl;
  wire[0:0] IDX_LOOP_f1_and_189_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_234_nl;
  wire[0:0] IDX_LOOP_f1_and_190_nl;
  wire[0:0] IDX_LOOP_f1_and_191_nl;
  wire[0:0] IDX_LOOP_f1_and_192_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_235_nl;
  wire[0:0] IDX_LOOP_f1_or_125_nl;
  wire[0:0] IDX_LOOP_f1_or_126_nl;
  wire[0:0] IDX_LOOP_f1_or_127_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_236_nl;
  wire[0:0] IDX_LOOP_f1_or_128_nl;
  wire[0:0] IDX_LOOP_f1_or_129_nl;
  wire[0:0] IDX_LOOP_f1_or_130_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_237_nl;
  wire[0:0] IDX_LOOP_f1_or_131_nl;
  wire[0:0] IDX_LOOP_f1_or_132_nl;
  wire[0:0] IDX_LOOP_f1_or_133_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_238_nl;
  wire[0:0] IDX_LOOP_f1_and_205_nl;
  wire[0:0] IDX_LOOP_f1_and_206_nl;
  wire[0:0] IDX_LOOP_f1_and_207_nl;
  wire[0:0] IDX_LOOP_f1_mux1h_239_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[64:0] acc_3_nl;
  wire[65:0] nl_acc_3_nl;
  wire[63:0] IDX_LOOP_mux_29_nl;
  wire[0:0] IDX_LOOP_or_12_nl;
  wire[0:0] IDX_LOOP_or_13_nl;
  wire[63:0] IDX_LOOP_mux1h_103_nl;
  wire[0:0] IDX_LOOP_or_14_nl;
  wire[0:0] IDX_LOOP_or_15_nl;
  wire [63:0] nl_IDX_LOOP_1_modulo_dev_cmp_base_rsc_dat;
  assign IDX_LOOP_or_12_nl = and_dcpl_604 | and_dcpl_607 | and_dcpl_610 | and_dcpl_612
      | and_dcpl_615 | and_dcpl_618 | and_dcpl_620 | and_dcpl_622;
  assign IDX_LOOP_mux_29_nl = MUX_v_64_2_2(z_out_4, tmp_10_lpi_4_dfm, IDX_LOOP_or_12_nl);
  assign IDX_LOOP_or_13_nl = (~ and_dcpl_604) | and_dcpl_601 | and_dcpl_607 | and_dcpl_610
      | and_dcpl_612 | and_dcpl_615 | and_dcpl_618 | and_dcpl_620 | and_dcpl_622;
  assign IDX_LOOP_or_14_nl = and_dcpl_607 | and_dcpl_612 | and_dcpl_618 | and_dcpl_622;
  assign IDX_LOOP_or_15_nl = and_dcpl_610 | and_dcpl_615 | and_dcpl_620;
  assign IDX_LOOP_mux1h_103_nl = MUX1HOT_v_64_4_2((~ IDX_LOOP_modulo_dev_return_1_sva),
      IDX_LOOP_modulo_dev_return_1_sva, (~ z_out_7), (~ z_out_8), {and_dcpl_601 ,
      and_dcpl_604 , IDX_LOOP_or_14_nl , IDX_LOOP_or_15_nl});
  assign nl_acc_3_nl = ({IDX_LOOP_mux_29_nl , IDX_LOOP_or_13_nl}) + ({IDX_LOOP_mux1h_103_nl
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[64:0];
  assign nl_IDX_LOOP_1_modulo_dev_cmp_base_rsc_dat = readslicef_65_64_1(acc_3_nl);
  wire [63:0] nl_IDX_LOOP_1_modulo_dev_cmp_m_rsc_dat;
  assign nl_IDX_LOOP_1_modulo_dev_cmp_m_rsc_dat = p_sva;
  wire [0:0] nl_IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat;
  assign nl_IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat = and_dcpl_103 & (~
      (fsm_output[1])) & (~ (fsm_output[8]));
  wire[6:0] STAGE_LOOP_gp_and_nl;
  wire[0:0] STAGE_LOOP_gp_not_1_nl;
  wire[0:0] STAGE_LOOP_gp_STAGE_LOOP_gp_or_nl;
  wire[0:0] STAGE_LOOP_gp_STAGE_LOOP_gp_or_1_nl;
  wire[0:0] STAGE_LOOP_gp_STAGE_LOOP_gp_or_2_nl;
  wire [9:0] nl_IDX_LOOP_1_lshift_rg_a;
  assign STAGE_LOOP_gp_not_1_nl = ~ and_636_ssc;
  assign STAGE_LOOP_gp_and_nl = MUX_v_7_2_2(7'b0000000, IDX_LOOP_t_10_3_sva_6_0,
      STAGE_LOOP_gp_not_1_nl);
  assign STAGE_LOOP_gp_STAGE_LOOP_gp_or_nl = (~(and_636_ssc | and_dcpl_544 | and_dcpl_547
      | and_dcpl_551 | and_dcpl_553)) | and_dcpl_555 | and_dcpl_557 | and_dcpl_561
      | and_dcpl_563;
  assign STAGE_LOOP_gp_STAGE_LOOP_gp_or_1_nl = (~(and_636_ssc | and_dcpl_544 | and_dcpl_547
      | and_dcpl_555 | and_dcpl_557)) | and_dcpl_551 | and_dcpl_553 | and_dcpl_561
      | and_dcpl_563;
  assign STAGE_LOOP_gp_STAGE_LOOP_gp_or_2_nl = (~(and_dcpl_544 | and_dcpl_551 | and_dcpl_555
      | and_dcpl_561)) | and_636_ssc | and_dcpl_547 | and_dcpl_553 | and_dcpl_557
      | and_dcpl_563;
  assign nl_IDX_LOOP_1_lshift_rg_a = {STAGE_LOOP_gp_and_nl , STAGE_LOOP_gp_STAGE_LOOP_gp_or_nl
      , STAGE_LOOP_gp_STAGE_LOOP_gp_or_1_nl , STAGE_LOOP_gp_STAGE_LOOP_gp_or_2_nl};
  wire[0:0] STAGE_LOOP_gp_or_nl;
  wire [3:0] nl_IDX_LOOP_1_lshift_rg_s;
  assign STAGE_LOOP_gp_or_nl = and_dcpl_544 | and_dcpl_547 | and_dcpl_551 | and_dcpl_553
      | and_dcpl_555 | and_dcpl_557 | and_dcpl_561 | and_dcpl_563;
  assign nl_IDX_LOOP_1_lshift_rg_s = MUX_v_4_2_2((z_out_1[3:0]), STAGE_LOOP_gp_acc_psp_sva,
      STAGE_LOOP_gp_or_nl);
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_33_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_33_tr0 = ~ IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_65_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_65_tr0 = ~ IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_97_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_97_tr0 = ~ IDX_LOOP_slc_IDX_LOOP_acc_8_itm;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_129_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_129_tr0 = ~ IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_161_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_161_tr0 = ~ IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_193_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_193_tr0 = ~ IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_225_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_225_tr0 = ~ IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_257_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_257_tr0 = ~ IDX_LOOP_1_slc_IDX_LOOP_acc_10_itm;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_GROUP_LOOP_C_0_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_GROUP_LOOP_C_0_tr0 = ~ z_out_2_10;
  wire [0:0] nl_DIT_RELOOP_core_core_fsm_inst_STAGE_LOOP_C_1_tr0;
  assign nl_DIT_RELOOP_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 = STAGE_LOOP_acc_itm_4_1;
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_7_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_6_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_5_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_4_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_3_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_2_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_1_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_0_obj (
      .ld(reg_twiddle_rsc_triosy_0_0_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_0_lz)
    );
  mgc_rem #(.width_a(32'sd128),
  .width_b(32'sd64),
  .signd(32'sd0)) IDX_LOOP_1_IDX_LOOP_rem_1_cmp (
      .a(IDX_LOOP_1_IDX_LOOP_rem_1_cmp_a),
      .b(reg_IDX_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse),
      .z(IDX_LOOP_1_IDX_LOOP_rem_1_cmp_z)
    );
  modulo_dev  IDX_LOOP_1_modulo_dev_cmp (
      .base_rsc_dat(nl_IDX_LOOP_1_modulo_dev_cmp_base_rsc_dat[63:0]),
      .m_rsc_dat(nl_IDX_LOOP_1_modulo_dev_cmp_m_rsc_dat[63:0]),
      .return_rsc_z(IDX_LOOP_1_modulo_dev_cmp_return_rsc_z),
      .ccs_ccore_start_rsc_dat(nl_IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat[0:0]),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_en)
    );
  mgc_shift_r_v5 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_op_rshift_rg (
      .a(11'b10000000000),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_op_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd10),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) IDX_LOOP_1_lshift_rg (
      .a(nl_IDX_LOOP_1_lshift_rg_a[9:0]),
      .s(nl_IDX_LOOP_1_lshift_rg_s[3:0]),
      .z(z_out_6)
    );
  DIT_RELOOP_core_wait_dp DIT_RELOOP_core_wait_dp_inst (
      .ensig_cgo_iro(nor_302_rmff),
      .ensig_cgo(reg_ensig_cgo_cse),
      .IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_en(IDX_LOOP_1_modulo_dev_cmp_ccs_ccore_en)
    );
  DIT_RELOOP_core_core_fsm DIT_RELOOP_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .IDX_LOOP_C_33_tr0(nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_33_tr0[0:0]),
      .IDX_LOOP_C_65_tr0(nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_65_tr0[0:0]),
      .IDX_LOOP_C_97_tr0(nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_97_tr0[0:0]),
      .IDX_LOOP_C_129_tr0(nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_129_tr0[0:0]),
      .IDX_LOOP_C_161_tr0(nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_161_tr0[0:0]),
      .IDX_LOOP_C_193_tr0(nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_193_tr0[0:0]),
      .IDX_LOOP_C_225_tr0(nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_225_tr0[0:0]),
      .IDX_LOOP_C_257_tr0(nl_DIT_RELOOP_core_core_fsm_inst_IDX_LOOP_C_257_tr0[0:0]),
      .GROUP_LOOP_C_0_tr0(nl_DIT_RELOOP_core_core_fsm_inst_GROUP_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_1_tr0(nl_DIT_RELOOP_core_core_fsm_inst_STAGE_LOOP_C_1_tr0[0:0])
    );
  assign or_676_cse = (fsm_output[7:0]!=8'b00000000);
  assign mux_188_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[2]);
  assign or_199_nl = (fsm_output[3:2]!=2'b01);
  assign mux_189_nl = MUX_s_1_2_2(mux_188_nl, or_199_nl, or_680_cse);
  assign nor_302_rmff = ~(mux_189_nl | (fsm_output[4]) | (fsm_output[8]));
  assign or_200_cse = (fsm_output[2:0]!=3'b000);
  assign mux_293_cse = MUX_s_1_2_2((fsm_output[0]), nor_tmp_55, IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm);
  assign mux_289_cse = MUX_s_1_2_2((fsm_output[0]), nor_tmp_55, IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm);
  assign mux_286_cse = MUX_s_1_2_2((fsm_output[0]), nor_tmp_55, IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm);
  assign or_347_cse = (IDX_LOOP_idx2_9_0_2_sva[1]) | nand_23_cse;
  assign and_513_cse = (fsm_output[6:5]==2'b11);
  assign or_90_cse = (fsm_output[7:5]!=3'b000) | or_tmp_3;
  assign mux_493_nl = MUX_s_1_2_2(or_tmp_502, (~ mux_tmp_461), fsm_output[7]);
  assign IDX_LOOP_f1_or_69_cse = ~(mux_493_nl & (~ (fsm_output[8])));
  assign mux_494_nl = MUX_s_1_2_2(not_tmp_296, mux_tmp_461, fsm_output[7]);
  assign IDX_LOOP_f1_or_70_cse = mux_494_nl | (fsm_output[8]);
  assign or_680_cse = (fsm_output[1:0]!=2'b00);
  assign and_448_cse = or_680_cse & (fsm_output[2]);
  assign IDX_LOOP_f2_IDX_LOOP_f2_nor_cse = ~((IDX_LOOP_idx2_acc_tmp[1:0]!=2'b00)
      | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign and_509_cse = (fsm_output[1:0]==2'b11);
  assign IDX_LOOP_f2_and_8_cse = (~ (IDX_LOOP_idx2_acc_1_psp_sva[1])) & and_dcpl_207;
  assign IDX_LOOP_f2_and_10_cse = (IDX_LOOP_idx2_acc_2_psp_sva[0]) & and_dcpl_219;
  assign IDX_LOOP_f2_and_14_cse = (IDX_LOOP_idx2_acc_3_psp_sva[0]) & and_dcpl_227;
  assign IDX_LOOP_f2_and_9_cse = (IDX_LOOP_idx2_acc_1_psp_sva[1]) & and_dcpl_207;
  assign IDX_LOOP_f2_and_11_cse = (~ (IDX_LOOP_idx2_acc_2_psp_sva[0])) & and_dcpl_219;
  assign IDX_LOOP_f2_and_15_cse = (~ (IDX_LOOP_idx2_acc_3_psp_sva[0])) & and_dcpl_227;
  assign IDX_LOOP_f1_or_64_tmp = and_dcpl_247 | and_dcpl_254 | and_dcpl_261 | and_dcpl_267;
  assign xnor_cse = ~((fsm_output[5]) ^ (fsm_output[7]));
  assign nl_STAGE_LOOP_i_3_0_sva_2 = STAGE_LOOP_i_3_0_sva + 4'b0001;
  assign STAGE_LOOP_i_3_0_sva_2 = nl_STAGE_LOOP_i_3_0_sva_2[3:0];
  assign nl_IDX_LOOP_idx2_acc_tmp = ({IDX_LOOP_idx1_acc_psp_8_sva_mx0w0 , (z_out_5[1:0])})
      + (STAGE_LOOP_op_rshift_psp_1_sva[9:1]);
  assign IDX_LOOP_idx2_acc_tmp = nl_IDX_LOOP_idx2_acc_tmp[8:0];
  assign nl_IDX_LOOP_idx1_acc_psp_8_sva_mx0w0 = (z_out_5[8:2]) + IDX_LOOP_t_10_3_sva_6_0;
  assign IDX_LOOP_idx1_acc_psp_8_sva_mx0w0 = nl_IDX_LOOP_idx1_acc_psp_8_sva_mx0w0[6:0];
  assign nl_IDX_LOOP_idx2_9_0_2_sva_mx0w0 = ({IDX_LOOP_idx1_acc_psp_8_sva_mx0w0 ,
      (z_out_5[1:0]) , 1'b1}) + STAGE_LOOP_op_rshift_psp_1_sva;
  assign IDX_LOOP_idx2_9_0_2_sva_mx0w0 = nl_IDX_LOOP_idx2_9_0_2_sva_mx0w0[9:0];
  assign IDX_LOOP_f1_equal_tmp_mx0w0 = ~((z_out_5[1:0]!=2'b00));
  assign IDX_LOOP_f1_equal_tmp_1_mx0w0 = (z_out_5[1:0]==2'b01);
  assign IDX_LOOP_f1_equal_tmp_2_mx0w0 = (z_out_5[1:0]==2'b10);
  assign IDX_LOOP_f1_equal_tmp_3_mx0w0 = (z_out_5[1:0]==2'b11);
  assign nl_IDX_LOOP_idx2_acc_1_psp_sva_mx0w0 = IDX_LOOP_idx1_acc_psp_3_sva_mx0w0
      + (STAGE_LOOP_op_rshift_psp_1_sva[9:1]);
  assign IDX_LOOP_idx2_acc_1_psp_sva_mx0w0 = nl_IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[8:0];
  assign nl_IDX_LOOP_idx1_acc_psp_3_sva_mx0w0 = (z_out_5[8:0]) + ({IDX_LOOP_t_10_3_sva_6_0
      , 2'b01});
  assign IDX_LOOP_idx1_acc_psp_3_sva_mx0w0 = nl_IDX_LOOP_idx1_acc_psp_3_sva_mx0w0[8:0];
  assign nl_IDX_LOOP_idx2_9_0_4_sva_mx0w0 = ({IDX_LOOP_idx1_acc_psp_3_sva_mx0w0 ,
      1'b1}) + STAGE_LOOP_op_rshift_psp_1_sva;
  assign IDX_LOOP_idx2_9_0_4_sva_mx0w0 = nl_IDX_LOOP_idx2_9_0_4_sva_mx0w0[9:0];
  assign nl_IDX_LOOP_idx2_acc_2_psp_sva_mx0w0 = ({IDX_LOOP_idx1_acc_2_psp_sva_mx0w0
      , (z_out_5[0])}) + (STAGE_LOOP_op_rshift_psp_1_sva[9:1]);
  assign IDX_LOOP_idx2_acc_2_psp_sva_mx0w0 = nl_IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[8:0];
  assign nl_IDX_LOOP_idx1_acc_2_psp_sva_mx0w0 = (z_out_5[8:1]) + ({IDX_LOOP_t_10_3_sva_6_0
      , 1'b1});
  assign IDX_LOOP_idx1_acc_2_psp_sva_mx0w0 = nl_IDX_LOOP_idx1_acc_2_psp_sva_mx0w0[7:0];
  assign nl_IDX_LOOP_idx2_9_0_6_sva_mx0w0 = ({IDX_LOOP_idx1_acc_2_psp_sva_mx0w0 ,
      (z_out_5[0]) , 1'b1}) + STAGE_LOOP_op_rshift_psp_1_sva;
  assign IDX_LOOP_idx2_9_0_6_sva_mx0w0 = nl_IDX_LOOP_idx2_9_0_6_sva_mx0w0[9:0];
  assign nl_IDX_LOOP_idx2_acc_3_psp_sva_mx0w0 = IDX_LOOP_idx1_acc_psp_7_sva_mx0w0
      + (STAGE_LOOP_op_rshift_psp_1_sva[9:1]);
  assign IDX_LOOP_idx2_acc_3_psp_sva_mx0w0 = nl_IDX_LOOP_idx2_acc_3_psp_sva_mx0w0[8:0];
  assign nl_IDX_LOOP_idx1_acc_psp_7_sva_mx0w0 = (z_out_5[8:0]) + ({IDX_LOOP_t_10_3_sva_6_0
      , 2'b11});
  assign IDX_LOOP_idx1_acc_psp_7_sva_mx0w0 = nl_IDX_LOOP_idx1_acc_psp_7_sva_mx0w0[8:0];
  assign nl_IDX_LOOP_idx2_9_0_sva_mx0w0 = ({IDX_LOOP_idx1_acc_psp_7_sva_mx0w0 , 1'b1})
      + STAGE_LOOP_op_rshift_psp_1_sva;
  assign IDX_LOOP_idx2_9_0_sva_mx0w0 = nl_IDX_LOOP_idx2_9_0_sva_mx0w0[9:0];
  assign IDX_LOOP_f2_nor_cse_1 = ~((IDX_LOOP_idx2_acc_psp_sva[1:0]!=2'b00));
  assign IDX_LOOP_f2_nor_1_cse_1 = ~((IDX_LOOP_idx2_acc_psp_sva[1]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign IDX_LOOP_f2_nor_2_cse_1 = ~((IDX_LOOP_idx2_acc_psp_sva[0]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign IDX_LOOP_IDX_LOOP_and_126_nl = (reg_IDX_LOOP_1_lshift_idiv_ftd_7==3'b001);
  assign IDX_LOOP_IDX_LOOP_and_128_nl = (reg_IDX_LOOP_1_lshift_idiv_ftd_7==3'b010);
  assign IDX_LOOP_IDX_LOOP_and_130_nl = (reg_IDX_LOOP_1_lshift_idiv_ftd_7==3'b100);
  assign IDX_LOOP_mux1h_68_itm_mx0w0 = MUX1HOT_v_64_8_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
      twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_5_i_q_d,
      twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d, {IDX_LOOP_IDX_LOOP_nor_12_itm
      , IDX_LOOP_IDX_LOOP_and_126_nl , IDX_LOOP_IDX_LOOP_and_128_nl , IDX_LOOP_IDX_LOOP_and_104_itm
      , IDX_LOOP_IDX_LOOP_and_130_nl , IDX_LOOP_IDX_LOOP_and_106_itm , IDX_LOOP_IDX_LOOP_and_107_itm
      , IDX_LOOP_IDX_LOOP_and_108_itm});
  assign IDX_LOOP_f2_nor_12_cse_1 = ~((IDX_LOOP_idx2_9_0_2_sva[2:1]!=2'b00));
  assign IDX_LOOP_f2_nor_13_cse_1 = ~((IDX_LOOP_idx2_9_0_2_sva[2]) | (IDX_LOOP_idx2_9_0_2_sva[0]));
  assign IDX_LOOP_f2_nor_14_cse_1 = ~((IDX_LOOP_idx2_9_0_2_sva[1:0]!=2'b00));
  assign IDX_LOOP_f2_nor_24_cse_1 = ~((IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b00));
  assign IDX_LOOP_f2_nor_25_cse_1 = ~((IDX_LOOP_idx2_acc_1_psp_sva[1]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign IDX_LOOP_f2_nor_26_cse_1 = ~((IDX_LOOP_idx2_acc_1_psp_sva[0]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign IDX_LOOP_f2_nor_36_cse_1 = ~((IDX_LOOP_idx2_9_0_4_sva[2:1]!=2'b00));
  assign IDX_LOOP_f2_nor_37_cse_1 = ~((IDX_LOOP_idx2_9_0_4_sva[2]) | (IDX_LOOP_idx2_9_0_4_sva[0]));
  assign IDX_LOOP_f2_nor_38_cse_1 = ~((IDX_LOOP_idx2_9_0_4_sva[1:0]!=2'b00));
  assign IDX_LOOP_f2_nor_48_cse_1 = ~((IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b00));
  assign IDX_LOOP_f2_nor_49_cse_1 = ~((IDX_LOOP_idx2_acc_2_psp_sva[1]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign IDX_LOOP_f2_nor_50_cse_1 = ~((IDX_LOOP_idx2_acc_2_psp_sva[0]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign IDX_LOOP_f2_nor_60_cse_1 = ~((IDX_LOOP_idx2_9_0_6_sva[2:1]!=2'b00));
  assign IDX_LOOP_f2_nor_61_cse_1 = ~((IDX_LOOP_idx2_9_0_6_sva[2]) | (IDX_LOOP_idx2_9_0_6_sva[0]));
  assign IDX_LOOP_f2_nor_62_cse_1 = ~((IDX_LOOP_idx2_9_0_6_sva[1:0]!=2'b00));
  assign IDX_LOOP_f2_nor_72_cse_1 = ~((IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b00));
  assign IDX_LOOP_f2_nor_73_cse_1 = ~((IDX_LOOP_idx2_acc_3_psp_sva[1]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign IDX_LOOP_f2_nor_74_cse_1 = ~((IDX_LOOP_idx2_acc_3_psp_sva[0]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign IDX_LOOP_f2_nor_84_cse_1 = ~((IDX_LOOP_idx2_9_0_sva[2:1]!=2'b00));
  assign IDX_LOOP_f2_nor_85_cse_1 = ~((IDX_LOOP_idx2_9_0_sva[2]) | (IDX_LOOP_idx2_9_0_sva[0]));
  assign IDX_LOOP_f2_nor_86_cse_1 = ~((IDX_LOOP_idx2_9_0_sva[1:0]!=2'b00));
  assign nl_STAGE_LOOP_acc_nl = ({1'b1 , (~ STAGE_LOOP_i_3_0_sva_2)}) + 5'b01011;
  assign STAGE_LOOP_acc_nl = nl_STAGE_LOOP_acc_nl[4:0];
  assign STAGE_LOOP_acc_itm_4_1 = readslicef_5_1_4(STAGE_LOOP_acc_nl);
  assign and_dcpl = ~((fsm_output[8:7]!=2'b00));
  assign and_dcpl_1 = (fsm_output[6:5]==2'b01);
  assign or_tmp_2 = (fsm_output[4:0]!=5'b00000);
  assign or_tmp_3 = and_509_cse | (fsm_output[4:2]!=3'b000);
  assign or_tmp_4 = (fsm_output[4:1]!=4'b0000);
  assign and_dcpl_15 = ~((fsm_output[8:6]!=3'b000));
  assign or_tmp_11 = and_448_cse | (fsm_output[4:3]!=2'b00);
  assign or_tmp_16 = ((fsm_output[2:1]==2'b11)) | (fsm_output[4:3]!=2'b00);
  assign or_tmp_19 = (fsm_output[6:5]!=2'b00) | or_tmp_3;
  assign or_40_cse = ((fsm_output[2:0]==3'b111)) | (fsm_output[4:3]!=2'b00);
  assign or_44_cse = (fsm_output[4:2]!=3'b000);
  assign or_47_cse = (fsm_output[6]) | or_tmp_3;
  assign or_51_cse = (fsm_output[4:3]!=2'b00);
  assign or_tmp_26 = (fsm_output[7:1]!=7'b0000000);
  assign and_dcpl_55 = (fsm_output[6:5]==2'b10);
  assign and_dcpl_66 = (fsm_output[8:7]==2'b01);
  assign or_677_cse = (fsm_output[7:6]!=2'b00);
  assign nor_236_nl = ~((fsm_output[7:5]!=3'b000) | or_tmp_11);
  assign mux_180_cse = MUX_s_1_2_2(or_tmp_26, nor_236_nl, fsm_output[8]);
  assign and_dcpl_93 = ~((fsm_output[6:5]!=2'b00));
  assign and_dcpl_94 = and_dcpl_93 & and_dcpl;
  assign and_dcpl_95 = ~((fsm_output[1:0]!=2'b00));
  assign and_dcpl_96 = ~((fsm_output[4:3]!=2'b00));
  assign and_dcpl_97 = and_dcpl_96 & (~ (fsm_output[2]));
  assign and_dcpl_101 = and_dcpl_93 & (fsm_output[8:7]==2'b10);
  assign and_dcpl_102 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_103 = and_dcpl_96 & (fsm_output[2]);
  assign and_dcpl_104 = and_dcpl_103 & and_dcpl_102;
  assign and_dcpl_108 = and_dcpl_103 & and_dcpl_95;
  assign and_dcpl_109 = and_dcpl_108 & and_dcpl_94;
  assign and_dcpl_113 = and_dcpl_1 & and_dcpl;
  assign and_dcpl_114 = and_dcpl_108 & and_dcpl_113;
  assign and_dcpl_116 = and_dcpl_55 & and_dcpl;
  assign and_dcpl_117 = and_dcpl_108 & and_dcpl_116;
  assign and_dcpl_119 = and_513_cse & and_dcpl;
  assign and_dcpl_120 = and_dcpl_108 & and_dcpl_119;
  assign and_dcpl_122 = and_dcpl_93 & and_dcpl_66;
  assign and_dcpl_123 = and_dcpl_108 & and_dcpl_122;
  assign and_dcpl_124 = and_dcpl_1 & and_dcpl_66;
  assign and_dcpl_125 = and_dcpl_108 & and_dcpl_124;
  assign and_dcpl_126 = and_dcpl_55 & and_dcpl_66;
  assign and_dcpl_127 = and_dcpl_108 & and_dcpl_126;
  assign and_dcpl_128 = and_513_cse & and_dcpl_66;
  assign and_dcpl_129 = and_dcpl_108 & and_dcpl_128;
  assign and_dcpl_134 = (fsm_output[4:3]==2'b01);
  assign and_dcpl_135 = and_dcpl_134 & (~ (fsm_output[2]));
  assign and_dcpl_138 = and_dcpl_135 & and_dcpl_95;
  assign and_dcpl_151 = ~((fsm_output[6:4]!=3'b000) | (~ and_dcpl));
  assign and_dcpl_153 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_154 = and_dcpl_97 & and_dcpl_153;
  assign and_dcpl_155 = and_dcpl_154 & and_dcpl_94;
  assign and_dcpl_157 = and_dcpl_97 & and_509_cse;
  assign and_dcpl_158 = and_dcpl_157 & and_dcpl_94;
  assign and_dcpl_159 = and_dcpl_104 & and_dcpl_94;
  assign not_tmp_162 = ~((z_out_6[1]) & (fsm_output[3]));
  assign not_tmp_164 = ~((z_out_6[0]) & (fsm_output[3]));
  assign nand_44_cse = ~((IDX_LOOP_idx2_9_0_2_sva[2:0]==3'b111));
  assign mux_256_cse = MUX_s_1_2_2((reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1]), (IDX_LOOP_idx1_acc_2_psp_sva[0]),
      fsm_output[7]);
  assign and_dcpl_176 = and_dcpl_97 & (fsm_output[1]) & (~ (fsm_output[8]));
  assign not_tmp_180 = ~((STAGE_LOOP_op_rshift_psp_1_sva[0]) & (fsm_output[0]));
  assign and_481_cse = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7==2'b11);
  assign or_290_cse = (~ (IDX_LOOP_idx1_acc_2_psp_sva[0])) | (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]))
      | (fsm_output[0]);
  assign or_288_cse = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b11) | (fsm_output[0]);
  assign or_286_cse = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b11) | (fsm_output[0]);
  assign and_dcpl_179 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_183 = and_dcpl_97 & and_dcpl_102;
  assign and_dcpl_184 = and_dcpl_183 & and_dcpl_113;
  assign and_dcpl_185 = and_dcpl_183 & and_dcpl_116;
  assign and_dcpl_187 = and_dcpl_183 & and_dcpl_119;
  assign and_dcpl_188 = and_dcpl_183 & and_dcpl_122;
  assign and_dcpl_190 = and_dcpl_183 & and_dcpl_124;
  assign and_dcpl_191 = and_dcpl_183 & and_dcpl_126;
  assign and_dcpl_193 = and_dcpl_183 & and_dcpl_128;
  assign and_dcpl_194 = and_dcpl_183 & and_dcpl_101;
  assign and_dcpl_198 = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1]) & (fsm_output[6:5]==2'b01)
      & and_dcpl;
  assign and_dcpl_200 = and_dcpl_97 & and_dcpl_153 & (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]);
  assign and_dcpl_202 = (fsm_output[1]) & (~ (fsm_output[6]));
  assign and_dcpl_203 = and_dcpl_202 & (fsm_output[5]);
  assign and_dcpl_204 = and_dcpl_203 & and_dcpl;
  assign or_dcpl_74 = (fsm_output[0]) | (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]));
  assign and_dcpl_207 = and_dcpl_157 & and_dcpl_116;
  assign and_dcpl_208 = (IDX_LOOP_idx1_acc_psp_3_sva[0]) & (fsm_output[6]);
  assign and_dcpl_210 = and_dcpl_208 & (fsm_output[5]) & and_dcpl;
  assign and_dcpl_212 = and_dcpl_97 & and_dcpl_153 & (IDX_LOOP_idx1_acc_psp_3_sva[1]);
  assign and_dcpl_214 = (fsm_output[1]) & (fsm_output[6]);
  assign and_dcpl_215 = and_dcpl_214 & (fsm_output[5]);
  assign and_dcpl_216 = and_dcpl_215 & and_dcpl;
  assign or_dcpl_76 = (fsm_output[0]) | (~ (IDX_LOOP_idx1_acc_psp_3_sva[1]));
  assign and_dcpl_217 = and_dcpl_97 & (or_dcpl_76 | (~ (IDX_LOOP_idx1_acc_psp_3_sva[0])));
  assign and_dcpl_219 = and_dcpl_157 & and_dcpl_122;
  assign and_dcpl_220 = (IDX_LOOP_idx1_acc_2_psp_sva[0]) & (~ (fsm_output[6]));
  assign and_dcpl_222 = and_dcpl_220 & (fsm_output[5]) & and_dcpl_66;
  assign and_dcpl_224 = and_dcpl_203 & and_dcpl_66;
  assign and_dcpl_225 = and_dcpl_97 & (or_dcpl_74 | (~ (IDX_LOOP_idx1_acc_2_psp_sva[0])));
  assign and_dcpl_227 = and_dcpl_157 & and_dcpl_126;
  assign and_dcpl_228 = (IDX_LOOP_idx1_acc_psp_7_sva[0]) & (fsm_output[6]);
  assign and_dcpl_230 = and_dcpl_228 & (fsm_output[5]) & and_dcpl_66;
  assign and_dcpl_232 = and_dcpl_97 & and_dcpl_153 & (IDX_LOOP_idx1_acc_psp_7_sva[1]);
  assign and_dcpl_234 = and_dcpl_215 & and_dcpl_66;
  assign or_dcpl_79 = (fsm_output[0]) | (~ (IDX_LOOP_idx1_acc_psp_7_sva[1]));
  assign and_dcpl_235 = and_dcpl_97 & (or_dcpl_79 | (~ (IDX_LOOP_idx1_acc_psp_7_sva[0])));
  assign nor_tmp_55 = (fsm_output[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0]);
  assign or_tmp_248 = (fsm_output[0]) | (STAGE_LOOP_op_rshift_psp_1_sva[0]);
  assign and_dcpl_241 = and_dcpl_96 & and_dcpl_179;
  assign and_dcpl_247 = and_dcpl_157 & and_dcpl_113;
  assign and_dcpl_249 = and_dcpl_208 & (~ (fsm_output[5])) & and_dcpl;
  assign and_dcpl_251 = and_dcpl_214 & (~ (fsm_output[5]));
  assign and_dcpl_252 = and_dcpl_251 & and_dcpl;
  assign and_dcpl_254 = and_dcpl_157 & and_dcpl_119;
  assign and_dcpl_256 = and_dcpl_220 & (~ (fsm_output[5])) & and_dcpl_66;
  assign and_dcpl_259 = and_dcpl_202 & (~ (fsm_output[5])) & and_dcpl_66;
  assign and_dcpl_261 = and_dcpl_157 & and_dcpl_124;
  assign and_dcpl_263 = and_dcpl_228 & (~ (fsm_output[5])) & and_dcpl_66;
  assign and_dcpl_265 = and_dcpl_251 & and_dcpl_66;
  assign and_dcpl_267 = and_dcpl_157 & and_dcpl_128;
  assign nand_23_cse = ~((IDX_LOOP_idx2_9_0_2_sva[2]) & (IDX_LOOP_idx2_9_0_2_sva[0]));
  assign or_362_cse = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7!=2'b10);
  assign and_dcpl_271 = and_dcpl_97 & and_dcpl_153 & (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]));
  assign or_dcpl_81 = (fsm_output[0]) | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]);
  assign and_dcpl_275 = (~ (IDX_LOOP_idx1_acc_psp_3_sva[0])) & (fsm_output[6]);
  assign and_dcpl_277 = and_dcpl_275 & (fsm_output[5]) & and_dcpl;
  assign or_dcpl_83 = or_dcpl_76 | (IDX_LOOP_idx1_acc_psp_3_sva[0]);
  assign and_dcpl_279 = and_dcpl_97 & or_dcpl_83;
  assign or_dcpl_84 = or_dcpl_81 | (~ (IDX_LOOP_idx1_acc_2_psp_sva[0]));
  assign and_dcpl_282 = and_dcpl_97 & or_dcpl_84;
  assign and_dcpl_284 = (~ (IDX_LOOP_idx1_acc_psp_7_sva[0])) & (fsm_output[6]);
  assign and_dcpl_286 = and_dcpl_284 & (fsm_output[5]) & and_dcpl_66;
  assign or_dcpl_85 = or_dcpl_79 | (IDX_LOOP_idx1_acc_psp_7_sva[0]);
  assign and_dcpl_288 = and_dcpl_97 & or_dcpl_85;
  assign and_dcpl_293 = and_dcpl_275 & (~ (fsm_output[5])) & and_dcpl;
  assign and_dcpl_299 = and_dcpl_284 & (~ (fsm_output[5])) & and_dcpl_66;
  assign or_425_cse = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b011);
  assign or_439_cse = (IDX_LOOP_idx1_acc_2_psp_sva[0]) | (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]))
      | (fsm_output[0]);
  assign or_437_cse = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b01) | (fsm_output[0]);
  assign or_435_cse = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b01) | (fsm_output[0]);
  assign and_dcpl_306 = (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1])) & (fsm_output[6:5]==2'b01)
      & and_dcpl;
  assign and_dcpl_311 = and_dcpl_97 & and_dcpl_153 & (~ (IDX_LOOP_idx1_acc_psp_3_sva[1]));
  assign or_dcpl_87 = (fsm_output[0]) | (IDX_LOOP_idx1_acc_psp_3_sva[1]);
  assign and_dcpl_313 = and_dcpl_97 & (or_dcpl_87 | (~ (IDX_LOOP_idx1_acc_psp_3_sva[0])));
  assign and_dcpl_315 = ~((IDX_LOOP_idx1_acc_2_psp_sva[0]) | (fsm_output[6]));
  assign and_dcpl_317 = and_dcpl_315 & (fsm_output[5]) & and_dcpl_66;
  assign and_dcpl_319 = and_dcpl_97 & (or_dcpl_74 | (IDX_LOOP_idx1_acc_2_psp_sva[0]));
  assign and_dcpl_322 = and_dcpl_97 & and_dcpl_153 & (~ (IDX_LOOP_idx1_acc_psp_7_sva[1]));
  assign or_dcpl_90 = (fsm_output[0]) | (IDX_LOOP_idx1_acc_psp_7_sva[1]);
  assign and_dcpl_324 = and_dcpl_97 & (or_dcpl_90 | (~ (IDX_LOOP_idx1_acc_psp_7_sva[0])));
  assign or_tmp_395 = (fsm_output[0]) | (IDX_LOOP_idx2_acc_tmp[1:0]!=2'b01) | (STAGE_LOOP_op_rshift_psp_1_sva[0]);
  assign and_dcpl_331 = and_dcpl_315 & (~ (fsm_output[5])) & and_dcpl_66;
  assign or_504_cse = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b001);
  assign or_520_cse = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7!=2'b00);
  assign or_519_cse = (IDX_LOOP_idx1_acc_2_psp_sva[0]) | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0])
      | (fsm_output[0]);
  assign or_517_cse = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b00) | (fsm_output[0]);
  assign or_515_cse = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b00) | (fsm_output[0]);
  assign and_dcpl_342 = and_dcpl_97 & (or_dcpl_87 | (IDX_LOOP_idx1_acc_psp_3_sva[0]));
  assign and_dcpl_345 = and_dcpl_97 & (or_dcpl_81 | (IDX_LOOP_idx1_acc_2_psp_sva[0]));
  assign and_dcpl_348 = and_dcpl_97 & (or_dcpl_90 | (IDX_LOOP_idx1_acc_psp_7_sva[0]));
  assign and_tmp_7 = (fsm_output[6:5]==2'b11) & or_44_cse;
  assign or_dcpl_103 = or_44_cse | (~ (fsm_output[1])) | (fsm_output[0]) | (fsm_output[6])
      | (fsm_output[5]) | (fsm_output[7]) | (fsm_output[8]);
  assign and_375_nl = (fsm_output[6]) & or_tmp_4;
  assign mux_462_nl = MUX_s_1_2_2(and_375_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_463_nl = MUX_s_1_2_2(or_tmp_19, (~ mux_462_nl), fsm_output[7]);
  assign and_dcpl_367 = mux_463_nl & (~ (fsm_output[8]));
  assign mux_464_nl = MUX_s_1_2_2(or_tmp_19, (~ and_tmp_7), fsm_output[7]);
  assign and_dcpl_368 = mux_464_nl & (~ (fsm_output[8]));
  assign and_tmp_9 = (fsm_output[6]) & or_tmp_2;
  assign mux_467_nl = MUX_s_1_2_2(or_tmp_3, (~ or_44_cse), fsm_output[5]);
  assign and_dcpl_374 = mux_467_nl & and_dcpl_15;
  assign and_tmp_10 = (fsm_output[6]) & or_tmp_3;
  assign mux_470_nl = MUX_s_1_2_2((~ or_tmp_3), or_44_cse, fsm_output[6]);
  assign mux_471_nl = MUX_s_1_2_2(mux_470_nl, (fsm_output[6]), fsm_output[5]);
  assign and_dcpl_377 = (~ mux_471_nl) & and_dcpl;
  assign and_tmp_11 = (fsm_output[6]) & or_44_cse;
  assign mux_474_nl = MUX_s_1_2_2(or_47_cse, (~ and_tmp_11), fsm_output[5]);
  assign and_dcpl_380 = mux_474_nl & and_dcpl;
  assign or_tmp_502 = (fsm_output[6:2]!=5'b00000);
  assign mux_479_nl = MUX_s_1_2_2(or_tmp_19, (~ or_tmp_502), fsm_output[7]);
  assign and_dcpl_383 = mux_479_nl & (~ (fsm_output[8]));
  assign or_tmp_505 = (fsm_output[6]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[3]);
  assign mux_tmp_457 = MUX_s_1_2_2((fsm_output[6]), or_tmp_505, fsm_output[5]);
  assign mux_485_nl = MUX_s_1_2_2(or_tmp_19, (~ mux_tmp_457), fsm_output[7]);
  assign and_dcpl_386 = mux_485_nl & (~ (fsm_output[8]));
  assign nand_14_nl = ~((fsm_output[6:5]==2'b11) & or_tmp_3);
  assign mux_487_nl = MUX_s_1_2_2(or_tmp_19, nand_14_nl, fsm_output[7]);
  assign and_dcpl_387 = mux_487_nl & (~ (fsm_output[8]));
  assign mux_tmp_461 = MUX_s_1_2_2(and_tmp_11, (fsm_output[6]), fsm_output[5]);
  assign mux_489_nl = MUX_s_1_2_2(or_tmp_19, (~ mux_tmp_461), fsm_output[7]);
  assign and_dcpl_388 = mux_489_nl & (~ (fsm_output[8]));
  assign not_tmp_290 = ~((fsm_output[6:5]!=2'b00) | or_tmp_16);
  assign and_dcpl_390 = ~((~(or_tmp_502 ^ (fsm_output[7]))) | (fsm_output[8]));
  assign or_587_nl = (fsm_output[2:1]!=2'b00);
  assign mux_491_nl = MUX_s_1_2_2((fsm_output[4]), or_51_cse, or_587_nl);
  assign not_tmp_292 = ~((fsm_output[6:5]!=2'b00) | mux_491_nl);
  assign not_tmp_296 = ~((fsm_output[6:5]!=2'b00) | or_tmp_11);
  assign not_tmp_298 = ~((fsm_output[6:5]!=2'b00) | or_40_cse);
  assign or_tmp_516 = (fsm_output[6:3]!=4'b0000);
  assign mux_502_nl = MUX_s_1_2_2((~ or_tmp_11), or_44_cse, fsm_output[6]);
  assign mux_503_nl = MUX_s_1_2_2(mux_502_nl, (fsm_output[6]), fsm_output[5]);
  assign and_dcpl_404 = (~ mux_503_nl) & and_dcpl;
  assign mux_505_nl = MUX_s_1_2_2(or_tmp_502, (~ mux_tmp_457), fsm_output[7]);
  assign and_dcpl_407 = mux_505_nl & (~ (fsm_output[8]));
  assign mux_506_nl = MUX_s_1_2_2(or_tmp_502, (~ and_tmp_7), fsm_output[7]);
  assign and_dcpl_408 = mux_506_nl & (~ (fsm_output[8]));
  assign and_dcpl_413 = and_dcpl_241 & (fsm_output[0]) & (fsm_output[5]) & (~ (fsm_output[8]));
  assign mux_515_nl = MUX_s_1_2_2(not_tmp_296, mux_tmp_457, fsm_output[7]);
  assign and_dcpl_416 = ~(mux_515_nl | (fsm_output[8]));
  assign mux_516_nl = MUX_s_1_2_2(not_tmp_296, and_tmp_7, fsm_output[7]);
  assign and_dcpl_417 = ~(mux_516_nl | (fsm_output[8]));
  assign mux_520_nl = MUX_s_1_2_2(not_tmp_290, and_tmp_7, fsm_output[7]);
  assign and_dcpl_419 = ~(mux_520_nl | (fsm_output[8]));
  assign and_tmp_14 = (fsm_output[6]) & or_51_cse;
  assign mux_523_nl = MUX_s_1_2_2((fsm_output[4]), or_51_cse, or_200_cse);
  assign nor_112_nl = ~((fsm_output[6:5]!=2'b00) | mux_523_nl);
  assign mux_524_nl = MUX_s_1_2_2(nor_112_nl, and_tmp_7, fsm_output[7]);
  assign and_dcpl_423 = ~(mux_524_nl | (fsm_output[8]));
  assign and_dcpl_430 = and_dcpl_97 & or_677_cse & and_509_cse & (~ (fsm_output[5]))
      & (~ (fsm_output[8]));
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_104 & and_dcpl_101;
  assign GROUP_LOOP_j_10_0_sva_9_0_mx0c0 = and_dcpl_183 & and_dcpl_94;
  assign IDX_LOOP_modulo_dev_return_1_sva_mx0c1 = and_dcpl_135 & and_dcpl_102 & (~
      (fsm_output[8]));
  assign and_359_nl = and_dcpl_311 & and_dcpl_293;
  assign and_360_nl = and_dcpl_342 & and_dcpl_252;
  assign and_361_nl = and_dcpl_271 & and_dcpl_331;
  assign and_362_nl = and_dcpl_345 & and_dcpl_259;
  assign and_363_nl = and_dcpl_322 & and_dcpl_299;
  assign and_364_nl = and_dcpl_348 & and_dcpl_265;
  assign vec_rsc_0_0_i_radr_d = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_tmp[8:2]), IDX_LOOP_idx1_acc_psp_8_sva,
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_155 , and_dcpl_158 , and_dcpl_247 ,
      and_359_nl , and_360_nl , and_dcpl_254 , and_361_nl , and_362_nl , and_dcpl_261
      , and_363_nl , and_364_nl , and_dcpl_267});
  assign and_247_nl = and_dcpl_154 & and_dcpl_113;
  assign and_248_nl = and_dcpl_154 & and_dcpl_119;
  assign and_249_nl = and_dcpl_154 & and_dcpl_124;
  assign and_250_nl = and_dcpl_154 & and_dcpl_128;
  assign vec_rsc_0_0_i_wadr_d_pff = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_psp_sva[8:2]),
      IDX_LOOP_idx1_acc_psp_8_sva, (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]),
      (IDX_LOOP_idx1_acc_psp_3_sva[8:2]), (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]),
      (IDX_LOOP_idx1_acc_2_psp_sva[7:1]), (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]),
      (IDX_LOOP_idx1_acc_psp_7_sva[8:2]), (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_184
      , and_247_nl , and_dcpl_185 , and_dcpl_187 , and_248_nl , and_dcpl_188 , and_dcpl_190
      , and_249_nl , and_dcpl_191 , and_dcpl_193 , and_250_nl , and_dcpl_194});
  assign and_246_nl = and_dcpl_241 & (~ (fsm_output[0])) & (fsm_output[5]) & (~ (fsm_output[8]));
  assign vec_rsc_0_0_i_d_d_pff = MUX_v_64_2_2(IDX_LOOP_1_IDX_LOOP_rem_1_cmp_z, IDX_LOOP_modulo_dev_return_1_sva,
      and_246_nl);
  assign or_549_nl = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1]) | (fsm_output[8]);
  assign or_548_nl = (IDX_LOOP_idx1_acc_2_psp_sva[0]) | (fsm_output[8]);
  assign mux_432_nl = MUX_s_1_2_2(or_549_nl, or_548_nl, fsm_output[7]);
  assign nor_130_nl = ~((reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]) | mux_432_nl);
  assign nor_131_nl = ~((IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b00) | (fsm_output[8]));
  assign nor_132_nl = ~((IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b00) | (fsm_output[8]));
  assign mux_431_nl = MUX_s_1_2_2(nor_131_nl, nor_132_nl, fsm_output[7]);
  assign mux_433_nl = MUX_s_1_2_2(nor_130_nl, mux_431_nl, fsm_output[6]);
  assign and_453_nl = (fsm_output[1]) & (fsm_output[5]) & mux_433_nl;
  assign or_544_nl = (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b000) | (~ (fsm_output[8]));
  assign or_542_nl = (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b000) | (fsm_output[8]);
  assign mux_428_nl = MUX_s_1_2_2(or_544_nl, or_542_nl, fsm_output[7]);
  assign or_541_nl = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b000) | (fsm_output[8]);
  assign or_540_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b000) | (fsm_output[8]);
  assign mux_427_nl = MUX_s_1_2_2(or_541_nl, or_540_nl, fsm_output[7]);
  assign mux_429_nl = MUX_s_1_2_2(mux_428_nl, mux_427_nl, fsm_output[6]);
  assign or_539_nl = (IDX_LOOP_idx2_acc_psp_sva[1:0]!=2'b00) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign or_538_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b00) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign mux_425_nl = MUX_s_1_2_2(or_539_nl, or_538_nl, fsm_output[7]);
  assign or_537_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b00) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign or_536_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b00) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign mux_424_nl = MUX_s_1_2_2(or_537_nl, or_536_nl, fsm_output[7]);
  assign mux_426_nl = MUX_s_1_2_2(mux_425_nl, mux_424_nl, fsm_output[6]);
  assign mux_430_nl = MUX_s_1_2_2(mux_429_nl, mux_426_nl, fsm_output[5]);
  assign nor_133_nl = ~((fsm_output[1]) | mux_430_nl);
  assign mux_434_nl = MUX_s_1_2_2(and_453_nl, nor_133_nl, fsm_output[0]);
  assign vec_rsc_0_0_i_we_d_pff = mux_434_nl & and_dcpl_97;
  assign nor_128_nl = ~((fsm_output[0]) | IDX_LOOP_f2_IDX_LOOP_f2_nor_cse);
  assign or_570_nl = (fsm_output[0]) | (IDX_LOOP_idx2_acc_tmp[1:0]!=2'b00) | (STAGE_LOOP_op_rshift_psp_1_sva[0]);
  assign mux_448_nl = MUX_s_1_2_2(nor_128_nl, or_570_nl, or_520_cse);
  assign or_568_nl = (IDX_LOOP_idx1_acc_2_psp_sva[0]) | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]);
  assign mux_446_nl = MUX_s_1_2_2(mux_293_cse, or_tmp_248, or_568_nl);
  assign or_566_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b00);
  assign mux_447_nl = MUX_s_1_2_2(mux_446_nl, or_519_cse, or_566_nl);
  assign mux_449_nl = MUX_s_1_2_2(mux_448_nl, mux_447_nl, fsm_output[7]);
  assign or_565_nl = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b00);
  assign mux_442_nl = MUX_s_1_2_2(mux_289_cse, or_tmp_248, or_565_nl);
  assign or_563_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b00);
  assign mux_443_nl = MUX_s_1_2_2(mux_442_nl, or_517_cse, or_563_nl);
  assign or_561_nl = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b00);
  assign mux_439_nl = MUX_s_1_2_2(mux_286_cse, or_tmp_248, or_561_nl);
  assign or_559_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b00);
  assign mux_440_nl = MUX_s_1_2_2(mux_439_nl, or_515_cse, or_559_nl);
  assign mux_444_nl = MUX_s_1_2_2(mux_443_nl, mux_440_nl, fsm_output[7]);
  assign mux_450_nl = MUX_s_1_2_2(mux_449_nl, mux_444_nl, fsm_output[6]);
  assign or_558_nl = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b000) | (~ IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0]));
  assign or_556_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b000) | (~ IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0]));
  assign mux_436_nl = MUX_s_1_2_2(or_558_nl, or_556_nl, fsm_output[7]);
  assign or_554_nl = (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b000) | (~ IDX_LOOP_slc_IDX_LOOP_acc_8_itm)
      | (~ (fsm_output[0]));
  assign or_552_nl = (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b000) | (~ IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm)
      | (~ (fsm_output[0]));
  assign mux_435_nl = MUX_s_1_2_2(or_554_nl, or_552_nl, fsm_output[7]);
  assign mux_437_nl = MUX_s_1_2_2(mux_436_nl, mux_435_nl, fsm_output[6]);
  assign mux_451_nl = MUX_s_1_2_2(mux_450_nl, mux_437_nl, fsm_output[5]);
  assign vec_rsc_0_0_i_re_d_pff = (~ mux_451_nl) & and_dcpl_176;
  assign and_345_nl = and_dcpl_271 & and_dcpl_306;
  assign and_347_nl = and_dcpl_97 & (or_dcpl_81 | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1]))
      & and_dcpl_204;
  assign and_348_nl = and_dcpl_311 & and_dcpl_277;
  assign and_350_nl = and_dcpl_342 & and_dcpl_216;
  assign and_351_nl = and_dcpl_271 & and_dcpl_317;
  assign and_353_nl = and_dcpl_345 & and_dcpl_224;
  assign and_354_nl = and_dcpl_322 & and_dcpl_286;
  assign and_356_nl = and_dcpl_348 & and_dcpl_234;
  assign vec_rsc_0_1_i_radr_d = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_tmp[8:2]), IDX_LOOP_idx1_acc_psp_8_sva,
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_155 , and_345_nl , and_347_nl , and_dcpl_207
      , and_348_nl , and_350_nl , and_dcpl_219 , and_351_nl , and_353_nl , and_dcpl_227
      , and_354_nl , and_356_nl});
  assign and_190_nl = and_dcpl_154 & and_dcpl_116;
  assign and_193_nl = and_dcpl_154 & and_dcpl_122;
  assign and_196_nl = and_dcpl_154 & and_dcpl_126;
  assign and_199_nl = and_dcpl_154 & and_dcpl_101;
  assign vec_rsc_0_1_i_wadr_d_pff = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), IDX_LOOP_idx1_acc_psp_8_sva, (IDX_LOOP_idx2_acc_1_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]), {and_dcpl_184
      , and_dcpl_185 , and_190_nl , and_dcpl_187 , and_dcpl_188 , and_193_nl , and_dcpl_190
      , and_dcpl_191 , and_196_nl , and_dcpl_193 , and_dcpl_194 , and_199_nl});
  assign and_186_nl = (or_677_cse ^ (fsm_output[8])) & and_dcpl_96 & and_dcpl_179
      & (~ (fsm_output[0])) & (~ (fsm_output[5]));
  assign vec_rsc_0_1_i_d_d_pff = MUX_v_64_2_2(IDX_LOOP_1_IDX_LOOP_rem_1_cmp_z, IDX_LOOP_modulo_dev_return_1_sva,
      and_186_nl);
  assign or_512_nl = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b00) | (~ (fsm_output[7]));
  assign or_510_nl = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]) | mux_256_cse;
  assign mux_409_nl = MUX_s_1_2_2(or_512_nl, or_510_nl, fsm_output[6]);
  assign or_509_nl = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b00) | (fsm_output[7:6]!=2'b00);
  assign mux_410_nl = MUX_s_1_2_2(mux_409_nl, or_509_nl, fsm_output[8]);
  assign nor_138_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | mux_410_nl);
  assign or_506_nl = (~ (fsm_output[7])) | (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b001);
  assign or_502_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b001);
  assign mux_404_nl = MUX_s_1_2_2(or_504_cse, or_502_nl, fsm_output[7]);
  assign mux_405_nl = MUX_s_1_2_2(or_506_nl, mux_404_nl, fsm_output[6]);
  assign or_500_nl = (fsm_output[7:6]!=2'b00) | (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b001);
  assign mux_406_nl = MUX_s_1_2_2(mux_405_nl, or_500_nl, fsm_output[8]);
  assign or_497_nl = (IDX_LOOP_idx2_acc_psp_sva[1:0]!=2'b00) | (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign or_495_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b00) | (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign mux_402_nl = MUX_s_1_2_2(or_497_nl, or_495_nl, fsm_output[7]);
  assign or_493_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b00) | (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign or_491_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b00) | (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign mux_401_nl = MUX_s_1_2_2(or_493_nl, or_491_nl, fsm_output[7]);
  assign mux_403_nl = MUX_s_1_2_2(mux_402_nl, mux_401_nl, fsm_output[6]);
  assign or_498_nl = (fsm_output[8]) | mux_403_nl;
  assign mux_407_nl = MUX_s_1_2_2(mux_406_nl, or_498_nl, fsm_output[5]);
  assign nor_139_nl = ~((fsm_output[1]) | mux_407_nl);
  assign mux_411_nl = MUX_s_1_2_2(nor_138_nl, nor_139_nl, fsm_output[0]);
  assign vec_rsc_0_1_i_we_d_pff = mux_411_nl & and_dcpl_97;
  assign nor_134_nl = ~((IDX_LOOP_idx2_acc_tmp[1:0]!=2'b00) | (fsm_output[0]));
  assign nor_135_nl = ~((IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b00) | (~ IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0])));
  assign mux_421_nl = MUX_s_1_2_2(nor_134_nl, nor_135_nl, fsm_output[7]);
  assign nor_136_nl = ~((IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b00) | (~ IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0])));
  assign nor_137_nl = ~((IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b00) | (~ IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0])));
  assign mux_420_nl = MUX_s_1_2_2(nor_136_nl, nor_137_nl, fsm_output[7]);
  assign mux_422_nl = MUX_s_1_2_2(mux_421_nl, mux_420_nl, fsm_output[6]);
  assign nand_10_nl = ~((STAGE_LOOP_op_rshift_psp_1_sva[0]) & mux_422_nl);
  assign and_343_nl = (fsm_output[0]) & or_504_cse;
  assign mux_416_nl = MUX_s_1_2_2((fsm_output[0]), and_343_nl, IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm);
  assign or_522_nl = (fsm_output[0]) | (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b001);
  assign mux_417_nl = MUX_s_1_2_2(mux_416_nl, or_522_nl, or_520_cse);
  assign and_454_nl = ((IDX_LOOP_idx1_acc_2_psp_sva[0]) | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0])
      | (~ IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm)) & (fsm_output[0]);
  assign nor_99_nl = ~((IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b001));
  assign mux_415_nl = MUX_s_1_2_2(or_519_cse, and_454_nl, nor_99_nl);
  assign mux_418_nl = MUX_s_1_2_2(mux_417_nl, mux_415_nl, fsm_output[7]);
  assign and_455_nl = ((IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b00) | (~ IDX_LOOP_slc_IDX_LOOP_acc_8_itm))
      & (fsm_output[0]);
  assign nor_97_nl = ~((IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b001));
  assign mux_413_nl = MUX_s_1_2_2(or_517_cse, and_455_nl, nor_97_nl);
  assign and_456_nl = ((IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b00) | (~ IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm))
      & (fsm_output[0]);
  assign nor_95_nl = ~((IDX_LOOP_idx2_9_0_sva[2:0]!=3'b001));
  assign mux_412_nl = MUX_s_1_2_2(or_515_cse, and_456_nl, nor_95_nl);
  assign mux_414_nl = MUX_s_1_2_2(mux_413_nl, mux_412_nl, fsm_output[7]);
  assign mux_419_nl = MUX_s_1_2_2(mux_418_nl, mux_414_nl, fsm_output[6]);
  assign mux_423_nl = MUX_s_1_2_2(nand_10_nl, mux_419_nl, fsm_output[5]);
  assign vec_rsc_0_1_i_re_d_pff = (~ mux_423_nl) & and_dcpl_176;
  assign and_334_nl = and_dcpl_311 & and_dcpl_249;
  assign and_335_nl = and_dcpl_313 & and_dcpl_252;
  assign and_338_nl = and_dcpl_200 & and_dcpl_331;
  assign and_339_nl = and_dcpl_319 & and_dcpl_259;
  assign and_340_nl = and_dcpl_322 & and_dcpl_263;
  assign and_341_nl = and_dcpl_324 & and_dcpl_265;
  assign vec_rsc_0_2_i_radr_d = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_tmp[8:2]), IDX_LOOP_idx1_acc_psp_8_sva,
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_155 , and_dcpl_158 , and_dcpl_247 ,
      and_334_nl , and_335_nl , and_dcpl_254 , and_338_nl , and_339_nl , and_dcpl_261
      , and_340_nl , and_341_nl , and_dcpl_267});
  assign nor_142_nl = ~((reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1]) | (fsm_output[8]));
  assign nor_143_nl = ~((IDX_LOOP_idx1_acc_2_psp_sva[0]) | (fsm_output[8]));
  assign mux_380_nl = MUX_s_1_2_2(nor_142_nl, nor_143_nl, fsm_output[7]);
  assign and_459_nl = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]) & mux_380_nl;
  assign nor_144_nl = ~((IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b01) | (fsm_output[8]));
  assign nor_145_nl = ~((IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b01) | (fsm_output[8]));
  assign mux_379_nl = MUX_s_1_2_2(nor_144_nl, nor_145_nl, fsm_output[7]);
  assign mux_381_nl = MUX_s_1_2_2(and_459_nl, mux_379_nl, fsm_output[6]);
  assign and_458_nl = (fsm_output[1]) & (fsm_output[5]) & mux_381_nl;
  assign or_465_nl = (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b010) | (~ (fsm_output[8]));
  assign or_463_nl = (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b010) | (fsm_output[8]);
  assign mux_376_nl = MUX_s_1_2_2(or_465_nl, or_463_nl, fsm_output[7]);
  assign or_462_nl = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b010) | (fsm_output[8]);
  assign or_461_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b010) | (fsm_output[8]);
  assign mux_375_nl = MUX_s_1_2_2(or_462_nl, or_461_nl, fsm_output[7]);
  assign mux_377_nl = MUX_s_1_2_2(mux_376_nl, mux_375_nl, fsm_output[6]);
  assign or_460_nl = (IDX_LOOP_idx2_acc_psp_sva[1:0]!=2'b01) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign or_459_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b01) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign mux_373_nl = MUX_s_1_2_2(or_460_nl, or_459_nl, fsm_output[7]);
  assign or_458_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b01) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign or_457_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b01) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign mux_372_nl = MUX_s_1_2_2(or_458_nl, or_457_nl, fsm_output[7]);
  assign mux_374_nl = MUX_s_1_2_2(mux_373_nl, mux_372_nl, fsm_output[6]);
  assign mux_378_nl = MUX_s_1_2_2(mux_377_nl, mux_374_nl, fsm_output[5]);
  assign nor_146_nl = ~((fsm_output[1]) | mux_378_nl);
  assign mux_382_nl = MUX_s_1_2_2(and_458_nl, nor_146_nl, fsm_output[0]);
  assign vec_rsc_0_2_i_we_d_pff = mux_382_nl & and_dcpl_97;
  assign nor_140_nl = ~((fsm_output[0]) | (~((IDX_LOOP_idx2_acc_tmp[1:0]!=2'b01)
      | (STAGE_LOOP_op_rshift_psp_1_sva[0]))));
  assign mux_396_nl = MUX_s_1_2_2(or_tmp_395, nor_140_nl, reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]);
  assign mux_397_nl = MUX_s_1_2_2(mux_396_nl, or_tmp_395, reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1]);
  assign nor_94_nl = ~((IDX_LOOP_idx1_acc_2_psp_sva[0]) | (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0])));
  assign mux_394_nl = MUX_s_1_2_2(or_tmp_248, mux_293_cse, nor_94_nl);
  assign or_485_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b01);
  assign mux_395_nl = MUX_s_1_2_2(mux_394_nl, or_439_cse, or_485_nl);
  assign mux_398_nl = MUX_s_1_2_2(mux_397_nl, mux_395_nl, fsm_output[7]);
  assign or_483_nl = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b01);
  assign mux_390_nl = MUX_s_1_2_2(mux_289_cse, or_tmp_248, or_483_nl);
  assign nor_93_nl = ~((IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b01));
  assign mux_391_nl = MUX_s_1_2_2(or_437_cse, mux_390_nl, nor_93_nl);
  assign or_481_nl = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b01);
  assign mux_387_nl = MUX_s_1_2_2(mux_286_cse, or_tmp_248, or_481_nl);
  assign or_479_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b01);
  assign mux_388_nl = MUX_s_1_2_2(mux_387_nl, or_435_cse, or_479_nl);
  assign mux_392_nl = MUX_s_1_2_2(mux_391_nl, mux_388_nl, fsm_output[7]);
  assign mux_399_nl = MUX_s_1_2_2(mux_398_nl, mux_392_nl, fsm_output[6]);
  assign or_478_nl = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b010) | (~ IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0]));
  assign or_476_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b010) | (~ IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0]));
  assign mux_384_nl = MUX_s_1_2_2(or_478_nl, or_476_nl, fsm_output[7]);
  assign or_474_nl = (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b010) | (~ IDX_LOOP_slc_IDX_LOOP_acc_8_itm)
      | (~ (fsm_output[0]));
  assign or_472_nl = (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b010) | (~ IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm)
      | (~ (fsm_output[0]));
  assign mux_383_nl = MUX_s_1_2_2(or_474_nl, or_472_nl, fsm_output[7]);
  assign mux_385_nl = MUX_s_1_2_2(mux_384_nl, mux_383_nl, fsm_output[6]);
  assign mux_400_nl = MUX_s_1_2_2(mux_399_nl, mux_385_nl, fsm_output[5]);
  assign vec_rsc_0_2_i_re_d_pff = (~ mux_400_nl) & and_dcpl_176;
  assign and_313_nl = and_dcpl_200 & and_dcpl_306;
  assign and_315_nl = and_dcpl_97 & (or_dcpl_74 | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1]))
      & and_dcpl_204;
  assign and_318_nl = and_dcpl_311 & and_dcpl_210;
  assign and_320_nl = and_dcpl_313 & and_dcpl_216;
  assign and_324_nl = and_dcpl_200 & and_dcpl_317;
  assign and_326_nl = and_dcpl_319 & and_dcpl_224;
  assign and_329_nl = and_dcpl_322 & and_dcpl_230;
  assign and_331_nl = and_dcpl_324 & and_dcpl_234;
  assign vec_rsc_0_3_i_radr_d = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_tmp[8:2]), IDX_LOOP_idx1_acc_psp_8_sva,
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_155 , and_313_nl , and_315_nl , and_dcpl_207
      , and_318_nl , and_320_nl , and_dcpl_219 , and_324_nl , and_326_nl , and_dcpl_227
      , and_329_nl , and_331_nl});
  assign or_432_nl = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b01) | (~ (fsm_output[7]));
  assign nand_6_nl = ~((reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]) & (~ mux_256_cse));
  assign mux_357_nl = MUX_s_1_2_2(or_432_nl, nand_6_nl, fsm_output[6]);
  assign or_430_nl = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b01) | (fsm_output[7:6]!=2'b00);
  assign mux_358_nl = MUX_s_1_2_2(mux_357_nl, or_430_nl, fsm_output[8]);
  assign nor_151_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | mux_358_nl);
  assign nand_16_nl = ~((fsm_output[7]) & (IDX_LOOP_idx2_9_0_4_sva[2:0]==3'b011));
  assign or_423_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b011);
  assign mux_352_nl = MUX_s_1_2_2(or_425_cse, or_423_nl, fsm_output[7]);
  assign mux_353_nl = MUX_s_1_2_2(nand_16_nl, mux_352_nl, fsm_output[6]);
  assign or_422_nl = (fsm_output[7:6]!=2'b00) | (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b011);
  assign mux_354_nl = MUX_s_1_2_2(mux_353_nl, or_422_nl, fsm_output[8]);
  assign or_419_nl = (IDX_LOOP_idx2_acc_psp_sva[1]) | (~((IDX_LOOP_idx2_acc_psp_sva[0])
      & (STAGE_LOOP_op_rshift_psp_1_sva[0])));
  assign or_418_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b01) | (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign mux_350_nl = MUX_s_1_2_2(or_419_nl, or_418_nl, fsm_output[7]);
  assign or_416_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1]) | (~((IDX_LOOP_idx2_acc_1_psp_sva[0])
      & (STAGE_LOOP_op_rshift_psp_1_sva[0])));
  assign or_415_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b01) | (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign mux_349_nl = MUX_s_1_2_2(or_416_nl, or_415_nl, fsm_output[7]);
  assign mux_351_nl = MUX_s_1_2_2(mux_350_nl, mux_349_nl, fsm_output[6]);
  assign or_420_nl = (fsm_output[8]) | mux_351_nl;
  assign mux_355_nl = MUX_s_1_2_2(mux_354_nl, or_420_nl, fsm_output[5]);
  assign nor_152_nl = ~((fsm_output[1]) | mux_355_nl);
  assign mux_359_nl = MUX_s_1_2_2(nor_151_nl, nor_152_nl, fsm_output[0]);
  assign vec_rsc_0_3_i_we_d_pff = mux_359_nl & and_dcpl_97;
  assign nor_147_nl = ~((IDX_LOOP_idx2_acc_tmp[1:0]!=2'b01) | (fsm_output[0]));
  assign and_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]==2'b01) & IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm
      & (fsm_output[0]);
  assign mux_369_nl = MUX_s_1_2_2(nor_147_nl, and_nl, fsm_output[7]);
  assign and_525_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]==2'b01) & IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm
      & (fsm_output[0]);
  assign and_526_nl = IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm & (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b01)
      & (fsm_output[0]);
  assign mux_368_nl = MUX_s_1_2_2(and_525_nl, and_526_nl, fsm_output[7]);
  assign mux_370_nl = MUX_s_1_2_2(mux_369_nl, mux_368_nl, fsm_output[6]);
  assign nand_7_nl = ~((STAGE_LOOP_op_rshift_psp_1_sva[0]) & mux_370_nl);
  assign or_443_nl = (fsm_output[0]) | (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b011);
  assign and_308_nl = (fsm_output[0]) & or_425_cse;
  assign mux_364_nl = MUX_s_1_2_2((fsm_output[0]), and_308_nl, IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm);
  assign nor_90_nl = ~((reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7!=2'b01));
  assign mux_365_nl = MUX_s_1_2_2(or_443_nl, mux_364_nl, nor_90_nl);
  assign and_460_nl = ((IDX_LOOP_idx1_acc_2_psp_sva[0]) | (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]))
      | (~ IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm)) & (fsm_output[0]);
  assign nor_88_nl = ~((IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b011));
  assign mux_363_nl = MUX_s_1_2_2(or_439_cse, and_460_nl, nor_88_nl);
  assign mux_366_nl = MUX_s_1_2_2(mux_365_nl, mux_363_nl, fsm_output[7]);
  assign and_461_nl = ((IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b01) | (~ IDX_LOOP_slc_IDX_LOOP_acc_8_itm))
      & (fsm_output[0]);
  assign nor_86_nl = ~((IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b011));
  assign mux_361_nl = MUX_s_1_2_2(or_437_cse, and_461_nl, nor_86_nl);
  assign and_462_nl = ((IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b01) | (~ IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm))
      & (fsm_output[0]);
  assign nor_84_nl = ~((IDX_LOOP_idx2_9_0_sva[2:0]!=3'b011));
  assign mux_360_nl = MUX_s_1_2_2(or_435_cse, and_462_nl, nor_84_nl);
  assign mux_362_nl = MUX_s_1_2_2(mux_361_nl, mux_360_nl, fsm_output[7]);
  assign mux_367_nl = MUX_s_1_2_2(mux_366_nl, mux_362_nl, fsm_output[6]);
  assign mux_371_nl = MUX_s_1_2_2(nand_7_nl, mux_367_nl, fsm_output[5]);
  assign vec_rsc_0_3_i_re_d_pff = (~ mux_371_nl) & and_dcpl_176;
  assign and_299_nl = and_dcpl_212 & and_dcpl_293;
  assign and_300_nl = and_dcpl_279 & and_dcpl_252;
  assign and_301_nl = and_dcpl_271 & and_dcpl_256;
  assign and_302_nl = and_dcpl_282 & and_dcpl_259;
  assign and_305_nl = and_dcpl_232 & and_dcpl_299;
  assign and_306_nl = and_dcpl_288 & and_dcpl_265;
  assign vec_rsc_0_4_i_radr_d = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_tmp[8:2]), IDX_LOOP_idx1_acc_psp_8_sva,
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_155 , and_dcpl_158 , and_dcpl_247 ,
      and_299_nl , and_300_nl , and_dcpl_254 , and_301_nl , and_302_nl , and_dcpl_261
      , and_305_nl , and_306_nl , and_dcpl_267});
  assign or_391_nl = (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1])) | (fsm_output[8]);
  assign or_390_nl = (~ (IDX_LOOP_idx1_acc_2_psp_sva[0])) | (fsm_output[8]);
  assign mux_331_nl = MUX_s_1_2_2(or_391_nl, or_390_nl, fsm_output[7]);
  assign nor_155_nl = ~((reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]) | mux_331_nl);
  assign nor_156_nl = ~((IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b10) | (fsm_output[8]));
  assign nor_157_nl = ~((IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b10) | (fsm_output[8]));
  assign mux_330_nl = MUX_s_1_2_2(nor_156_nl, nor_157_nl, fsm_output[7]);
  assign mux_332_nl = MUX_s_1_2_2(nor_155_nl, mux_330_nl, fsm_output[6]);
  assign and_466_nl = (fsm_output[1]) & (fsm_output[5]) & mux_332_nl;
  assign or_386_nl = (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b100) | (~ (fsm_output[8]));
  assign or_384_nl = (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b100) | (fsm_output[8]);
  assign mux_327_nl = MUX_s_1_2_2(or_386_nl, or_384_nl, fsm_output[7]);
  assign or_383_nl = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b100) | (fsm_output[8]);
  assign or_382_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b100) | (fsm_output[8]);
  assign mux_326_nl = MUX_s_1_2_2(or_383_nl, or_382_nl, fsm_output[7]);
  assign mux_328_nl = MUX_s_1_2_2(mux_327_nl, mux_326_nl, fsm_output[6]);
  assign or_381_nl = (IDX_LOOP_idx2_acc_psp_sva[1:0]!=2'b10) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign or_380_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b10) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign mux_324_nl = MUX_s_1_2_2(or_381_nl, or_380_nl, fsm_output[7]);
  assign or_379_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b10) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign or_378_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b10) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign mux_323_nl = MUX_s_1_2_2(or_379_nl, or_378_nl, fsm_output[7]);
  assign mux_325_nl = MUX_s_1_2_2(mux_324_nl, mux_323_nl, fsm_output[6]);
  assign mux_329_nl = MUX_s_1_2_2(mux_328_nl, mux_325_nl, fsm_output[5]);
  assign nor_158_nl = ~((fsm_output[1]) | mux_329_nl);
  assign mux_333_nl = MUX_s_1_2_2(and_466_nl, nor_158_nl, fsm_output[0]);
  assign vec_rsc_0_4_i_we_d_pff = mux_333_nl & and_dcpl_97;
  assign or_413_nl = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7!=2'b10) | (~ (fsm_output[0]));
  assign nor_153_nl = ~((~((IDX_LOOP_idx2_acc_tmp[0]) | (STAGE_LOOP_op_rshift_psp_1_sva[0])))
      | (fsm_output[0]));
  assign or_409_nl = (IDX_LOOP_idx2_acc_tmp[0]) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[0]);
  assign mux_344_nl = MUX_s_1_2_2(nor_153_nl, or_409_nl, or_362_cse);
  assign mux_345_nl = MUX_s_1_2_2(or_413_nl, mux_344_nl, IDX_LOOP_idx2_acc_tmp[1]);
  assign and_463_nl = ((~ IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm) | (STAGE_LOOP_op_rshift_psp_1_sva[0]))
      & (fsm_output[0]);
  assign nor_79_nl = ~((IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b10));
  assign mux_342_nl = MUX_s_1_2_2(or_tmp_248, and_463_nl, nor_79_nl);
  assign or_406_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b10);
  assign mux_343_nl = MUX_s_1_2_2(mux_342_nl, or_dcpl_83, or_406_nl);
  assign mux_346_nl = MUX_s_1_2_2(mux_345_nl, mux_343_nl, fsm_output[6]);
  assign or_405_nl = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b100) | (~ IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0]));
  assign or_403_nl = (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b100) | (~ IDX_LOOP_slc_IDX_LOOP_acc_8_itm)
      | (~ (fsm_output[0]));
  assign mux_341_nl = MUX_s_1_2_2(or_405_nl, or_403_nl, fsm_output[6]);
  assign mux_347_nl = MUX_s_1_2_2(mux_346_nl, mux_341_nl, fsm_output[5]);
  assign and_464_nl = ((~ IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm) | (STAGE_LOOP_op_rshift_psp_1_sva[0]))
      & (fsm_output[0]);
  assign or_399_nl = (~ (IDX_LOOP_idx1_acc_2_psp_sva[0])) | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]);
  assign mux_337_nl = MUX_s_1_2_2(and_464_nl, or_tmp_248, or_399_nl);
  assign nor_77_nl = ~((IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b10));
  assign mux_338_nl = MUX_s_1_2_2(or_dcpl_84, mux_337_nl, nor_77_nl);
  assign or_398_nl = (~ (IDX_LOOP_idx2_acc_3_psp_sva[1])) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[0]);
  assign and_465_nl = ((~ (IDX_LOOP_idx2_acc_3_psp_sva[1])) | (~ IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm)
      | (STAGE_LOOP_op_rshift_psp_1_sva[0])) & (fsm_output[0]);
  assign nor_75_nl = ~((IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b10));
  assign mux_335_nl = MUX_s_1_2_2(or_398_nl, and_465_nl, nor_75_nl);
  assign mux_336_nl = MUX_s_1_2_2(mux_335_nl, or_dcpl_85, IDX_LOOP_idx2_acc_3_psp_sva[0]);
  assign mux_339_nl = MUX_s_1_2_2(mux_338_nl, mux_336_nl, fsm_output[6]);
  assign or_396_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b100) | (~ IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm)
      | (~ (fsm_output[0]));
  assign or_394_nl = (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b100) | (~ IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm)
      | (~ (fsm_output[0]));
  assign mux_334_nl = MUX_s_1_2_2(or_396_nl, or_394_nl, fsm_output[6]);
  assign mux_340_nl = MUX_s_1_2_2(mux_339_nl, mux_334_nl, fsm_output[5]);
  assign mux_348_nl = MUX_s_1_2_2(mux_347_nl, mux_340_nl, fsm_output[7]);
  assign vec_rsc_0_4_i_re_d_pff = (~ mux_348_nl) & and_dcpl_176;
  assign and_277_nl = and_dcpl_271 & and_dcpl_198;
  assign and_279_nl = and_dcpl_97 & (or_dcpl_81 | (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1])))
      & and_dcpl_204;
  assign and_283_nl = and_dcpl_212 & and_dcpl_277;
  assign and_285_nl = and_dcpl_279 & and_dcpl_216;
  assign and_286_nl = and_dcpl_271 & and_dcpl_222;
  assign and_288_nl = and_dcpl_282 & and_dcpl_224;
  assign and_292_nl = and_dcpl_232 & and_dcpl_286;
  assign and_294_nl = and_dcpl_288 & and_dcpl_234;
  assign vec_rsc_0_5_i_radr_d = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_tmp[8:2]), IDX_LOOP_idx1_acc_psp_8_sva,
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_155 , and_277_nl , and_279_nl , and_dcpl_207
      , and_283_nl , and_285_nl , and_dcpl_219 , and_286_nl , and_288_nl , and_dcpl_227
      , and_292_nl , and_294_nl});
  assign or_354_nl = (IDX_LOOP_idx1_acc_psp_3_sva[0]) | (~((IDX_LOOP_idx1_acc_psp_3_sva[1])
      & (fsm_output[7])));
  assign or_353_nl = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]) | (~ mux_256_cse);
  assign mux_308_nl = MUX_s_1_2_2(or_354_nl, or_353_nl, fsm_output[6]);
  assign or_352_nl = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b10) | (fsm_output[7:6]!=2'b00);
  assign mux_309_nl = MUX_s_1_2_2(mux_308_nl, or_352_nl, fsm_output[8]);
  assign nor_163_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | mux_309_nl);
  assign or_349_nl = (~ (fsm_output[7])) | (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b101);
  assign or_346_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b101);
  assign mux_303_nl = MUX_s_1_2_2(or_347_cse, or_346_nl, fsm_output[7]);
  assign mux_304_nl = MUX_s_1_2_2(or_349_nl, mux_303_nl, fsm_output[6]);
  assign or_344_nl = (fsm_output[7:6]!=2'b00) | (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b101);
  assign mux_305_nl = MUX_s_1_2_2(mux_304_nl, or_344_nl, fsm_output[8]);
  assign or_341_nl = (IDX_LOOP_idx2_acc_psp_sva[1:0]!=2'b10) | (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign or_339_nl = (IDX_LOOP_idx2_acc_2_psp_sva[0]) | (~((IDX_LOOP_idx2_acc_2_psp_sva[1])
      & (STAGE_LOOP_op_rshift_psp_1_sva[0])));
  assign mux_301_nl = MUX_s_1_2_2(or_341_nl, or_339_nl, fsm_output[7]);
  assign or_338_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b10) | (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign or_336_nl = (IDX_LOOP_idx2_acc_3_psp_sva[0]) | (~((IDX_LOOP_idx2_acc_3_psp_sva[1])
      & (STAGE_LOOP_op_rshift_psp_1_sva[0])));
  assign mux_300_nl = MUX_s_1_2_2(or_338_nl, or_336_nl, fsm_output[7]);
  assign mux_302_nl = MUX_s_1_2_2(mux_301_nl, mux_300_nl, fsm_output[6]);
  assign or_342_nl = (fsm_output[8]) | mux_302_nl;
  assign mux_306_nl = MUX_s_1_2_2(mux_305_nl, or_342_nl, fsm_output[5]);
  assign nor_164_nl = ~((fsm_output[1]) | mux_306_nl);
  assign mux_310_nl = MUX_s_1_2_2(nor_163_nl, nor_164_nl, fsm_output[0]);
  assign vec_rsc_0_5_i_we_d_pff = mux_310_nl & and_dcpl_97;
  assign nor_159_nl = ~((IDX_LOOP_idx2_acc_tmp[1:0]!=2'b10) | (fsm_output[0]));
  assign and_522_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]==2'b10) & IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm
      & (fsm_output[0]);
  assign mux_320_nl = MUX_s_1_2_2(nor_159_nl, and_522_nl, fsm_output[7]);
  assign and_523_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]==2'b10) & IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm
      & (fsm_output[0]);
  assign and_524_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b10) & IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm
      & (fsm_output[0]);
  assign mux_319_nl = MUX_s_1_2_2(and_523_nl, and_524_nl, fsm_output[7]);
  assign mux_321_nl = MUX_s_1_2_2(mux_320_nl, mux_319_nl, fsm_output[6]);
  assign nand_4_nl = ~((STAGE_LOOP_op_rshift_psp_1_sva[0]) & mux_321_nl);
  assign and_273_nl = (fsm_output[0]) & or_347_cse;
  assign mux_315_nl = MUX_s_1_2_2((fsm_output[0]), and_273_nl, IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm);
  assign or_364_nl = (fsm_output[0]) | (IDX_LOOP_idx2_9_0_2_sva[1]) | nand_23_cse;
  assign mux_316_nl = MUX_s_1_2_2(mux_315_nl, or_364_nl, or_362_cse);
  assign or_361_nl = (~ (IDX_LOOP_idx1_acc_2_psp_sva[0])) | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0])
      | (fsm_output[0]);
  assign and_467_nl = ((~ (IDX_LOOP_idx1_acc_2_psp_sva[0])) | (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0])
      | (~ IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm)) & (fsm_output[0]);
  assign nor_71_nl = ~((IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b101));
  assign mux_314_nl = MUX_s_1_2_2(or_361_nl, and_467_nl, nor_71_nl);
  assign mux_317_nl = MUX_s_1_2_2(mux_316_nl, mux_314_nl, fsm_output[7]);
  assign or_359_nl = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b10) | (fsm_output[0]);
  assign and_468_nl = ((IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b10) | (~ IDX_LOOP_slc_IDX_LOOP_acc_8_itm))
      & (fsm_output[0]);
  assign nor_69_nl = ~((IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b101));
  assign mux_312_nl = MUX_s_1_2_2(or_359_nl, and_468_nl, nor_69_nl);
  assign or_357_nl = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b10) | (fsm_output[0]);
  assign and_469_nl = ((IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b10) | (~ IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm))
      & (fsm_output[0]);
  assign nor_67_nl = ~((IDX_LOOP_idx2_9_0_sva[2:0]!=3'b101));
  assign mux_311_nl = MUX_s_1_2_2(or_357_nl, and_469_nl, nor_67_nl);
  assign mux_313_nl = MUX_s_1_2_2(mux_312_nl, mux_311_nl, fsm_output[7]);
  assign mux_318_nl = MUX_s_1_2_2(mux_317_nl, mux_313_nl, fsm_output[6]);
  assign mux_322_nl = MUX_s_1_2_2(nand_4_nl, mux_318_nl, fsm_output[5]);
  assign vec_rsc_0_5_i_re_d_pff = (~ mux_322_nl) & and_dcpl_176;
  assign and_254_nl = and_dcpl_212 & and_dcpl_249;
  assign and_257_nl = and_dcpl_217 & and_dcpl_252;
  assign and_261_nl = and_dcpl_200 & and_dcpl_256;
  assign and_264_nl = and_dcpl_225 & and_dcpl_259;
  assign and_268_nl = and_dcpl_232 & and_dcpl_263;
  assign and_270_nl = and_dcpl_235 & and_dcpl_265;
  assign vec_rsc_0_6_i_radr_d = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_tmp[8:2]), IDX_LOOP_idx1_acc_psp_8_sva,
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_155 , and_dcpl_158 , and_dcpl_247 ,
      and_254_nl , and_257_nl , and_dcpl_254 , and_261_nl , and_264_nl , and_dcpl_261
      , and_268_nl , and_270_nl , and_dcpl_267});
  assign nor_167_nl = ~((~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1])) | (fsm_output[8]));
  assign nor_168_nl = ~((~ (IDX_LOOP_idx1_acc_2_psp_sva[0])) | (fsm_output[8]));
  assign mux_280_nl = MUX_s_1_2_2(nor_167_nl, nor_168_nl, fsm_output[7]);
  assign and_479_nl = (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]) & mux_280_nl;
  assign nor_169_nl = ~((IDX_LOOP_idx1_acc_psp_3_sva[1:0]!=2'b11) | (fsm_output[8]));
  assign nor_170_nl = ~((IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b11) | (fsm_output[8]));
  assign mux_279_nl = MUX_s_1_2_2(nor_169_nl, nor_170_nl, fsm_output[7]);
  assign mux_281_nl = MUX_s_1_2_2(and_479_nl, mux_279_nl, fsm_output[6]);
  assign and_478_nl = (fsm_output[1]) & (fsm_output[5]) & mux_281_nl;
  assign nand_31_nl = ~((IDX_LOOP_idx2_9_0_sva[2:0]==3'b110) & (fsm_output[8]));
  assign or_313_nl = (IDX_LOOP_idx2_9_0_4_sva[2:0]!=3'b110) | (fsm_output[8]);
  assign mux_276_nl = MUX_s_1_2_2(nand_31_nl, or_313_nl, fsm_output[7]);
  assign or_312_nl = (IDX_LOOP_idx2_9_0_2_sva[2:0]!=3'b110) | (fsm_output[8]);
  assign or_311_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]!=3'b110) | (fsm_output[8]);
  assign mux_275_nl = MUX_s_1_2_2(or_312_nl, or_311_nl, fsm_output[7]);
  assign mux_277_nl = MUX_s_1_2_2(mux_276_nl, mux_275_nl, fsm_output[6]);
  assign or_310_nl = (IDX_LOOP_idx2_acc_psp_sva[1:0]!=2'b11) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign or_309_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]!=2'b11) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign mux_273_nl = MUX_s_1_2_2(or_310_nl, or_309_nl, fsm_output[7]);
  assign or_308_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]!=2'b11) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign or_307_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]!=2'b11) | (STAGE_LOOP_op_rshift_psp_1_sva[0])
      | (fsm_output[8]);
  assign mux_272_nl = MUX_s_1_2_2(or_308_nl, or_307_nl, fsm_output[7]);
  assign mux_274_nl = MUX_s_1_2_2(mux_273_nl, mux_272_nl, fsm_output[6]);
  assign mux_278_nl = MUX_s_1_2_2(mux_277_nl, mux_274_nl, fsm_output[5]);
  assign nor_171_nl = ~((fsm_output[1]) | mux_278_nl);
  assign mux_282_nl = MUX_s_1_2_2(and_478_nl, nor_171_nl, fsm_output[0]);
  assign vec_rsc_0_6_i_we_d_pff = mux_282_nl & and_dcpl_97;
  assign or_674_nl = (fsm_output[0]) | (IDX_LOOP_idx2_acc_tmp[1:0]!=2'b11) | (STAGE_LOOP_op_rshift_psp_1_sva[0]);
  assign nor_165_nl = ~((fsm_output[0]) | (~((IDX_LOOP_idx2_acc_tmp[1:0]!=2'b11)
      | (STAGE_LOOP_op_rshift_psp_1_sva[0]))));
  assign mux_296_nl = MUX_s_1_2_2(or_674_nl, nor_165_nl, and_481_cse);
  assign and_471_nl = (IDX_LOOP_idx1_acc_2_psp_sva[0]) & (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]);
  assign mux_294_nl = MUX_s_1_2_2(or_tmp_248, mux_293_cse, and_471_nl);
  assign and_472_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]==2'b11);
  assign mux_295_nl = MUX_s_1_2_2(or_290_cse, mux_294_nl, and_472_nl);
  assign mux_297_nl = MUX_s_1_2_2(mux_296_nl, mux_295_nl, fsm_output[7]);
  assign and_473_nl = (IDX_LOOP_idx1_acc_psp_3_sva[1:0]==2'b11);
  assign mux_290_nl = MUX_s_1_2_2(or_tmp_248, mux_289_cse, and_473_nl);
  assign and_474_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]==2'b11);
  assign mux_291_nl = MUX_s_1_2_2(or_288_cse, mux_290_nl, and_474_nl);
  assign and_475_nl = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]==2'b11);
  assign mux_287_nl = MUX_s_1_2_2(or_tmp_248, mux_286_cse, and_475_nl);
  assign and_476_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11);
  assign mux_288_nl = MUX_s_1_2_2(or_286_cse, mux_287_nl, and_476_nl);
  assign mux_292_nl = MUX_s_1_2_2(mux_291_nl, mux_288_nl, fsm_output[7]);
  assign mux_298_nl = MUX_s_1_2_2(mux_297_nl, mux_292_nl, fsm_output[6]);
  assign nand_68_nl = ~((IDX_LOOP_idx2_9_0_2_sva[2:0]==3'b110) & IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm
      & (fsm_output[0]));
  assign nand_69_nl = ~((IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b110) & IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm
      & (fsm_output[0]));
  assign mux_284_nl = MUX_s_1_2_2(nand_68_nl, nand_69_nl, fsm_output[7]);
  assign nand_67_nl = ~((IDX_LOOP_idx2_9_0_4_sva[2:0]==3'b110) & IDX_LOOP_slc_IDX_LOOP_acc_8_itm
      & (fsm_output[0]));
  assign nand_66_nl = ~((IDX_LOOP_idx2_9_0_sva[2:0]==3'b110) & IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm
      & (fsm_output[0]));
  assign mux_283_nl = MUX_s_1_2_2(nand_67_nl, nand_66_nl, fsm_output[7]);
  assign mux_285_nl = MUX_s_1_2_2(mux_284_nl, mux_283_nl, fsm_output[6]);
  assign mux_299_nl = MUX_s_1_2_2(mux_298_nl, mux_285_nl, fsm_output[5]);
  assign vec_rsc_0_6_i_re_d_pff = (~ mux_299_nl) & and_dcpl_176;
  assign and_205_nl = and_dcpl_200 & and_dcpl_198;
  assign and_210_nl = and_dcpl_97 & (or_dcpl_74 | (~ (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[1])))
      & and_dcpl_204;
  assign and_217_nl = and_dcpl_212 & and_dcpl_210;
  assign and_222_nl = and_dcpl_217 & and_dcpl_216;
  assign and_227_nl = and_dcpl_200 & and_dcpl_222;
  assign and_230_nl = and_dcpl_225 & and_dcpl_224;
  assign and_237_nl = and_dcpl_232 & and_dcpl_230;
  assign and_240_nl = and_dcpl_235 & and_dcpl_234;
  assign vec_rsc_0_7_i_radr_d = MUX1HOT_v_7_12_2((IDX_LOOP_idx2_acc_tmp[8:2]), IDX_LOOP_idx1_acc_psp_8_sva,
      (IDX_LOOP_idx2_9_0_2_sva[9:3]), (IDX_LOOP_idx2_acc_1_psp_sva[8:2]), (IDX_LOOP_idx1_acc_psp_3_sva[8:2]),
      (IDX_LOOP_idx2_9_0_4_sva[9:3]), (IDX_LOOP_idx2_acc_2_psp_sva[8:2]), (IDX_LOOP_idx1_acc_2_psp_sva[7:1]),
      (IDX_LOOP_idx2_9_0_6_sva[9:3]), (IDX_LOOP_idx2_acc_3_psp_sva[8:2]), (IDX_LOOP_idx1_acc_psp_7_sva[8:2]),
      (IDX_LOOP_idx2_9_0_sva[9:3]), {and_dcpl_155 , and_205_nl , and_210_nl , and_dcpl_207
      , and_217_nl , and_222_nl , and_dcpl_219 , and_227_nl , and_230_nl , and_dcpl_227
      , and_237_nl , and_240_nl});
  assign nand_41_nl = ~((IDX_LOOP_idx1_acc_psp_3_sva[1:0]==2'b11) & (fsm_output[7]));
  assign nand_42_nl = ~((reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0]) & mux_256_cse);
  assign mux_257_nl = MUX_s_1_2_2(nand_41_nl, nand_42_nl, fsm_output[6]);
  assign or_283_nl = (IDX_LOOP_idx1_acc_psp_7_sva[1:0]!=2'b11) | (fsm_output[7:6]!=2'b00);
  assign mux_258_nl = MUX_s_1_2_2(mux_257_nl, or_283_nl, fsm_output[8]);
  assign nor_172_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | mux_258_nl);
  assign nand_43_nl = ~((fsm_output[7]) & (IDX_LOOP_idx2_9_0_4_sva[2:0]==3'b111));
  assign nand_45_nl = ~((IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b111));
  assign mux_252_nl = MUX_s_1_2_2(nand_44_cse, nand_45_nl, fsm_output[7]);
  assign mux_253_nl = MUX_s_1_2_2(nand_43_nl, mux_252_nl, fsm_output[6]);
  assign or_280_nl = (fsm_output[7:6]!=2'b00) | (IDX_LOOP_idx2_9_0_sva[2:0]!=3'b111);
  assign mux_254_nl = MUX_s_1_2_2(mux_253_nl, or_280_nl, fsm_output[8]);
  assign nand_47_nl = ~((IDX_LOOP_idx2_acc_psp_sva[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign nand_48_nl = ~((IDX_LOOP_idx2_acc_2_psp_sva[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign mux_250_nl = MUX_s_1_2_2(nand_47_nl, nand_48_nl, fsm_output[7]);
  assign nand_49_nl = ~((IDX_LOOP_idx2_acc_1_psp_sva[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign nand_50_nl = ~((IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0]));
  assign mux_249_nl = MUX_s_1_2_2(nand_49_nl, nand_50_nl, fsm_output[7]);
  assign mux_251_nl = MUX_s_1_2_2(mux_250_nl, mux_249_nl, fsm_output[6]);
  assign or_278_nl = (fsm_output[8]) | mux_251_nl;
  assign mux_255_nl = MUX_s_1_2_2(mux_254_nl, or_278_nl, fsm_output[5]);
  assign nor_173_nl = ~((fsm_output[1]) | mux_255_nl);
  assign mux_259_nl = MUX_s_1_2_2(nor_172_nl, nor_173_nl, fsm_output[0]);
  assign vec_rsc_0_7_i_we_d_pff = mux_259_nl & and_dcpl_97;
  assign nand_32_nl = ~((IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (fsm_output[0])));
  assign or_297_nl = (~((IDX_LOOP_idx2_acc_2_psp_sva[1:0]==2'b11) & IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm))
      | not_tmp_180;
  assign mux_269_nl = MUX_s_1_2_2(nand_32_nl, or_297_nl, fsm_output[7]);
  assign or_295_nl = (~((IDX_LOOP_idx2_acc_1_psp_sva[1:0]==2'b11) & IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm))
      | not_tmp_180;
  assign or_293_nl = (~((IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11) & IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm))
      | not_tmp_180;
  assign mux_268_nl = MUX_s_1_2_2(or_295_nl, or_293_nl, fsm_output[7]);
  assign mux_270_nl = MUX_s_1_2_2(mux_269_nl, mux_268_nl, fsm_output[6]);
  assign or_291_nl = (fsm_output[0]) | nand_44_cse;
  assign and_480_nl = (fsm_output[0]) & nand_44_cse;
  assign mux_264_nl = MUX_s_1_2_2((fsm_output[0]), and_480_nl, IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm);
  assign mux_265_nl = MUX_s_1_2_2(or_291_nl, mux_264_nl, and_481_cse);
  assign and_482_nl = (~((IDX_LOOP_idx1_acc_2_psp_sva[0]) & (reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7[0])
      & IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm)) & (fsm_output[0]);
  assign and_483_nl = (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b111);
  assign mux_263_nl = MUX_s_1_2_2(or_290_cse, and_482_nl, and_483_nl);
  assign mux_266_nl = MUX_s_1_2_2(mux_265_nl, mux_263_nl, fsm_output[7]);
  assign and_484_nl = (~((IDX_LOOP_idx1_acc_psp_3_sva[1:0]==2'b11) & IDX_LOOP_slc_IDX_LOOP_acc_8_itm))
      & (fsm_output[0]);
  assign and_485_nl = (IDX_LOOP_idx2_9_0_4_sva[2:0]==3'b111);
  assign mux_261_nl = MUX_s_1_2_2(or_288_cse, and_484_nl, and_485_nl);
  assign and_486_nl = (~((IDX_LOOP_idx1_acc_psp_7_sva[1:0]==2'b11) & IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm))
      & (fsm_output[0]);
  assign and_487_nl = (IDX_LOOP_idx2_9_0_sva[2:0]==3'b111);
  assign mux_260_nl = MUX_s_1_2_2(or_286_cse, and_486_nl, and_487_nl);
  assign mux_262_nl = MUX_s_1_2_2(mux_261_nl, mux_260_nl, fsm_output[7]);
  assign mux_267_nl = MUX_s_1_2_2(mux_266_nl, mux_262_nl, fsm_output[6]);
  assign mux_271_nl = MUX_s_1_2_2(mux_270_nl, mux_267_nl, fsm_output[5]);
  assign vec_rsc_0_7_i_re_d_pff = (~ mux_271_nl) & and_dcpl_176;
  assign twiddle_rsc_0_0_i_radr_d_pff = z_out_6[9:3];
  assign nor_175_cse = ~((z_out_6[2:0]!=3'b000) | (fsm_output[3]));
  assign nor_174_nl = ~((z_out_6[2:0]!=3'b000) | (~ (fsm_output[3])));
  assign mux_246_nl = MUX_s_1_2_2(nor_174_nl, nor_175_cse, fsm_output[2]);
  assign mux_247_nl = MUX_s_1_2_2(mux_246_nl, nor_175_cse, fsm_output[1]);
  assign twiddle_rsc_0_0_i_re_d_pff = mux_247_nl & and_dcpl_151;
  assign nor_183_cse = ~((z_out_6[2:0]!=3'b001) | (fsm_output[3]));
  assign nor_182_nl = ~((z_out_6[2:0]!=3'b001) | (~ (fsm_output[3])));
  assign mux_239_nl = MUX_s_1_2_2(nor_182_nl, nor_183_cse, fsm_output[2]);
  assign mux_240_nl = MUX_s_1_2_2(mux_239_nl, nor_183_cse, fsm_output[1]);
  assign nor_186_nl = ~((z_out_6[2:1]!=2'b00) | not_tmp_164);
  assign mux_236_nl = MUX_s_1_2_2(nor_186_nl, nor_183_cse, fsm_output[2]);
  assign mux_237_nl = MUX_s_1_2_2(mux_236_nl, nor_183_cse, fsm_output[1]);
  assign mux_241_nl = MUX_s_1_2_2(mux_240_nl, mux_237_nl, fsm_output[0]);
  assign twiddle_rsc_0_1_i_re_d_pff = mux_241_nl & and_dcpl_151;
  assign nor_191_cse = ~((z_out_6[2:0]!=3'b010) | (fsm_output[3]));
  assign nor_190_nl = ~((z_out_6[2]) | (z_out_6[0]) | not_tmp_162);
  assign mux_232_nl = MUX_s_1_2_2(nor_190_nl, nor_191_cse, fsm_output[2]);
  assign mux_233_nl = MUX_s_1_2_2(mux_232_nl, nor_191_cse, fsm_output[1]);
  assign nor_194_nl = ~((z_out_6[2:0]!=3'b010) | (~ (fsm_output[3])));
  assign mux_229_nl = MUX_s_1_2_2(nor_194_nl, nor_191_cse, fsm_output[2]);
  assign mux_230_nl = MUX_s_1_2_2(mux_229_nl, nor_191_cse, fsm_output[1]);
  assign mux_234_nl = MUX_s_1_2_2(mux_233_nl, mux_230_nl, fsm_output[0]);
  assign twiddle_rsc_0_2_i_re_d_pff = mux_234_nl & and_dcpl_151;
  assign nor_199_cse = ~((z_out_6[2:0]!=3'b011) | (fsm_output[3]));
  assign nor_198_nl = ~((z_out_6[2]) | (~((z_out_6[1:0]==2'b11) & (fsm_output[3]))));
  assign mux_225_nl = MUX_s_1_2_2(nor_198_nl, nor_199_cse, fsm_output[2]);
  assign mux_226_nl = MUX_s_1_2_2(mux_225_nl, nor_199_cse, fsm_output[1]);
  assign twiddle_rsc_0_3_i_re_d_pff = mux_226_nl & and_dcpl_151;
  assign nor_207_cse = ~((z_out_6[2:0]!=3'b100) | (fsm_output[3]));
  assign nor_206_nl = ~((z_out_6[2:0]!=3'b100) | (~ (fsm_output[3])));
  assign mux_218_nl = MUX_s_1_2_2(nor_206_nl, nor_207_cse, fsm_output[2]);
  assign mux_219_nl = MUX_s_1_2_2(mux_218_nl, nor_207_cse, fsm_output[1]);
  assign twiddle_rsc_0_4_i_re_d_pff = mux_219_nl & and_dcpl_151;
  assign nor_215_cse = ~((z_out_6[2:0]!=3'b101) | (fsm_output[3]));
  assign and_520_nl = (z_out_6[2:0]==3'b101) & (fsm_output[3]);
  assign mux_211_nl = MUX_s_1_2_2(and_520_nl, nor_215_cse, fsm_output[2]);
  assign mux_212_nl = MUX_s_1_2_2(mux_211_nl, nor_215_cse, fsm_output[1]);
  assign nor_218_nl = ~((z_out_6[2:1]!=2'b10) | not_tmp_164);
  assign mux_208_nl = MUX_s_1_2_2(nor_218_nl, nor_215_cse, fsm_output[2]);
  assign mux_209_nl = MUX_s_1_2_2(mux_208_nl, nor_215_cse, fsm_output[1]);
  assign mux_213_nl = MUX_s_1_2_2(mux_212_nl, mux_209_nl, fsm_output[0]);
  assign twiddle_rsc_0_5_i_re_d_pff = mux_213_nl & and_dcpl_151;
  assign nor_223_cse = ~((z_out_6[2:0]!=3'b110) | (fsm_output[3]));
  assign nor_222_nl = ~((~ (z_out_6[2])) | (z_out_6[0]) | not_tmp_162);
  assign mux_204_nl = MUX_s_1_2_2(nor_222_nl, nor_223_cse, fsm_output[2]);
  assign mux_205_nl = MUX_s_1_2_2(mux_204_nl, nor_223_cse, fsm_output[1]);
  assign and_519_nl = (z_out_6[2:0]==3'b110) & (fsm_output[3]);
  assign mux_201_nl = MUX_s_1_2_2(and_519_nl, nor_223_cse, fsm_output[2]);
  assign mux_202_nl = MUX_s_1_2_2(mux_201_nl, nor_223_cse, fsm_output[1]);
  assign mux_206_nl = MUX_s_1_2_2(mux_205_nl, mux_202_nl, fsm_output[0]);
  assign twiddle_rsc_0_6_i_re_d_pff = mux_206_nl & and_dcpl_151;
  assign and_489_cse = (z_out_6[2:0]==3'b111) & (~ (fsm_output[3]));
  assign and_488_nl = (z_out_6[2:0]==3'b111) & (fsm_output[3]);
  assign mux_197_nl = MUX_s_1_2_2(and_488_nl, and_489_cse, fsm_output[2]);
  assign mux_198_nl = MUX_s_1_2_2(mux_197_nl, and_489_cse, fsm_output[1]);
  assign twiddle_rsc_0_7_i_re_d_pff = mux_198_nl & and_dcpl_151;
  assign and_dcpl_431 = ~((fsm_output[5]) | (fsm_output[7]));
  assign and_dcpl_436 = ~((fsm_output[0]) | (fsm_output[4]) | (fsm_output[3]));
  assign and_dcpl_443 = and_dcpl_436 & (fsm_output[2]) & (~ (fsm_output[1])) & (~
      (fsm_output[6])) & (fsm_output[8]) & and_dcpl_431;
  assign nor_327_cse = ~((fsm_output[6]) | (fsm_output[8]));
  assign nor_326_cse = ~((fsm_output[4:2]!=3'b000));
  assign and_dcpl_454 = nor_326_cse & (fsm_output[1:0]==2'b10) & nor_327_cse & and_dcpl_431;
  assign and_dcpl_468 = and_dcpl_96 & (fsm_output[2]) & (~ (fsm_output[1])) & (~
      (fsm_output[0])) & (~ (fsm_output[6])) & (fsm_output[8]) & and_dcpl_431;
  assign and_dcpl_469 = (fsm_output[5]) & (~ (fsm_output[7]));
  assign and_dcpl_475 = nor_326_cse & (fsm_output[1:0]==2'b11);
  assign and_dcpl_476 = and_dcpl_475 & nor_327_cse & and_dcpl_469;
  assign and_dcpl_477 = (fsm_output[6]) & (~ (fsm_output[8]));
  assign and_dcpl_479 = and_dcpl_475 & and_dcpl_477 & and_dcpl_469;
  assign and_dcpl_480 = (fsm_output[5]) & (fsm_output[7]);
  assign and_dcpl_482 = and_dcpl_475 & nor_327_cse & and_dcpl_480;
  assign and_dcpl_484 = and_dcpl_475 & and_dcpl_477 & and_dcpl_480;
  assign and_dcpl_491 = and_dcpl_96 & (fsm_output[2:0]==3'b011);
  assign and_dcpl_492 = and_dcpl_491 & and_dcpl_477 & and_dcpl_431;
  assign and_dcpl_493 = (~ (fsm_output[5])) & (fsm_output[7]);
  assign and_dcpl_496 = and_dcpl_491 & nor_327_cse & and_dcpl_493;
  assign and_dcpl_498 = and_dcpl_491 & and_dcpl_477 & and_dcpl_493;
  assign and_dcpl_503 = and_dcpl_96 & (fsm_output[2]) & and_dcpl_95 & nor_327_cse
      & and_dcpl_431;
  assign and_dcpl_509 = ~((fsm_output[4:0]!=5'b01000));
  assign and_dcpl_533 = (fsm_output[4:0]==5'b00010) & nor_327_cse & and_dcpl_431;
  assign and_dcpl_536 = nor_327_cse & and_dcpl_431;
  assign and_dcpl_544 = and_dcpl_97 & and_dcpl_153 & and_dcpl_536;
  assign and_dcpl_547 = and_dcpl_97 & and_509_cse & and_dcpl_536;
  assign and_dcpl_551 = and_dcpl_103 & and_dcpl_95 & and_dcpl_536;
  assign and_dcpl_553 = and_dcpl_103 & and_dcpl_102 & and_dcpl_536;
  assign and_dcpl_555 = and_dcpl_103 & and_dcpl_153 & and_dcpl_536;
  assign and_dcpl_557 = and_dcpl_103 & and_509_cse & and_dcpl_536;
  assign and_dcpl_559 = (fsm_output[4:2]==3'b010);
  assign and_dcpl_561 = and_dcpl_559 & and_dcpl_95 & and_dcpl_536;
  assign and_dcpl_563 = and_dcpl_559 & and_dcpl_102 & and_dcpl_536;
  assign and_dcpl_570 = and_dcpl_96 & (fsm_output[2]) & and_dcpl_95;
  assign and_dcpl_571 = and_dcpl_570 & nor_327_cse & and_dcpl_469;
  assign and_dcpl_574 = and_dcpl_570 & and_dcpl_477 & and_dcpl_469;
  assign and_dcpl_577 = and_dcpl_570 & nor_327_cse & and_dcpl_480;
  assign and_dcpl_579 = and_dcpl_570 & and_dcpl_477 & and_dcpl_480;
  assign and_dcpl_587 = and_dcpl_570 & and_dcpl_477 & (~ (fsm_output[5])) & (~ (fsm_output[7]));
  assign and_dcpl_591 = and_dcpl_570 & (~ (fsm_output[6])) & (~ (fsm_output[8]))
      & and_dcpl_493;
  assign and_dcpl_593 = and_dcpl_570 & and_dcpl_477 & and_dcpl_493;
  assign and_dcpl_600 = and_dcpl_103 & (fsm_output[1:0]==2'b00);
  assign and_dcpl_601 = and_dcpl_600 & nor_327_cse & and_dcpl_431;
  assign and_dcpl_604 = and_dcpl_103 & (~ (fsm_output[1])) & (fsm_output[0]) & (~
      (fsm_output[8]));
  assign and_dcpl_607 = and_dcpl_600 & nor_327_cse & and_dcpl_469;
  assign and_dcpl_610 = and_dcpl_600 & and_dcpl_477 & and_dcpl_431;
  assign and_dcpl_612 = and_dcpl_600 & and_dcpl_477 & and_dcpl_469;
  assign and_dcpl_615 = and_dcpl_600 & nor_327_cse & and_dcpl_493;
  assign and_dcpl_618 = and_dcpl_600 & nor_327_cse & and_dcpl_480;
  assign and_dcpl_620 = and_dcpl_600 & and_dcpl_477 & and_dcpl_493;
  assign and_dcpl_622 = and_dcpl_600 & and_dcpl_477 & and_dcpl_480;
  assign and_636_ssc = and_dcpl_97 & and_dcpl_102 & and_dcpl_536;
  assign or_tmp = (fsm_output[8:5]!=4'b0111);
  assign or_698_nl = (fsm_output[6:5]!=2'b00);
  assign nand_71_nl = ~((fsm_output[6:5]==2'b11));
  assign mux_nl = MUX_s_1_2_2(or_698_nl, nand_71_nl, fsm_output[7]);
  assign or_tmp_545 = (fsm_output[8]) | mux_nl;
  always @(posedge clk) begin
    if ( rst ) begin
      STAGE_LOOP_i_3_0_sva <= 4'b0000;
    end
    else if ( (and_dcpl_97 & and_dcpl_95 & and_dcpl_94) | STAGE_LOOP_i_3_0_sva_mx0c1
        ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, STAGE_LOOP_i_3_0_sva_2, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      p_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ mux_187_nl ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_IDX_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      reg_ensig_cgo_cse <= 1'b0;
      IDX_LOOP_1_IDX_LOOP_rem_1_cmp_a <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      reg_twiddle_rsc_triosy_0_0_obj_ld_cse <= 1'b0;
      IDX_LOOP_IDX_LOOP_and_106_itm <= 1'b0;
      IDX_LOOP_IDX_LOOP_and_107_itm <= 1'b0;
      IDX_LOOP_IDX_LOOP_and_108_itm <= 1'b0;
      IDX_LOOP_IDX_LOOP_nor_12_itm <= 1'b0;
      reg_cse <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      reg_1_cse <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      reg_2_cse <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tmp_11_sva_29 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tmp_11_sva_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tmp_11_sva_5 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tmp_11_sva_7 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      tmp_11_sva_9 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      reg_IDX_LOOP_1_lshift_idiv_ftd_7 <= 3'b000;
    end
    else begin
      reg_IDX_LOOP_1_modulo_dev_cmp_m_rsc_dat_cse <= p_sva;
      reg_ensig_cgo_cse <= nor_302_rmff;
      IDX_LOOP_1_IDX_LOOP_rem_1_cmp_a <= MUX_v_128_2_2(IDX_LOOP_1_mul_mut, z_out_5,
          mux_192_nl);
      reg_twiddle_rsc_triosy_0_0_obj_ld_cse <= and_dcpl_104 & and_dcpl_93 & (fsm_output[8:7]==2'b10)
          & STAGE_LOOP_acc_itm_4_1;
      IDX_LOOP_IDX_LOOP_and_106_itm <= (z_out_6[2:0]==3'b101);
      IDX_LOOP_IDX_LOOP_and_107_itm <= (z_out_6[2:0]==3'b110);
      IDX_LOOP_IDX_LOOP_and_108_itm <= (z_out_6[2:0]==3'b111);
      IDX_LOOP_IDX_LOOP_nor_12_itm <= ~((z_out_6[2:0]!=3'b000));
      reg_cse <= MUX_v_64_2_2(vec_rsc_0_7_i_q_d, vec_rsc_0_6_i_q_d, and_dcpl_430);
      reg_1_cse <= MUX_v_64_2_2(vec_rsc_0_1_i_q_d, vec_rsc_0_0_i_q_d, and_dcpl_430);
      reg_2_cse <= MUX1HOT_v_64_3_2(vec_rsc_0_3_i_q_d, vec_rsc_0_2_i_q_d, vec_rsc_0_4_i_q_d,
          {and_dcpl_413 , IDX_LOOP_f2_or_5_nl , IDX_LOOP_f2_or_6_nl});
      tmp_11_sva_29 <= MUX_v_64_2_2(vec_rsc_0_5_i_q_d, vec_rsc_0_6_i_q_d, and_dcpl_430);
      tmp_11_sva_3 <= MUX_v_64_2_2(vec_rsc_0_3_i_q_d, vec_rsc_0_0_i_q_d, and_dcpl_430);
      tmp_11_sva_5 <= vec_rsc_0_5_i_q_d;
      tmp_11_sva_7 <= vec_rsc_0_7_i_q_d;
      tmp_11_sva_9 <= vec_rsc_0_1_i_q_d;
      reg_IDX_LOOP_1_lshift_idiv_ftd_7 <= z_out_6[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      STAGE_LOOP_op_rshift_psp_1_sva <= 10'b0000000000;
    end
    else if ( ~ mux_180_cse ) begin
      STAGE_LOOP_op_rshift_psp_1_sva <= STAGE_LOOP_op_rshift_itm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      STAGE_LOOP_gp_lshift_psp_sva <= 10'b0000000000;
    end
    else if ( ~ mux_180_cse ) begin
      STAGE_LOOP_gp_lshift_psp_sva <= z_out_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      GROUP_LOOP_j_10_0_sva_9_0 <= 10'b0000000000;
    end
    else if ( GROUP_LOOP_j_10_0_sva_9_0_mx0c0 | (and_dcpl_108 & and_dcpl_101) ) begin
      GROUP_LOOP_j_10_0_sva_9_0 <= MUX_v_10_2_2(10'b0000000000, (z_out[9:0]), GROUP_LOOP_j_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_t_10_3_sva_6_0 <= 7'b0000000;
    end
    else if ( MUX_s_1_2_2(mux_532_nl, or_tmp, fsm_output[4]) ) begin
      IDX_LOOP_t_10_3_sva_6_0 <= MUX_v_7_2_2(7'b0000000, reg_IDX_LOOP_t_10_3_ftd_1,
          or_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      STAGE_LOOP_gp_acc_psp_sva <= 4'b0000;
    end
    else if ( ~ mux_180_cse ) begin
      STAGE_LOOP_gp_acc_psp_sva <= z_out_1[3:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx2_acc_psp_sva <= 9'b000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      IDX_LOOP_idx2_acc_psp_sva <= IDX_LOOP_idx2_acc_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx1_acc_psp_8_sva <= 7'b0000000;
    end
    else if ( ~((~ mux_459_nl) & and_dcpl) ) begin
      IDX_LOOP_idx1_acc_psp_8_sva <= IDX_LOOP_idx1_acc_psp_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx2_9_0_2_sva <= 10'b0000000000;
    end
    else if ( ~((~ mux_461_nl) & and_dcpl) ) begin
      IDX_LOOP_idx2_9_0_2_sva <= IDX_LOOP_idx2_9_0_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      IDX_LOOP_2_slc_IDX_LOOP_acc_10_itm <= z_out[10];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_equal_tmp <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f1_equal_tmp <= IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_equal_tmp_1 <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f1_equal_tmp_1 <= IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_equal_tmp_2 <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f1_equal_tmp_2 <= IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_equal_tmp_3 <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f1_equal_tmp_3 <= IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx2_acc_1_psp_sva <= 9'b000000000;
    end
    else if ( ~(mux_465_nl & and_dcpl) ) begin
      IDX_LOOP_idx2_acc_1_psp_sva <= IDX_LOOP_idx2_acc_1_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx1_acc_psp_3_sva <= 9'b000000000;
    end
    else if ( ~(mux_466_nl & (~ (fsm_output[8]))) ) begin
      IDX_LOOP_idx1_acc_psp_3_sva <= IDX_LOOP_idx1_acc_psp_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm <= 1'b0;
    end
    else if ( ~(((or_44_cse | and_509_cse | (fsm_output[5])) ^ (fsm_output[6])) &
        and_dcpl) ) begin
      IDX_LOOP_3_slc_IDX_LOOP_acc_10_itm <= readslicef_11_1_10(IDX_LOOP_3_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_4_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_4_itm <= ~((IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_30_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_30_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_32_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_32_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_33_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_33_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_34_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_34_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_37_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_37_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_39_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_39_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_40_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_40_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_41_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_41_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_44_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_44_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_46_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_46_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_47_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_47_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_48_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_48_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_51_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_51_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_53_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_53_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_54_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_54_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_55_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_374 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_55_itm <= (IDX_LOOP_idx2_9_0_2_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx2_9_0_4_sva <= 10'b0000000000;
    end
    else if ( ~(mux_468_nl & (~ (fsm_output[8]))) ) begin
      IDX_LOOP_idx2_9_0_4_sva <= IDX_LOOP_idx2_9_0_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_slc_IDX_LOOP_acc_8_itm <= 1'b0;
    end
    else if ( ~(mux_469_nl & and_dcpl) ) begin
      IDX_LOOP_slc_IDX_LOOP_acc_8_itm <= readslicef_9_1_8(IDX_LOOP_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_8_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_8_itm <= ~((IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1:0]!=2'b00)
          | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_39_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_39_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1])) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_41_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_41_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[0])) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_42_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_42_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1:0]==2'b11) &
          (~ (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_43_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_43_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1:0]==2'b11) &
          (STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_47_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_47_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1])) & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_49_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_49_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[0])) & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_50_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_50_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1:0]==2'b11) &
          (~ (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_55_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_55_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1])) & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_58_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_58_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1:0]==2'b11) &
          (~ (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_59_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_59_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1:0]==2'b11) &
          (STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_63_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_63_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1])) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_66_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_66_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1:0]==2'b11) &
          (~ (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_67_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_377 ) begin
      IDX_LOOP_f1_and_67_itm <= (IDX_LOOP_idx2_acc_1_psp_sva_mx0w0[1:0]==2'b11) &
          (STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx2_acc_2_psp_sva <= 9'b000000000;
    end
    else if ( ~(mux_473_nl & (~ (fsm_output[8]))) ) begin
      IDX_LOOP_idx2_acc_2_psp_sva <= IDX_LOOP_idx2_acc_2_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx1_acc_2_psp_sva <= 8'b00000000;
    end
    else if ( ~ and_dcpl_367 ) begin
      IDX_LOOP_idx1_acc_2_psp_sva <= IDX_LOOP_idx1_acc_2_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm <= 1'b0;
    end
    else if ( (~(or_tmp_19 ^ (fsm_output[7]))) | (fsm_output[8]) ) begin
      IDX_LOOP_5_slc_IDX_LOOP_acc_10_itm <= readslicef_11_1_10(IDX_LOOP_5_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_12_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_12_itm <= ~((IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_88_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_88_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_89_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_89_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_93_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_93_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_95_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_95_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_96_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_96_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_97_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_97_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_100_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_100_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_102_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_102_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_103_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_103_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_104_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_104_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_107_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_107_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_109_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_109_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_110_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_110_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_111_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_380 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_111_itm <= (IDX_LOOP_idx2_9_0_4_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx2_9_0_6_sva <= 10'b0000000000;
    end
    else if ( ~(mux_476_nl & (~ (fsm_output[8]))) ) begin
      IDX_LOOP_idx2_9_0_6_sva <= IDX_LOOP_idx2_9_0_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm <= 1'b0;
    end
    else if ( ~(mux_478_nl & (~ (fsm_output[8]))) ) begin
      IDX_LOOP_6_slc_IDX_LOOP_acc_10_itm <= readslicef_11_1_10(IDX_LOOP_6_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_16_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_16_itm <= ~((IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1:0]!=2'b00)
          | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_75_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_75_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1])) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_77_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_77_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[0])) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_78_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_78_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1:0]==2'b11) &
          (~ (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_79_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_79_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1:0]==2'b11) &
          (STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_83_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_83_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1])) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_85_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_85_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[0])) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_86_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_86_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1:0]==2'b11) &
          (~ (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_87_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_87_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1:0]==2'b11) &
          (STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_91_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_91_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1])) & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_93_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_93_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[0])) & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_94_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_94_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1:0]==2'b11) &
          (~ (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_95_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_383 ) begin
      IDX_LOOP_f1_and_95_itm <= (IDX_LOOP_idx2_acc_2_psp_sva_mx0w0[1:0]==2'b11) &
          (STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx2_acc_3_psp_sva <= 9'b000000000;
    end
    else if ( ~(mux_480_nl & (~ (fsm_output[8]))) ) begin
      IDX_LOOP_idx2_acc_3_psp_sva <= IDX_LOOP_idx2_acc_3_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx1_acc_psp_7_sva <= 9'b000000000;
    end
    else if ( MUX_s_1_2_2((~ or_90_cse), or_tmp_26, fsm_output[8]) ) begin
      IDX_LOOP_idx1_acc_psp_7_sva <= IDX_LOOP_idx1_acc_psp_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm <= 1'b0;
    end
    else if ( ~(mux_483_nl & (~ (fsm_output[8]))) ) begin
      IDX_LOOP_7_slc_IDX_LOOP_acc_10_itm <= readslicef_11_1_10(IDX_LOOP_7_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_21_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_386 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_21_itm <= ~((IDX_LOOP_idx2_9_0_6_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_144_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_386 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_144_itm <= (IDX_LOOP_idx2_9_0_6_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_146_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_386 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_146_itm <= (IDX_LOOP_idx2_9_0_6_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_151_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_386 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_151_itm <= (IDX_LOOP_idx2_9_0_6_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_152_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_386 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_152_itm <= (IDX_LOOP_idx2_9_0_6_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_153_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_386 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_153_itm <= (IDX_LOOP_idx2_9_0_6_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_163_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_386 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_163_itm <= (IDX_LOOP_idx2_9_0_6_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_165_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_386 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_165_itm <= (IDX_LOOP_idx2_9_0_6_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_idx2_9_0_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2((~ or_90_cse), or_676_cse, fsm_output[8]) ) begin
      IDX_LOOP_idx2_9_0_sva <= IDX_LOOP_idx2_9_0_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_387 ) begin
      IDX_LOOP_slc_IDX_LOOP_acc_5_7_itm <= readslicef_8_1_7(IDX_LOOP_acc_5_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_24_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_388 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_24_itm <= ~((IDX_LOOP_idx2_acc_3_psp_sva_mx0w0[1:0]!=2'b00)
          | (STAGE_LOOP_op_rshift_psp_1_sva[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_121_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_388 ) begin
      IDX_LOOP_f1_and_121_itm <= (IDX_LOOP_idx2_acc_3_psp_sva_mx0w0[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_3_psp_sva_mx0w0[0])) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_123_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_388 ) begin
      IDX_LOOP_f1_and_123_itm <= (IDX_LOOP_idx2_acc_3_psp_sva_mx0w0[1:0]==2'b11)
          & (STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_131_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_388 ) begin
      IDX_LOOP_f1_and_131_itm <= (IDX_LOOP_idx2_acc_3_psp_sva_mx0w0[1:0]==2'b11)
          & (STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_1_slc_IDX_LOOP_acc_10_itm <= 1'b0;
    end
    else if ( ~(or_90_cse ^ (fsm_output[8])) ) begin
      IDX_LOOP_1_slc_IDX_LOOP_acc_10_itm <= z_out_2_10;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_28_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_nor_28_itm <= ~((IDX_LOOP_idx2_9_0_sva_mx0w0[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_208_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_208_itm <= (IDX_LOOP_idx2_9_0_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_209_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_209_itm <= (IDX_LOOP_idx2_9_0_sva_mx0w0[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_214_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_214_itm <= (IDX_LOOP_idx2_9_0_sva_mx0w0[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_219_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_219_itm <= (IDX_LOOP_idx2_9_0_sva_mx0w0[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_222_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_368 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_222_itm <= (IDX_LOOP_idx2_9_0_sva_mx0w0[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_101_itm <= 1'b0;
    end
    else if ( mux_490_nl | (fsm_output[8]) ) begin
      IDX_LOOP_f1_and_101_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_11_nl, IDX_LOOP_f1_and_101_nl,
          and_dcpl_159);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_102_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_390 ) begin
      IDX_LOOP_f1_and_102_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_13_nl, IDX_LOOP_f1_and_102_nl,
          and_dcpl_158);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_103_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_390 ) begin
      IDX_LOOP_f1_and_103_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_14_nl, IDX_LOOP_f1_and_103_nl,
          and_dcpl_158);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_111_itm <= 1'b0;
    end
    else if ( mux_492_nl | (fsm_output[8]) ) begin
      IDX_LOOP_f1_and_111_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_15_nl, IDX_LOOP_f1_and_111_nl,
          and_169_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_113_itm <= 1'b0;
      IDX_LOOP_f1_and_115_itm <= 1'b0;
      IDX_LOOP_f1_and_135_itm <= 1'b0;
      IDX_LOOP_f1_and_138_itm <= 1'b0;
      IDX_LOOP_f1_and_139_itm <= 1'b0;
    end
    else if ( IDX_LOOP_f1_or_69_cse ) begin
      IDX_LOOP_f1_and_113_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_19_nl, IDX_LOOP_f1_and_113_nl,
          and_dcpl_158);
      IDX_LOOP_f1_and_115_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_22_nl, IDX_LOOP_f1_and_115_nl,
          and_dcpl_158);
      IDX_LOOP_f1_and_135_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_31_nl, IDX_LOOP_f1_and_135_nl,
          and_dcpl_158);
      IDX_LOOP_f1_and_138_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_6_nl, IDX_LOOP_f1_and_138_nl,
          and_dcpl_158);
      IDX_LOOP_f1_and_139_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_7_nl, IDX_LOOP_f1_and_139_nl,
          and_dcpl_158);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_114_itm <= 1'b0;
      IDX_LOOP_f1_and_119_itm <= 1'b0;
      IDX_LOOP_f1_and_127_itm <= 1'b0;
    end
    else if ( IDX_LOOP_f1_or_70_cse ) begin
      IDX_LOOP_f1_and_114_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_21_nl, IDX_LOOP_f1_and_114_nl,
          and_dcpl_109);
      IDX_LOOP_f1_and_119_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_23_nl, IDX_LOOP_f1_and_119_nl,
          and_dcpl_109);
      IDX_LOOP_f1_and_127_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_29_nl, IDX_LOOP_f1_and_127_nl,
          and_dcpl_109);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_122_itm <= 1'b0;
    end
    else if ( mux_495_nl | (fsm_output[8]) ) begin
      IDX_LOOP_f1_and_122_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_27_nl, IDX_LOOP_f1_and_122_nl,
          and_164_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_129_itm <= 1'b0;
    end
    else if ( ~(mux_496_nl & (~ (fsm_output[8]))) ) begin
      IDX_LOOP_f1_and_129_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_3_nl, IDX_LOOP_f1_and_129_nl,
          and_166_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_130_itm <= 1'b0;
    end
    else if ( mux_497_nl | (fsm_output[8]) ) begin
      IDX_LOOP_f1_and_130_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_30_nl, IDX_LOOP_f1_and_130_nl,
          and_dcpl_159);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_137_itm <= 1'b0;
    end
    else if ( mux_499_nl | (fsm_output[8]) ) begin
      IDX_LOOP_f1_and_137_itm <= MUX_s_1_2_2(IDX_LOOP_f1_and_5_nl, IDX_LOOP_f1_and_137_nl,
          and_412_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_IDX_LOOP_and_104_itm <= 1'b0;
    end
    else if ( mux_501_nl | (fsm_output[8]) ) begin
      IDX_LOOP_IDX_LOOP_and_104_itm <= MUX_s_1_2_2(IDX_LOOP_IDX_LOOP_and_2_nl, IDX_LOOP_f2_IDX_LOOP_f2_and_215_nl,
          and_416_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_51_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_404 ) begin
      IDX_LOOP_f1_and_51_itm <= MUX_s_1_2_2(IDX_LOOP_f2_IDX_LOOP_f2_nor_cse, IDX_LOOP_f1_and_51_nl,
          and_dcpl_109);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_57_itm <= 1'b0;
    end
    else if ( ~(((or_51_cse | (fsm_output[2]) | (fsm_output[5])) ^ (fsm_output[6]))
        & and_dcpl) ) begin
      IDX_LOOP_f1_and_57_itm <= (IDX_LOOP_idx2_acc_1_psp_sva[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_1_psp_sva[0])) & IDX_LOOP_f1_equal_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_90_itm <= 1'b0;
    end
    else if ( ~(mux_504_nl & and_dcpl) ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_90_itm <= (IDX_LOOP_idx2_9_0_4_sva[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_99_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_390 ) begin
      IDX_LOOP_f1_and_99_itm <= (IDX_LOOP_idx2_acc_2_psp_sva[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_2_psp_sva[1])) & IDX_LOOP_f1_equal_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_142_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_142_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_149_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_149_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_156_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_156_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_159_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_159_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_160_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_160_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_166_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_166_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_200_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_408 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_200_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_223_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_408 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_223_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_mux1h_5_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_509_nl | (fsm_output[8]) ) begin
      IDX_LOOP_mux1h_5_itm <= IDX_LOOP_mux1h_68_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_modulo_dev_return_1_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_dcpl_158 | IDX_LOOP_modulo_dev_return_1_sva_mx0c1 | and_dcpl_413
        | and_dcpl_114 | and_dcpl_207 | and_dcpl_117 | and_dcpl_120 | and_dcpl_219
        | and_dcpl_123 | and_dcpl_125 | and_dcpl_227 | and_dcpl_127 | and_dcpl_129
        ) begin
      IDX_LOOP_modulo_dev_return_1_sva <= MUX1HOT_v_64_11_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
          vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
          vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, IDX_LOOP_1_modulo_dev_cmp_return_rsc_z,
          z_out_7, z_out_8, {IDX_LOOP_f2_and_nl , IDX_LOOP_f2_and_1_nl , IDX_LOOP_f2_or_nl
          , IDX_LOOP_f2_and_3_nl , IDX_LOOP_f2_or_1_nl , IDX_LOOP_f2_or_4_nl , IDX_LOOP_f2_and_6_nl
          , IDX_LOOP_f2_and_7_nl , IDX_LOOP_modulo_dev_return_1_sva_mx0c1 , IDX_LOOP_f2_or_2_nl
          , IDX_LOOP_f2_or_3_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_mux1h_1_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(mux_513_nl & and_dcpl_15) ) begin
      IDX_LOOP_mux1h_1_itm <= IDX_LOOP_mux1h_68_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f1_and_65_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_404 ) begin
      IDX_LOOP_f1_and_65_itm <= (IDX_LOOP_idx2_acc_1_psp_sva[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
          & (~ (IDX_LOOP_idx2_acc_1_psp_sva[0])) & IDX_LOOP_f1_equal_tmp_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_86_itm <= 1'b0;
    end
    else if ( ~((~ mux_514_nl) & and_dcpl) ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_86_itm <= (IDX_LOOP_idx2_9_0_4_sva[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_145_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_416 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_145_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_158_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_416 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_158_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_212_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_417 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_212_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_221_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_417 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_221_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_10_lpi_4_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_dcpl_109 | and_dcpl_247 | and_dcpl_207 | and_dcpl_254 | and_dcpl_219
        | and_dcpl_261 | and_dcpl_227 | and_dcpl_267 ) begin
      tmp_10_lpi_4_dfm <= MUX1HOT_v_64_5_2(z_out_4, vec_rsc_0_1_i_q_d, vec_rsc_0_3_i_q_d,
          vec_rsc_0_5_i_q_d, vec_rsc_0_7_i_q_d, {(~ IDX_LOOP_f1_or_64_tmp) , IDX_LOOP_f1_and_208_nl
          , IDX_LOOP_f1_and_209_nl , IDX_LOOP_f1_and_210_nl , IDX_LOOP_f1_and_211_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_mux1h_2_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~((~ mux_519_nl) & and_dcpl) ) begin
      IDX_LOOP_mux1h_2_itm <= IDX_LOOP_mux1h_68_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_201_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_419 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_201_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b110)
          & IDX_LOOP_f1_equal_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_202_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_419 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_202_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_216_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_419 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_216_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_mux1h_3_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~((~ mux_521_nl) & and_dcpl) ) begin
      IDX_LOOP_mux1h_3_itm <= IDX_LOOP_mux1h_68_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_167_itm <= 1'b0;
    end
    else if ( mux_522_nl | (fsm_output[8]) ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_167_itm <= (IDX_LOOP_idx2_9_0_6_sva[2:0]==3'b111)
          & IDX_LOOP_f1_equal_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_mux1h_4_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( (~(or_tmp_516 ^ (fsm_output[7]))) | (fsm_output[8]) ) begin
      IDX_LOOP_mux1h_4_itm <= IDX_LOOP_mux1h_68_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_1_mul_mut <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( (and_dcpl_135 & xnor_cse & and_dcpl_95 & (~ (fsm_output[6])) & (~ (fsm_output[8])))
        | (and_dcpl_138 & and_dcpl_113) | (and_dcpl_138 & and_dcpl_116) | (and_dcpl_138
        & and_dcpl_119) | (and_dcpl_138 & and_dcpl_122) | (and_dcpl_138 & and_dcpl_126)
        | (and_dcpl_138 & and_dcpl_128) ) begin
      IDX_LOOP_1_mul_mut <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_205_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_423 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_205_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_207_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_423 ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_207_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b101)
          & IDX_LOOP_f1_equal_tmp_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_mux1h_6_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_526_nl | (fsm_output[8]) ) begin
      IDX_LOOP_mux1h_6_itm <= IDX_LOOP_mux1h_68_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_198_itm <= 1'b0;
    end
    else if ( mux_527_nl | (fsm_output[8]) ) begin
      IDX_LOOP_f2_IDX_LOOP_f2_and_198_itm <= (IDX_LOOP_idx2_9_0_sva[2:0]==3'b011)
          & IDX_LOOP_f1_equal_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      IDX_LOOP_mux1h_7_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_529_nl | (fsm_output[8]) ) begin
      IDX_LOOP_mux1h_7_itm <= IDX_LOOP_mux1h_68_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7 <= 2'b00;
    end
    else if ( ~ and_dcpl_367 ) begin
      reg_IDX_LOOP_1_idx1_mul_sdt_ftd_7 <= z_out_5[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_IDX_LOOP_t_10_3_ftd_1 <= 7'b0000000;
    end
    else if ( ~ and_dcpl_387 ) begin
      reg_IDX_LOOP_t_10_3_ftd_1 <= z_out_1[6:0];
    end
  end
  assign nor_230_nl = ~((fsm_output[7:5]!=3'b000) | or_tmp_16);
  assign mux_187_nl = MUX_s_1_2_2(or_676_cse, nor_230_nl, fsm_output[8]);
  assign or_202_nl = (fsm_output[7:5]!=3'b000);
  assign mux_190_nl = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), or_202_nl);
  assign or_203_nl = (fsm_output[3]) | mux_190_nl;
  assign or_201_nl = (~ (fsm_output[3])) | (fsm_output[8]);
  assign mux_191_nl = MUX_s_1_2_2(or_203_nl, or_201_nl, or_200_cse);
  assign mux_192_nl = MUX_s_1_2_2(mux_191_nl, (fsm_output[8]), fsm_output[4]);
  assign IDX_LOOP_f2_or_5_nl = IDX_LOOP_f2_and_8_cse | IDX_LOOP_f2_and_10_cse | IDX_LOOP_f2_and_14_cse;
  assign IDX_LOOP_f2_or_6_nl = IDX_LOOP_f2_and_9_cse | IDX_LOOP_f2_and_11_cse | IDX_LOOP_f2_and_15_cse;
  assign GROUP_LOOP_j_not_1_nl = ~ GROUP_LOOP_j_10_0_sva_9_0_mx0c0;
  assign or_690_nl = (~ (fsm_output[0])) | (fsm_output[2]);
  assign or_691_nl = (fsm_output[0]) | (~ (fsm_output[2]));
  assign mux_182_nl = MUX_s_1_2_2(or_690_nl, or_691_nl, fsm_output[8]);
  assign or_nl = mux_182_nl | (~ and_dcpl_96) | (fsm_output[1]) | (fsm_output[6])
      | (fsm_output[5]) | (fsm_output[7]);
  assign or_697_nl = (~((fsm_output[1]) | (fsm_output[8]))) | (fsm_output[7:5]!=3'b000);
  assign mux_531_nl = MUX_s_1_2_2(or_697_nl, or_tmp_545, fsm_output[2]);
  assign mux_530_nl = MUX_s_1_2_2(or_tmp_545, or_tmp, or_200_cse);
  assign mux_532_nl = MUX_s_1_2_2(mux_531_nl, mux_530_nl, fsm_output[3]);
  assign mux_29_nl = MUX_s_1_2_2((~ or_tmp_3), or_tmp_4, fsm_output[6]);
  assign mux_459_nl = MUX_s_1_2_2(mux_29_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_27_nl = MUX_s_1_2_2((~ or_tmp_3), or_tmp_2, fsm_output[6]);
  assign mux_461_nl = MUX_s_1_2_2(mux_27_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_465_nl = MUX_s_1_2_2(or_47_cse, (~ and_tmp_9), fsm_output[5]);
  assign nor_300_nl = ~((fsm_output[6:1]!=6'b000000));
  assign mux_466_nl = MUX_s_1_2_2(or_tmp_19, nor_300_nl, fsm_output[7]);
  assign nl_IDX_LOOP_3_acc_nl = ({1'b1 , (~ STAGE_LOOP_op_rshift_psp_1_sva)}) + conv_u2s_10_11({IDX_LOOP_t_10_3_sva_6_0
      , 3'b010}) + 11'b00000000001;
  assign IDX_LOOP_3_acc_nl = nl_IDX_LOOP_3_acc_nl[10:0];
  assign nor_251_nl = ~((fsm_output[6:0]!=7'b0000000));
  assign mux_468_nl = MUX_s_1_2_2(or_tmp_19, nor_251_nl, fsm_output[7]);
  assign nl_IDX_LOOP_acc_nl = ({1'b1 , (~ (STAGE_LOOP_op_rshift_psp_1_sva[9:2]))})
      + conv_u2u_8_9({IDX_LOOP_t_10_3_sva_6_0 , 1'b0}) + 9'b000000001;
  assign IDX_LOOP_acc_nl = nl_IDX_LOOP_acc_nl[8:0];
  assign mux_469_nl = MUX_s_1_2_2(or_47_cse, (~ and_tmp_10), fsm_output[5]);
  assign or_35_nl = (fsm_output[6]) | (fsm_output[1]) | (fsm_output[0]) | (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[4]);
  assign mux_472_nl = MUX_s_1_2_2((fsm_output[6]), or_35_nl, fsm_output[5]);
  assign mux_473_nl = MUX_s_1_2_2(or_tmp_19, (~ mux_472_nl), fsm_output[7]);
  assign nl_IDX_LOOP_5_acc_nl = ({1'b1 , (~ STAGE_LOOP_op_rshift_psp_1_sva)}) + conv_u2s_10_11({IDX_LOOP_t_10_3_sva_6_0
      , 3'b100}) + 11'b00000000001;
  assign IDX_LOOP_5_acc_nl = nl_IDX_LOOP_5_acc_nl[10:0];
  assign mux_475_nl = MUX_s_1_2_2(and_tmp_9, (fsm_output[6]), fsm_output[5]);
  assign mux_476_nl = MUX_s_1_2_2(or_tmp_19, (~ mux_475_nl), fsm_output[7]);
  assign nl_IDX_LOOP_6_acc_nl = ({1'b1 , (~ STAGE_LOOP_op_rshift_psp_1_sva)}) + conv_u2s_10_11({IDX_LOOP_t_10_3_sva_6_0
      , 3'b101}) + 11'b00000000001;
  assign IDX_LOOP_6_acc_nl = nl_IDX_LOOP_6_acc_nl[10:0];
  assign mux_477_nl = MUX_s_1_2_2((fsm_output[6]), or_47_cse, fsm_output[5]);
  assign mux_478_nl = MUX_s_1_2_2(or_tmp_19, (~ mux_477_nl), fsm_output[7]);
  assign nand_15_nl = ~((fsm_output[6:5]==2'b11) & or_tmp_2);
  assign mux_480_nl = MUX_s_1_2_2(or_tmp_19, nand_15_nl, fsm_output[7]);
  assign nl_IDX_LOOP_7_acc_nl = ({1'b1 , (~ STAGE_LOOP_op_rshift_psp_1_sva)}) + conv_u2s_10_11({IDX_LOOP_t_10_3_sva_6_0
      , 3'b110}) + 11'b00000000001;
  assign IDX_LOOP_7_acc_nl = nl_IDX_LOOP_7_acc_nl[10:0];
  assign mux_482_nl = MUX_s_1_2_2(and_tmp_10, (fsm_output[6]), fsm_output[5]);
  assign mux_483_nl = MUX_s_1_2_2(or_tmp_19, (~ mux_482_nl), fsm_output[7]);
  assign nl_IDX_LOOP_acc_5_nl = ({1'b1 , (~ (STAGE_LOOP_op_rshift_psp_1_sva[9:3]))})
      + conv_u2u_7_8(IDX_LOOP_t_10_3_sva_6_0) + 8'b00000001;
  assign IDX_LOOP_acc_5_nl = nl_IDX_LOOP_acc_5_nl[7:0];
  assign IDX_LOOP_f1_and_11_nl = (IDX_LOOP_idx2_acc_tmp[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_tmp[1])) & IDX_LOOP_f1_equal_tmp_1_mx0w0;
  assign IDX_LOOP_f1_and_101_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_2_psp_sva[0])) & IDX_LOOP_f1_equal_tmp_1;
  assign mux_490_nl = MUX_s_1_2_2(not_tmp_290, or_tmp_502, fsm_output[7]);
  assign IDX_LOOP_f1_and_13_nl = (IDX_LOOP_idx2_acc_tmp[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_tmp[0])) & IDX_LOOP_f1_equal_tmp_1_mx0w0;
  assign IDX_LOOP_f1_and_102_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]==2'b11) & (~
      (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f1_and_14_nl = (IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]))
      & IDX_LOOP_f1_equal_tmp_1_mx0w0;
  assign IDX_LOOP_f1_and_103_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f1_and_15_nl = (IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & IDX_LOOP_f1_equal_tmp_1_mx0w0;
  assign IDX_LOOP_f1_and_111_nl = (IDX_LOOP_idx2_acc_3_psp_sva[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_3_psp_sva[1])) & IDX_LOOP_f1_equal_tmp_1;
  assign and_169_nl = and_dcpl_135 & and_dcpl_102 & and_dcpl_94;
  assign mux_492_nl = MUX_s_1_2_2(not_tmp_292, mux_tmp_461, fsm_output[7]);
  assign IDX_LOOP_f1_and_19_nl = (IDX_LOOP_idx2_acc_tmp[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_tmp[1])) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
  assign IDX_LOOP_f1_and_113_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_3_psp_sva[0])) & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f1_and_22_nl = (IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]))
      & IDX_LOOP_f1_equal_tmp_2_mx0w0;
  assign IDX_LOOP_f1_and_115_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f1_and_31_nl = (IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & IDX_LOOP_f1_equal_tmp_3_mx0w0;
  assign IDX_LOOP_f1_and_135_nl = (IDX_LOOP_idx2_acc_3_psp_sva[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_3_psp_sva[1])) & IDX_LOOP_f1_equal_tmp;
  assign IDX_LOOP_f1_and_6_nl = (IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]))
      & IDX_LOOP_f1_equal_tmp_mx0w0;
  assign IDX_LOOP_f1_and_138_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11) & (~
      (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp;
  assign IDX_LOOP_f1_and_7_nl = (IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & IDX_LOOP_f1_equal_tmp_mx0w0;
  assign IDX_LOOP_f1_and_139_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & IDX_LOOP_f1_equal_tmp;
  assign IDX_LOOP_f1_and_21_nl = (IDX_LOOP_idx2_acc_tmp[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_tmp[0])) & IDX_LOOP_f1_equal_tmp_2_mx0w0;
  assign IDX_LOOP_f1_and_114_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11) & (~
      (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f1_and_23_nl = (IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & IDX_LOOP_f1_equal_tmp_2_mx0w0;
  assign IDX_LOOP_f1_and_119_nl = (IDX_LOOP_idx2_acc_3_psp_sva[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_3_psp_sva[1])) & IDX_LOOP_f1_equal_tmp_2;
  assign IDX_LOOP_f1_and_29_nl = (IDX_LOOP_idx2_acc_tmp[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_tmp[0])) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
  assign IDX_LOOP_f1_and_127_nl = (IDX_LOOP_idx2_acc_3_psp_sva[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_3_psp_sva[1])) & IDX_LOOP_f1_equal_tmp_3;
  assign IDX_LOOP_f1_and_27_nl = (IDX_LOOP_idx2_acc_tmp[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_tmp[1])) & IDX_LOOP_f1_equal_tmp_3_mx0w0;
  assign IDX_LOOP_f1_and_122_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11) & (~
      (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_2;
  assign and_164_nl = and_dcpl_103 & and_dcpl_153 & and_dcpl_94;
  assign mux_495_nl = MUX_s_1_2_2(not_tmp_298, mux_tmp_461, fsm_output[7]);
  assign IDX_LOOP_f1_and_3_nl = (IDX_LOOP_idx2_acc_tmp[0]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_tmp[1])) & IDX_LOOP_f1_equal_tmp_mx0w0;
  assign IDX_LOOP_f1_and_129_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_3_psp_sva[0])) & IDX_LOOP_f1_equal_tmp_3;
  assign and_166_nl = and_dcpl_103 & and_509_cse & and_dcpl_94;
  assign mux_496_nl = MUX_s_1_2_2(or_tmp_516, (~ mux_tmp_461), fsm_output[7]);
  assign IDX_LOOP_f1_and_30_nl = (IDX_LOOP_idx2_acc_tmp[1:0]==2'b11) & (~ (STAGE_LOOP_op_rshift_psp_1_sva[0]))
      & IDX_LOOP_f1_equal_tmp_3_mx0w0;
  assign IDX_LOOP_f1_and_130_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1:0]==2'b11) & (~
      (STAGE_LOOP_op_rshift_psp_1_sva[0])) & IDX_LOOP_f1_equal_tmp_3;
  assign mux_497_nl = MUX_s_1_2_2(not_tmp_290, mux_tmp_461, fsm_output[7]);
  assign IDX_LOOP_f1_and_5_nl = (IDX_LOOP_idx2_acc_tmp[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_tmp[0])) & IDX_LOOP_f1_equal_tmp_mx0w0;
  assign IDX_LOOP_f1_and_137_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1]) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & (~ (IDX_LOOP_idx2_acc_3_psp_sva[0])) & IDX_LOOP_f1_equal_tmp;
  assign and_412_nl = and_dcpl_135 & and_509_cse & and_dcpl_94;
  assign mux_498_nl = MUX_s_1_2_2((fsm_output[4]), or_51_cse, fsm_output[2]);
  assign nor_117_nl = ~((fsm_output[6:5]!=2'b00) | mux_498_nl);
  assign mux_499_nl = MUX_s_1_2_2(nor_117_nl, mux_tmp_461, fsm_output[7]);
  assign IDX_LOOP_IDX_LOOP_and_2_nl = (z_out_6[2:0]==3'b011);
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_215_nl = (IDX_LOOP_idx2_9_0_sva[2:0]==3'b110)
      & IDX_LOOP_f1_equal_tmp_3;
  assign and_416_nl = and_dcpl_134 & (fsm_output[2]) & and_dcpl_95 & and_dcpl_94;
  assign mux_500_nl = MUX_s_1_2_2((fsm_output[4]), or_51_cse, and_448_cse);
  assign nor_116_nl = ~((fsm_output[6:5]!=2'b00) | mux_500_nl);
  assign mux_501_nl = MUX_s_1_2_2(nor_116_nl, and_tmp_7, fsm_output[7]);
  assign IDX_LOOP_f1_and_51_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1:0]==2'b11) & (STAGE_LOOP_op_rshift_psp_1_sva[0])
      & IDX_LOOP_f1_equal_tmp;
  assign mux_504_nl = MUX_s_1_2_2(or_tmp_505, (~ and_tmp_11), fsm_output[5]);
  assign or_633_nl = (fsm_output[2]) | (fsm_output[4]);
  assign mux_508_nl = MUX_s_1_2_2(or_633_nl, or_44_cse, or_680_cse);
  assign nor_115_nl = ~((fsm_output[6:5]!=2'b00) | mux_508_nl);
  assign or_630_nl = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[3]);
  assign mux_507_nl = MUX_s_1_2_2((fsm_output[6]), or_630_nl, fsm_output[5]);
  assign mux_509_nl = MUX_s_1_2_2(nor_115_nl, mux_507_nl, fsm_output[7]);
  assign IDX_LOOP_f2_and_nl = ((IDX_LOOP_f1_and_51_itm & IDX_LOOP_f1_equal_tmp) |
      (IDX_LOOP_f1_and_51_itm & IDX_LOOP_f1_equal_tmp_1) | (IDX_LOOP_f1_and_51_itm
      & IDX_LOOP_f1_equal_tmp_2) | (IDX_LOOP_f1_and_51_itm & IDX_LOOP_f1_equal_tmp_3))
      & and_dcpl_158;
  assign IDX_LOOP_f2_and_1_nl = (((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_cse_1
      & IDX_LOOP_f1_equal_tmp_3)) & and_dcpl_158;
  assign IDX_LOOP_f2_or_nl = ((((IDX_LOOP_idx2_acc_psp_sva[0]) & IDX_LOOP_f2_nor_1_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_acc_psp_sva[0]) & IDX_LOOP_f2_nor_1_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_acc_psp_sva[0]) & IDX_LOOP_f2_nor_1_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_acc_psp_sva[0]) & IDX_LOOP_f2_nor_1_cse_1
      & IDX_LOOP_f1_equal_tmp_3)) & and_dcpl_158) | IDX_LOOP_f2_and_8_cse | IDX_LOOP_f2_and_10_cse
      | IDX_LOOP_f2_and_14_cse;
  assign IDX_LOOP_f2_and_3_nl = (IDX_LOOP_f1_and_129_itm | IDX_LOOP_f1_and_101_itm
      | IDX_LOOP_f1_and_113_itm | IDX_LOOP_f1_and_122_itm) & and_dcpl_158;
  assign IDX_LOOP_f2_or_1_nl = ((((IDX_LOOP_idx2_acc_psp_sva[1]) & IDX_LOOP_f2_nor_2_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_acc_psp_sva[1]) & IDX_LOOP_f2_nor_2_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_acc_psp_sva[1]) & IDX_LOOP_f2_nor_2_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_acc_psp_sva[1]) & IDX_LOOP_f2_nor_2_cse_1
      & IDX_LOOP_f1_equal_tmp_3)) & and_dcpl_158) | IDX_LOOP_f2_and_9_cse | IDX_LOOP_f2_and_11_cse
      | IDX_LOOP_f2_and_15_cse;
  assign IDX_LOOP_f2_or_4_nl = ((IDX_LOOP_f1_and_137_itm | IDX_LOOP_f1_and_102_itm
      | IDX_LOOP_f1_and_114_itm | IDX_LOOP_f1_and_127_itm) & and_dcpl_158) | and_dcpl_413;
  assign IDX_LOOP_f2_and_6_nl = (IDX_LOOP_f1_and_138_itm | IDX_LOOP_f1_and_103_itm
      | IDX_LOOP_f1_and_115_itm | IDX_LOOP_f1_and_130_itm) & and_dcpl_158;
  assign IDX_LOOP_f2_and_7_nl = (IDX_LOOP_f1_and_139_itm | IDX_LOOP_f1_and_111_itm
      | IDX_LOOP_f1_and_119_itm | IDX_LOOP_f1_and_135_itm) & and_dcpl_158;
  assign IDX_LOOP_f2_or_2_nl = and_dcpl_114 | and_dcpl_120 | and_dcpl_125 | and_dcpl_129;
  assign IDX_LOOP_f2_or_3_nl = and_dcpl_117 | and_dcpl_123 | and_dcpl_127;
  assign mux_513_nl = MUX_s_1_2_2(or_tmp_11, (~ or_51_cse), fsm_output[5]);
  assign nor_114_nl = ~((fsm_output[6]) | or_tmp_11);
  assign mux_514_nl = MUX_s_1_2_2(nor_114_nl, and_tmp_11, fsm_output[5]);
  assign IDX_LOOP_f1_mux1h_201_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_equal_tmp, IDX_LOOP_f1_equal_tmp_3,
      IDX_LOOP_f1_equal_tmp_2, IDX_LOOP_f1_equal_tmp_1, {and_dcpl_476 , and_dcpl_479
      , and_dcpl_482 , and_dcpl_484});
  assign IDX_LOOP_f1_and_208_nl = IDX_LOOP_f1_mux1h_201_nl & IDX_LOOP_f1_or_64_tmp;
  assign IDX_LOOP_f1_mux1h_202_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_equal_tmp_1, IDX_LOOP_f1_equal_tmp,
      IDX_LOOP_f1_equal_tmp_3, IDX_LOOP_f1_equal_tmp_2, {and_dcpl_476 , and_dcpl_479
      , and_dcpl_482 , and_dcpl_484});
  assign IDX_LOOP_f1_and_209_nl = IDX_LOOP_f1_mux1h_202_nl & IDX_LOOP_f1_or_64_tmp;
  assign IDX_LOOP_f1_mux1h_203_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_equal_tmp_2, IDX_LOOP_f1_equal_tmp_1,
      IDX_LOOP_f1_equal_tmp, IDX_LOOP_f1_equal_tmp_3, {and_dcpl_476 , and_dcpl_479
      , and_dcpl_482 , and_dcpl_484});
  assign IDX_LOOP_f1_and_210_nl = IDX_LOOP_f1_mux1h_203_nl & IDX_LOOP_f1_or_64_tmp;
  assign IDX_LOOP_f1_mux1h_204_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_equal_tmp_3, IDX_LOOP_f1_equal_tmp_2,
      IDX_LOOP_f1_equal_tmp_1, IDX_LOOP_f1_equal_tmp, {and_dcpl_476 , and_dcpl_479
      , and_dcpl_482 , and_dcpl_484});
  assign IDX_LOOP_f1_and_211_nl = IDX_LOOP_f1_mux1h_204_nl & IDX_LOOP_f1_or_64_tmp;
  assign mux_518_nl = MUX_s_1_2_2((~ or_tmp_16), or_51_cse, fsm_output[6]);
  assign mux_519_nl = MUX_s_1_2_2(mux_518_nl, (fsm_output[6]), fsm_output[5]);
  assign nor_113_nl = ~((fsm_output[6]) | or_40_cse);
  assign mux_521_nl = MUX_s_1_2_2(nor_113_nl, and_tmp_14, fsm_output[5]);
  assign mux_522_nl = MUX_s_1_2_2(not_tmp_298, mux_tmp_457, fsm_output[7]);
  assign mux_525_nl = MUX_s_1_2_2(and_tmp_14, (fsm_output[6]), fsm_output[5]);
  assign mux_526_nl = MUX_s_1_2_2(not_tmp_292, mux_525_nl, fsm_output[7]);
  assign mux_527_nl = MUX_s_1_2_2(not_tmp_292, and_tmp_7, fsm_output[7]);
  assign or_657_nl = and_509_cse | (fsm_output[2]);
  assign mux_528_nl = MUX_s_1_2_2((fsm_output[4]), or_51_cse, or_657_nl);
  assign nor_260_nl = ~((fsm_output[6:5]!=2'b00) | mux_528_nl);
  assign and_521_nl = (fsm_output[6:5]==2'b11) & or_51_cse;
  assign mux_529_nl = MUX_s_1_2_2(nor_260_nl, and_521_nl, fsm_output[7]);
  assign IDX_LOOP_mux_25_nl = MUX_v_10_2_2((~ STAGE_LOOP_op_rshift_psp_1_sva), GROUP_LOOP_j_10_0_sva_9_0,
      and_dcpl_443);
  assign IDX_LOOP_IDX_LOOP_nand_1_nl = ~(and_dcpl_443 & (~(and_dcpl_436 & (fsm_output[2:1]==2'b01)
      & nor_327_cse & and_dcpl_431)));
  assign not_1293_nl = ~ and_dcpl_443;
  assign IDX_LOOP_IDX_LOOP_and_132_nl = MUX_v_7_2_2(7'b0000000, IDX_LOOP_t_10_3_sva_6_0,
      not_1293_nl);
  assign nl_acc_nl = ({(~ and_dcpl_443) , IDX_LOOP_mux_25_nl , IDX_LOOP_IDX_LOOP_nand_1_nl})
      + conv_u2u_11_12({IDX_LOOP_IDX_LOOP_and_132_nl , 4'b0011});
  assign acc_nl = nl_acc_nl[11:0];
  assign z_out = readslicef_12_11_1(acc_nl);
  assign STAGE_LOOP_gp_mux_5_nl = MUX_v_7_2_2(({3'b000 , STAGE_LOOP_i_3_0_sva}),
      IDX_LOOP_t_10_3_sva_6_0, and_dcpl_454);
  assign nl_z_out_1 = conv_u2u_7_8(STAGE_LOOP_gp_mux_5_nl) + conv_s2u_2_8({(~ and_dcpl_454)
      , 1'b1});
  assign z_out_1 = nl_z_out_1[7:0];
  assign IDX_LOOP_mux_26_nl = MUX_v_11_2_2(({z_out_1 , 3'b000}), z_out, and_dcpl_468);
  assign IDX_LOOP_mux_27_nl = MUX_v_10_2_2((~ STAGE_LOOP_op_rshift_psp_1_sva), (~
      STAGE_LOOP_gp_lshift_psp_sva), and_dcpl_468);
  assign nl_acc_2_nl = ({IDX_LOOP_mux_26_nl , 1'b1}) + ({1'b1 , IDX_LOOP_mux_27_nl
      , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[11:0];
  assign z_out_2_10 = readslicef_12_1_11(acc_2_nl);
  assign and_719_nl = and_dcpl_509 & nor_327_cse & xnor_cse;
  assign and_720_nl = and_dcpl_509 & nor_327_cse & and_dcpl_469;
  assign and_721_nl = and_dcpl_509 & and_dcpl_477 & and_dcpl_431;
  assign and_722_nl = and_dcpl_509 & and_dcpl_477 & and_dcpl_469;
  assign and_723_nl = and_dcpl_509 & nor_327_cse & and_dcpl_493;
  assign and_724_nl = and_dcpl_509 & and_dcpl_477 & and_dcpl_493;
  assign and_725_nl = and_dcpl_509 & and_dcpl_477 & (fsm_output[5]) & (fsm_output[7]);
  assign IDX_LOOP_mux1h_102_nl = MUX1HOT_v_64_8_2(IDX_LOOP_mux1h_5_itm, IDX_LOOP_mux1h_1_itm,
      IDX_LOOP_mux1h_2_itm, IDX_LOOP_mux1h_3_itm, IDX_LOOP_mux1h_4_itm, IDX_LOOP_mux1h_6_itm,
      IDX_LOOP_mux1h_7_itm, ({55'b0000000000000000000000000000000000000000000000000000000
      , (GROUP_LOOP_j_10_0_sva_9_0[8:0])}), {and_719_nl , and_720_nl , and_721_nl
      , and_722_nl , and_723_nl , and_724_nl , and_725_nl , and_dcpl_533});
  assign IDX_LOOP_mux_28_nl = MUX_v_64_2_2(IDX_LOOP_1_modulo_dev_cmp_return_rsc_z,
      ({55'b0000000000000000000000000000000000000000000000000000000 , (STAGE_LOOP_op_rshift_psp_1_sva[8:0])}),
      and_dcpl_533);
  assign z_out_5 = conv_u2u_128_128(IDX_LOOP_mux1h_102_nl * IDX_LOOP_mux_28_nl);
  assign IDX_LOOP_f1_mux1h_205_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_equal_tmp_3, IDX_LOOP_f1_equal_tmp_2,
      IDX_LOOP_f1_equal_tmp_1, IDX_LOOP_f1_equal_tmp, {and_dcpl_492 , and_dcpl_496
      , and_dcpl_498 , and_dcpl_503});
  assign IDX_LOOP_f1_mux1h_206_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_equal_tmp, IDX_LOOP_f1_equal_tmp_3,
      IDX_LOOP_f1_equal_tmp_2, IDX_LOOP_f1_equal_tmp_1, {and_dcpl_492 , and_dcpl_496
      , and_dcpl_498 , and_dcpl_503});
  assign IDX_LOOP_f1_mux1h_207_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_equal_tmp_1, IDX_LOOP_f1_equal_tmp,
      IDX_LOOP_f1_equal_tmp_3, IDX_LOOP_f1_equal_tmp_2, {and_dcpl_492 , and_dcpl_496
      , and_dcpl_498 , and_dcpl_503});
  assign IDX_LOOP_f1_mux1h_208_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_equal_tmp_2, IDX_LOOP_f1_equal_tmp_1,
      IDX_LOOP_f1_equal_tmp, IDX_LOOP_f1_equal_tmp_3, {and_dcpl_492 , and_dcpl_496
      , and_dcpl_498 , and_dcpl_503});
  assign z_out_4 = MUX1HOT_v_64_4_2(vec_rsc_0_0_i_q_d, vec_rsc_0_2_i_q_d, vec_rsc_0_4_i_q_d,
      vec_rsc_0_6_i_q_d, {IDX_LOOP_f1_mux1h_205_nl , IDX_LOOP_f1_mux1h_206_nl , IDX_LOOP_f1_mux1h_207_nl
      , IDX_LOOP_f1_mux1h_208_nl});
  assign IDX_LOOP_f1_or_82_nl = (IDX_LOOP_f2_IDX_LOOP_f2_nor_4_itm & IDX_LOOP_f1_equal_tmp)
      | (IDX_LOOP_f2_IDX_LOOP_f2_nor_4_itm & IDX_LOOP_f1_equal_tmp_1) | (IDX_LOOP_f2_IDX_LOOP_f2_nor_4_itm
      & IDX_LOOP_f1_equal_tmp_2) | (IDX_LOOP_f2_IDX_LOOP_f2_nor_4_itm & IDX_LOOP_f1_equal_tmp_3);
  assign IDX_LOOP_f1_or_83_nl = (IDX_LOOP_f2_IDX_LOOP_f2_nor_12_itm & IDX_LOOP_f1_equal_tmp_3)
      | (IDX_LOOP_f2_IDX_LOOP_f2_nor_12_itm & IDX_LOOP_f1_equal_tmp) | (IDX_LOOP_f2_IDX_LOOP_f2_nor_12_itm
      & IDX_LOOP_f1_equal_tmp_1) | (IDX_LOOP_f2_IDX_LOOP_f2_nor_12_itm & IDX_LOOP_f1_equal_tmp_2);
  assign IDX_LOOP_f1_or_84_nl = (IDX_LOOP_f2_IDX_LOOP_f2_nor_21_itm & IDX_LOOP_f1_equal_tmp_2)
      | (IDX_LOOP_f2_IDX_LOOP_f2_nor_21_itm & IDX_LOOP_f1_equal_tmp_3) | (IDX_LOOP_f2_IDX_LOOP_f2_nor_21_itm
      & IDX_LOOP_f1_equal_tmp) | (IDX_LOOP_f2_IDX_LOOP_f2_nor_21_itm & IDX_LOOP_f1_equal_tmp_1);
  assign IDX_LOOP_f1_or_85_nl = (IDX_LOOP_f2_IDX_LOOP_f2_nor_28_itm & IDX_LOOP_f1_equal_tmp_1)
      | (IDX_LOOP_f2_IDX_LOOP_f2_nor_28_itm & IDX_LOOP_f1_equal_tmp_2) | (IDX_LOOP_f2_IDX_LOOP_f2_nor_28_itm
      & IDX_LOOP_f1_equal_tmp_3) | (IDX_LOOP_f2_IDX_LOOP_f2_nor_28_itm & IDX_LOOP_f1_equal_tmp);
  assign IDX_LOOP_f1_mux1h_209_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_or_82_nl, IDX_LOOP_f1_or_83_nl,
      IDX_LOOP_f1_or_84_nl, IDX_LOOP_f1_or_85_nl, {and_dcpl_571 , and_dcpl_574 ,
      and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_224_nl = (IDX_LOOP_idx2_9_0_2_sva[0]) & IDX_LOOP_f2_nor_12_cse_1
      & IDX_LOOP_f1_equal_tmp;
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_225_nl = (IDX_LOOP_idx2_9_0_4_sva[0]) & IDX_LOOP_f2_nor_36_cse_1
      & IDX_LOOP_f1_equal_tmp_3;
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_226_nl = (IDX_LOOP_idx2_9_0_6_sva[0]) & IDX_LOOP_f2_nor_60_cse_1
      & IDX_LOOP_f1_equal_tmp_2;
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_227_nl = (IDX_LOOP_idx2_9_0_sva[0]) & IDX_LOOP_f2_nor_84_cse_1
      & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f1_mux1h_210_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_224_nl,
      IDX_LOOP_f2_IDX_LOOP_f2_and_225_nl, IDX_LOOP_f2_IDX_LOOP_f2_and_226_nl, IDX_LOOP_f2_IDX_LOOP_f2_and_227_nl,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_or_86_nl = ((IDX_LOOP_idx2_9_0_2_sva[1]) & IDX_LOOP_f2_nor_13_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_9_0_2_sva[1]) & IDX_LOOP_f2_nor_13_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_9_0_2_sva[1]) & IDX_LOOP_f2_nor_13_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_9_0_2_sva[1]) & IDX_LOOP_f2_nor_13_cse_1
      & IDX_LOOP_f1_equal_tmp_3);
  assign IDX_LOOP_f1_or_87_nl = ((IDX_LOOP_idx2_9_0_4_sva[1]) & IDX_LOOP_f2_nor_37_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_9_0_4_sva[1]) & IDX_LOOP_f2_nor_37_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_9_0_4_sva[1]) & IDX_LOOP_f2_nor_37_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_9_0_4_sva[1]) & IDX_LOOP_f2_nor_37_cse_1
      & IDX_LOOP_f1_equal_tmp_2);
  assign IDX_LOOP_f1_or_88_nl = ((IDX_LOOP_idx2_9_0_6_sva[1]) & IDX_LOOP_f2_nor_61_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_9_0_6_sva[1]) & IDX_LOOP_f2_nor_61_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_9_0_6_sva[1]) & IDX_LOOP_f2_nor_61_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_9_0_6_sva[1]) & IDX_LOOP_f2_nor_61_cse_1
      & IDX_LOOP_f1_equal_tmp_1);
  assign IDX_LOOP_f1_or_89_nl = ((IDX_LOOP_idx2_9_0_sva[1]) & IDX_LOOP_f2_nor_85_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_9_0_sva[1]) & IDX_LOOP_f2_nor_85_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_9_0_sva[1]) & IDX_LOOP_f2_nor_85_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_9_0_sva[1]) & IDX_LOOP_f2_nor_85_cse_1
      & IDX_LOOP_f1_equal_tmp);
  assign IDX_LOOP_f1_mux1h_211_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_or_86_nl, IDX_LOOP_f1_or_87_nl,
      IDX_LOOP_f1_or_88_nl, IDX_LOOP_f1_or_89_nl, {and_dcpl_571 , and_dcpl_574 ,
      and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_mux1h_212_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_30_itm,
      IDX_LOOP_f2_IDX_LOOP_f2_and_86_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_142_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_198_itm,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_or_90_nl = ((IDX_LOOP_idx2_9_0_2_sva[2]) & IDX_LOOP_f2_nor_14_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_9_0_2_sva[2]) & IDX_LOOP_f2_nor_14_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_9_0_2_sva[2]) & IDX_LOOP_f2_nor_14_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_9_0_2_sva[2]) & IDX_LOOP_f2_nor_14_cse_1
      & IDX_LOOP_f1_equal_tmp_3);
  assign IDX_LOOP_f1_or_91_nl = ((IDX_LOOP_idx2_9_0_4_sva[2]) & IDX_LOOP_f2_nor_38_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_9_0_4_sva[2]) & IDX_LOOP_f2_nor_38_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_9_0_4_sva[2]) & IDX_LOOP_f2_nor_38_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_9_0_4_sva[2]) & IDX_LOOP_f2_nor_38_cse_1
      & IDX_LOOP_f1_equal_tmp_2);
  assign IDX_LOOP_f1_or_92_nl = ((IDX_LOOP_idx2_9_0_6_sva[2]) & IDX_LOOP_f2_nor_62_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_9_0_6_sva[2]) & IDX_LOOP_f2_nor_62_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_9_0_6_sva[2]) & IDX_LOOP_f2_nor_62_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_9_0_6_sva[2]) & IDX_LOOP_f2_nor_62_cse_1
      & IDX_LOOP_f1_equal_tmp_1);
  assign IDX_LOOP_f1_or_93_nl = ((IDX_LOOP_idx2_9_0_sva[2]) & IDX_LOOP_f2_nor_86_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_9_0_sva[2]) & IDX_LOOP_f2_nor_86_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_9_0_sva[2]) & IDX_LOOP_f2_nor_86_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_9_0_sva[2]) & IDX_LOOP_f2_nor_86_cse_1
      & IDX_LOOP_f1_equal_tmp);
  assign IDX_LOOP_f1_mux1h_213_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_or_90_nl, IDX_LOOP_f1_or_91_nl,
      IDX_LOOP_f1_or_92_nl, IDX_LOOP_f1_or_93_nl, {and_dcpl_571 , and_dcpl_574 ,
      and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_mux1h_214_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_32_itm,
      IDX_LOOP_f2_IDX_LOOP_f2_and_88_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_144_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_200_itm,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_or_94_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_33_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_40_itm
      | IDX_LOOP_f2_IDX_LOOP_f2_and_47_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_54_itm;
  assign IDX_LOOP_f1_or_95_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_89_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_96_itm
      | IDX_LOOP_f2_IDX_LOOP_f2_and_103_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_110_itm;
  assign IDX_LOOP_f1_or_96_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_145_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_152_itm
      | IDX_LOOP_f2_IDX_LOOP_f2_and_159_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_166_itm;
  assign IDX_LOOP_f1_or_97_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_201_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_208_itm
      | IDX_LOOP_IDX_LOOP_and_104_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_222_itm;
  assign IDX_LOOP_f1_mux1h_215_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_or_94_nl, IDX_LOOP_f1_or_95_nl,
      IDX_LOOP_f1_or_96_nl, IDX_LOOP_f1_or_97_nl, {and_dcpl_571 , and_dcpl_574 ,
      and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_mux1h_216_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_34_itm,
      IDX_LOOP_f2_IDX_LOOP_f2_and_90_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_146_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_202_itm,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_260_nl = (IDX_LOOP_idx2_9_0_2_sva[0]) & IDX_LOOP_f2_nor_12_cse_1
      & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_261_nl = (IDX_LOOP_idx2_9_0_4_sva[0]) & IDX_LOOP_f2_nor_36_cse_1
      & IDX_LOOP_f1_equal_tmp;
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_262_nl = (IDX_LOOP_idx2_9_0_6_sva[0]) & IDX_LOOP_f2_nor_60_cse_1
      & IDX_LOOP_f1_equal_tmp_3;
  assign IDX_LOOP_f2_IDX_LOOP_f2_and_263_nl = (IDX_LOOP_idx2_9_0_sva[0]) & IDX_LOOP_f2_nor_84_cse_1
      & IDX_LOOP_f1_equal_tmp_2;
  assign IDX_LOOP_f1_mux1h_217_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_260_nl,
      IDX_LOOP_f2_IDX_LOOP_f2_and_261_nl, IDX_LOOP_f2_IDX_LOOP_f2_and_262_nl, IDX_LOOP_f2_IDX_LOOP_f2_and_263_nl,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_mux1h_218_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_37_itm,
      IDX_LOOP_f2_IDX_LOOP_f2_and_93_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_149_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_205_itm,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_mux1h_219_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_39_itm,
      IDX_LOOP_f2_IDX_LOOP_f2_and_95_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_151_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_207_itm,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_or_98_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_41_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_48_itm;
  assign IDX_LOOP_f1_or_99_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_97_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_104_itm;
  assign IDX_LOOP_f1_or_100_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_153_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_160_itm;
  assign IDX_LOOP_f1_or_101_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_209_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_216_itm;
  assign IDX_LOOP_f1_mux1h_220_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_or_98_nl, IDX_LOOP_f1_or_99_nl,
      IDX_LOOP_f1_or_100_nl, IDX_LOOP_f1_or_101_nl, {and_dcpl_571 , and_dcpl_574
      , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_or_102_nl = ((IDX_LOOP_idx2_9_0_2_sva[0]) & IDX_LOOP_f2_nor_12_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_9_0_2_sva[0]) & IDX_LOOP_f2_nor_12_cse_1
      & IDX_LOOP_f1_equal_tmp_3);
  assign IDX_LOOP_f1_or_103_nl = ((IDX_LOOP_idx2_9_0_4_sva[0]) & IDX_LOOP_f2_nor_36_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_9_0_4_sva[0]) & IDX_LOOP_f2_nor_36_cse_1
      & IDX_LOOP_f1_equal_tmp_2);
  assign IDX_LOOP_f1_or_104_nl = ((IDX_LOOP_idx2_9_0_6_sva[0]) & IDX_LOOP_f2_nor_60_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_9_0_6_sva[0]) & IDX_LOOP_f2_nor_60_cse_1
      & IDX_LOOP_f1_equal_tmp_1);
  assign IDX_LOOP_f1_or_105_nl = ((IDX_LOOP_idx2_9_0_sva[0]) & IDX_LOOP_f2_nor_84_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_9_0_sva[0]) & IDX_LOOP_f2_nor_84_cse_1
      & IDX_LOOP_f1_equal_tmp);
  assign IDX_LOOP_f1_mux1h_221_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_or_102_nl, IDX_LOOP_f1_or_103_nl,
      IDX_LOOP_f1_or_104_nl, IDX_LOOP_f1_or_105_nl, {and_dcpl_571 , and_dcpl_574
      , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_or_106_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_44_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_51_itm;
  assign IDX_LOOP_f1_or_107_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_100_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_107_itm;
  assign IDX_LOOP_f1_or_108_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_156_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_163_itm;
  assign IDX_LOOP_f1_or_109_nl = IDX_LOOP_f2_IDX_LOOP_f2_and_212_itm | IDX_LOOP_f2_IDX_LOOP_f2_and_219_itm;
  assign IDX_LOOP_f1_mux1h_222_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f1_or_106_nl, IDX_LOOP_f1_or_107_nl,
      IDX_LOOP_f1_or_108_nl, IDX_LOOP_f1_or_109_nl, {and_dcpl_571 , and_dcpl_574
      , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_mux1h_223_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_46_itm,
      IDX_LOOP_f2_IDX_LOOP_f2_and_102_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_158_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_214_itm,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_mux1h_224_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_53_itm,
      IDX_LOOP_f2_IDX_LOOP_f2_and_109_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_165_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_221_itm,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign IDX_LOOP_f1_mux1h_225_nl = MUX1HOT_s_1_4_2(IDX_LOOP_f2_IDX_LOOP_f2_and_55_itm,
      IDX_LOOP_f2_IDX_LOOP_f2_and_111_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_167_itm, IDX_LOOP_f2_IDX_LOOP_f2_and_223_itm,
      {and_dcpl_571 , and_dcpl_574 , and_dcpl_577 , and_dcpl_579});
  assign z_out_7 = MUX1HOT_v_64_17_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d, vec_rsc_0_2_i_q_d,
      tmp_11_sva_3, vec_rsc_0_4_i_q_d, tmp_11_sva_5, vec_rsc_0_6_i_q_d, tmp_11_sva_7,
      tmp_11_sva_9, vec_rsc_0_3_i_q_d, IDX_LOOP_modulo_dev_return_1_sva, reg_cse,
      reg_1_cse, reg_2_cse, vec_rsc_0_5_i_q_d, tmp_11_sva_29, vec_rsc_0_7_i_q_d,
      {IDX_LOOP_f1_mux1h_209_nl , IDX_LOOP_f1_mux1h_210_nl , IDX_LOOP_f1_mux1h_211_nl
      , IDX_LOOP_f1_mux1h_212_nl , IDX_LOOP_f1_mux1h_213_nl , IDX_LOOP_f1_mux1h_214_nl
      , IDX_LOOP_f1_mux1h_215_nl , IDX_LOOP_f1_mux1h_216_nl , IDX_LOOP_f1_mux1h_217_nl
      , IDX_LOOP_f1_mux1h_218_nl , IDX_LOOP_f1_mux1h_219_nl , IDX_LOOP_f1_mux1h_220_nl
      , IDX_LOOP_f1_mux1h_221_nl , IDX_LOOP_f1_mux1h_222_nl , IDX_LOOP_f1_mux1h_223_nl
      , IDX_LOOP_f1_mux1h_224_nl , IDX_LOOP_f1_mux1h_225_nl});
  assign IDX_LOOP_f1_and_160_nl = IDX_LOOP_f2_IDX_LOOP_f2_nor_8_itm & IDX_LOOP_f1_equal_tmp_3;
  assign IDX_LOOP_f1_and_161_nl = IDX_LOOP_f2_IDX_LOOP_f2_nor_16_itm & IDX_LOOP_f1_equal_tmp_2;
  assign IDX_LOOP_f1_and_162_nl = IDX_LOOP_f2_IDX_LOOP_f2_nor_24_itm & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f1_mux1h_226_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_and_160_nl, IDX_LOOP_f1_and_161_nl,
      IDX_LOOP_f1_and_162_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_or_110_nl = ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_24_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_24_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_24_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_24_cse_1
      & IDX_LOOP_f1_equal_tmp_2);
  assign IDX_LOOP_f1_or_111_nl = ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_48_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_48_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_48_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_48_cse_1
      & IDX_LOOP_f1_equal_tmp_1);
  assign IDX_LOOP_f1_or_112_nl = ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_72_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_72_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_72_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((STAGE_LOOP_op_rshift_psp_1_sva[0]) & IDX_LOOP_f2_nor_72_cse_1
      & IDX_LOOP_f1_equal_tmp);
  assign IDX_LOOP_f1_mux1h_227_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_or_110_nl, IDX_LOOP_f1_or_111_nl,
      IDX_LOOP_f1_or_112_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_or_113_nl = ((IDX_LOOP_idx2_acc_1_psp_sva[0]) & IDX_LOOP_f2_nor_25_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_acc_1_psp_sva[1]) & IDX_LOOP_f2_nor_26_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_acc_1_psp_sva[1]) & IDX_LOOP_f2_nor_26_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_acc_1_psp_sva[0]) & IDX_LOOP_f2_nor_25_cse_1
      & IDX_LOOP_f1_equal_tmp_2);
  assign IDX_LOOP_f1_or_114_nl = ((IDX_LOOP_idx2_acc_2_psp_sva[0]) & IDX_LOOP_f2_nor_49_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_acc_2_psp_sva[1]) & IDX_LOOP_f2_nor_50_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_acc_2_psp_sva[1]) & IDX_LOOP_f2_nor_50_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_acc_2_psp_sva[0]) & IDX_LOOP_f2_nor_49_cse_1
      & IDX_LOOP_f1_equal_tmp_1);
  assign IDX_LOOP_f1_or_115_nl = ((IDX_LOOP_idx2_acc_3_psp_sva[0]) & IDX_LOOP_f2_nor_73_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_acc_3_psp_sva[1]) & IDX_LOOP_f2_nor_74_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_acc_3_psp_sva[1]) & IDX_LOOP_f2_nor_74_cse_1
      & IDX_LOOP_f1_equal_tmp_1) | ((IDX_LOOP_idx2_acc_3_psp_sva[0]) & IDX_LOOP_f2_nor_73_cse_1
      & IDX_LOOP_f1_equal_tmp);
  assign IDX_LOOP_f1_mux1h_228_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_or_113_nl, IDX_LOOP_f1_or_114_nl,
      IDX_LOOP_f1_or_115_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_or_116_nl = IDX_LOOP_f1_and_39_itm | IDX_LOOP_f1_and_47_itm
      | IDX_LOOP_f1_and_55_itm | IDX_LOOP_f1_and_63_itm;
  assign IDX_LOOP_f1_or_117_nl = IDX_LOOP_f1_and_75_itm | IDX_LOOP_f1_and_83_itm
      | IDX_LOOP_f1_and_91_itm | IDX_LOOP_f1_and_99_itm;
  assign IDX_LOOP_f1_or_118_nl = IDX_LOOP_f1_and_111_itm | IDX_LOOP_f1_and_119_itm
      | IDX_LOOP_f1_and_127_itm | IDX_LOOP_f1_and_135_itm;
  assign IDX_LOOP_f1_mux1h_229_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_or_116_nl, IDX_LOOP_f1_or_117_nl,
      IDX_LOOP_f1_or_118_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_or_119_nl = IDX_LOOP_f1_and_41_itm | IDX_LOOP_f1_and_49_itm
      | IDX_LOOP_f1_and_57_itm | IDX_LOOP_f1_and_65_itm;
  assign IDX_LOOP_f1_or_120_nl = IDX_LOOP_f1_and_77_itm | IDX_LOOP_f1_and_85_itm
      | IDX_LOOP_f1_and_93_itm | IDX_LOOP_f1_and_101_itm;
  assign IDX_LOOP_f1_or_121_nl = IDX_LOOP_f1_and_113_itm | IDX_LOOP_f1_and_121_itm
      | IDX_LOOP_f1_and_129_itm | IDX_LOOP_f1_and_137_itm;
  assign IDX_LOOP_f1_mux1h_230_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_or_119_nl, IDX_LOOP_f1_or_120_nl,
      IDX_LOOP_f1_or_121_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_mux1h_231_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_and_42_itm, IDX_LOOP_f1_and_78_itm,
      IDX_LOOP_f1_and_114_itm, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_or_122_nl = IDX_LOOP_f1_and_43_itm | IDX_LOOP_f1_and_51_itm
      | IDX_LOOP_f1_and_59_itm | IDX_LOOP_f1_and_67_itm;
  assign IDX_LOOP_f1_or_123_nl = IDX_LOOP_f1_and_79_itm | IDX_LOOP_f1_and_87_itm
      | IDX_LOOP_f1_and_95_itm | IDX_LOOP_f1_and_103_itm;
  assign IDX_LOOP_f1_or_124_nl = IDX_LOOP_f1_and_115_itm | IDX_LOOP_f1_and_123_itm
      | IDX_LOOP_f1_and_131_itm | IDX_LOOP_f1_and_139_itm;
  assign IDX_LOOP_f1_mux1h_232_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_or_122_nl, IDX_LOOP_f1_or_123_nl,
      IDX_LOOP_f1_or_124_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_and_187_nl = IDX_LOOP_f2_IDX_LOOP_f2_nor_8_itm & IDX_LOOP_f1_equal_tmp;
  assign IDX_LOOP_f1_and_188_nl = IDX_LOOP_f2_IDX_LOOP_f2_nor_16_itm & IDX_LOOP_f1_equal_tmp_3;
  assign IDX_LOOP_f1_and_189_nl = IDX_LOOP_f2_IDX_LOOP_f2_nor_24_itm & IDX_LOOP_f1_equal_tmp_2;
  assign IDX_LOOP_f1_mux1h_233_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_and_187_nl, IDX_LOOP_f1_and_188_nl,
      IDX_LOOP_f1_and_189_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_and_190_nl = (IDX_LOOP_idx2_acc_1_psp_sva[0]) & IDX_LOOP_f2_nor_25_cse_1
      & IDX_LOOP_f1_equal_tmp;
  assign IDX_LOOP_f1_and_191_nl = (IDX_LOOP_idx2_acc_2_psp_sva[0]) & IDX_LOOP_f2_nor_49_cse_1
      & IDX_LOOP_f1_equal_tmp_3;
  assign IDX_LOOP_f1_and_192_nl = (IDX_LOOP_idx2_acc_3_psp_sva[0]) & IDX_LOOP_f2_nor_73_cse_1
      & IDX_LOOP_f1_equal_tmp_2;
  assign IDX_LOOP_f1_mux1h_234_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_and_190_nl, IDX_LOOP_f1_and_191_nl,
      IDX_LOOP_f1_and_192_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_or_125_nl = ((IDX_LOOP_idx2_acc_1_psp_sva[1]) & IDX_LOOP_f2_nor_26_cse_1
      & IDX_LOOP_f1_equal_tmp) | ((IDX_LOOP_idx2_acc_1_psp_sva[0]) & IDX_LOOP_f2_nor_25_cse_1
      & IDX_LOOP_f1_equal_tmp_1);
  assign IDX_LOOP_f1_or_126_nl = ((IDX_LOOP_idx2_acc_2_psp_sva[1]) & IDX_LOOP_f2_nor_50_cse_1
      & IDX_LOOP_f1_equal_tmp_3) | ((IDX_LOOP_idx2_acc_2_psp_sva[0]) & IDX_LOOP_f2_nor_49_cse_1
      & IDX_LOOP_f1_equal_tmp);
  assign IDX_LOOP_f1_or_127_nl = ((IDX_LOOP_idx2_acc_3_psp_sva[1]) & IDX_LOOP_f2_nor_74_cse_1
      & IDX_LOOP_f1_equal_tmp_2) | ((IDX_LOOP_idx2_acc_3_psp_sva[0]) & IDX_LOOP_f2_nor_73_cse_1
      & IDX_LOOP_f1_equal_tmp_3);
  assign IDX_LOOP_f1_mux1h_235_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_or_125_nl, IDX_LOOP_f1_or_126_nl,
      IDX_LOOP_f1_or_127_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_or_128_nl = IDX_LOOP_f1_and_50_itm | IDX_LOOP_f1_and_58_itm;
  assign IDX_LOOP_f1_or_129_nl = IDX_LOOP_f1_and_86_itm | IDX_LOOP_f1_and_94_itm;
  assign IDX_LOOP_f1_or_130_nl = IDX_LOOP_f1_and_122_itm | IDX_LOOP_f1_and_130_itm;
  assign IDX_LOOP_f1_mux1h_236_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_or_128_nl, IDX_LOOP_f1_or_129_nl,
      IDX_LOOP_f1_or_130_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_or_131_nl = (IDX_LOOP_f2_IDX_LOOP_f2_nor_8_itm & IDX_LOOP_f1_equal_tmp_1)
      | (IDX_LOOP_f2_IDX_LOOP_f2_nor_8_itm & IDX_LOOP_f1_equal_tmp_2);
  assign IDX_LOOP_f1_or_132_nl = (IDX_LOOP_f2_IDX_LOOP_f2_nor_16_itm & IDX_LOOP_f1_equal_tmp)
      | (IDX_LOOP_f2_IDX_LOOP_f2_nor_16_itm & IDX_LOOP_f1_equal_tmp_1);
  assign IDX_LOOP_f1_or_133_nl = (IDX_LOOP_f2_IDX_LOOP_f2_nor_24_itm & IDX_LOOP_f1_equal_tmp_3)
      | (IDX_LOOP_f2_IDX_LOOP_f2_nor_24_itm & IDX_LOOP_f1_equal_tmp);
  assign IDX_LOOP_f1_mux1h_237_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_or_131_nl, IDX_LOOP_f1_or_132_nl,
      IDX_LOOP_f1_or_133_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_and_205_nl = (IDX_LOOP_idx2_acc_1_psp_sva[1]) & IDX_LOOP_f2_nor_26_cse_1
      & IDX_LOOP_f1_equal_tmp_1;
  assign IDX_LOOP_f1_and_206_nl = (IDX_LOOP_idx2_acc_2_psp_sva[1]) & IDX_LOOP_f2_nor_50_cse_1
      & IDX_LOOP_f1_equal_tmp;
  assign IDX_LOOP_f1_and_207_nl = (IDX_LOOP_idx2_acc_3_psp_sva[1]) & IDX_LOOP_f2_nor_74_cse_1
      & IDX_LOOP_f1_equal_tmp_3;
  assign IDX_LOOP_f1_mux1h_238_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_and_205_nl, IDX_LOOP_f1_and_206_nl,
      IDX_LOOP_f1_and_207_nl, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign IDX_LOOP_f1_mux1h_239_nl = MUX1HOT_s_1_3_2(IDX_LOOP_f1_and_66_itm, IDX_LOOP_f1_and_102_itm,
      IDX_LOOP_f1_and_138_itm, {and_dcpl_587 , and_dcpl_591 , and_dcpl_593});
  assign z_out_8 = MUX1HOT_v_64_14_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d, reg_2_cse,
      vec_rsc_0_3_i_q_d, vec_rsc_0_5_i_q_d, tmp_11_sva_29, vec_rsc_0_7_i_q_d, tmp_11_sva_3,
      vec_rsc_0_2_i_q_d, IDX_LOOP_modulo_dev_return_1_sva, reg_cse, reg_1_cse, vec_rsc_0_4_i_q_d,
      vec_rsc_0_6_i_q_d, {IDX_LOOP_f1_mux1h_226_nl , IDX_LOOP_f1_mux1h_227_nl , IDX_LOOP_f1_mux1h_228_nl
      , IDX_LOOP_f1_mux1h_229_nl , IDX_LOOP_f1_mux1h_230_nl , IDX_LOOP_f1_mux1h_231_nl
      , IDX_LOOP_f1_mux1h_232_nl , IDX_LOOP_f1_mux1h_233_nl , IDX_LOOP_f1_mux1h_234_nl
      , IDX_LOOP_f1_mux1h_235_nl , IDX_LOOP_f1_mux1h_236_nl , IDX_LOOP_f1_mux1h_237_nl
      , IDX_LOOP_f1_mux1h_238_nl , IDX_LOOP_f1_mux1h_239_nl});

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_11_2;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [10:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    MUX1HOT_v_64_11_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_14_2;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [13:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    MUX1HOT_v_64_14_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_17_2;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [16:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    MUX1HOT_v_64_17_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_5_2;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [4:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    MUX1HOT_v_64_5_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_8_2;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [7:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    MUX1HOT_v_64_8_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_12_2;
    input [6:0] input_11;
    input [6:0] input_10;
    input [6:0] input_9;
    input [6:0] input_8;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [11:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    result = result | ( input_4 & {7{sel[4]}});
    result = result | ( input_5 & {7{sel[5]}});
    result = result | ( input_6 & {7{sel[6]}});
    result = result | ( input_7 & {7{sel[7]}});
    result = result | ( input_8 & {7{sel[8]}});
    result = result | ( input_9 & {7{sel[9]}});
    result = result | ( input_10 & {7{sel[10]}});
    result = result | ( input_11 & {7{sel[11]}});
    MUX1HOT_v_7_12_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] readslicef_12_11_1;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_12_11_1 = tmp[10:0];
  end
  endfunction


  function automatic [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [63:0] readslicef_65_64_1;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_65_64_1 = tmp[63:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [7:0] conv_s2u_2_8 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_8 = {{6{vector[1]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction


  function automatic [127:0] conv_u2u_128_128 ;
    input [127:0]  vector ;
  begin
    conv_u2u_128_128 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    DIT_RELOOP
// ------------------------------------------------------------------


module DIT_RELOOP (
  clk, rst, vec_rsc_0_0_radr, vec_rsc_0_0_re, vec_rsc_0_0_q, vec_rsc_0_0_wadr, vec_rsc_0_0_d,
      vec_rsc_0_0_we, vec_rsc_triosy_0_0_lz, vec_rsc_0_1_radr, vec_rsc_0_1_re, vec_rsc_0_1_q,
      vec_rsc_0_1_wadr, vec_rsc_0_1_d, vec_rsc_0_1_we, vec_rsc_triosy_0_1_lz, vec_rsc_0_2_radr,
      vec_rsc_0_2_re, vec_rsc_0_2_q, vec_rsc_0_2_wadr, vec_rsc_0_2_d, vec_rsc_0_2_we,
      vec_rsc_triosy_0_2_lz, vec_rsc_0_3_radr, vec_rsc_0_3_re, vec_rsc_0_3_q, vec_rsc_0_3_wadr,
      vec_rsc_0_3_d, vec_rsc_0_3_we, vec_rsc_triosy_0_3_lz, vec_rsc_0_4_radr, vec_rsc_0_4_re,
      vec_rsc_0_4_q, vec_rsc_0_4_wadr, vec_rsc_0_4_d, vec_rsc_0_4_we, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_radr, vec_rsc_0_5_re, vec_rsc_0_5_q, vec_rsc_0_5_wadr, vec_rsc_0_5_d,
      vec_rsc_0_5_we, vec_rsc_triosy_0_5_lz, vec_rsc_0_6_radr, vec_rsc_0_6_re, vec_rsc_0_6_q,
      vec_rsc_0_6_wadr, vec_rsc_0_6_d, vec_rsc_0_6_we, vec_rsc_triosy_0_6_lz, vec_rsc_0_7_radr,
      vec_rsc_0_7_re, vec_rsc_0_7_q, vec_rsc_0_7_wadr, vec_rsc_0_7_d, vec_rsc_0_7_we,
      vec_rsc_triosy_0_7_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      twiddle_rsc_0_0_radr, twiddle_rsc_0_0_re, twiddle_rsc_0_0_q, twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_0_1_radr, twiddle_rsc_0_1_re, twiddle_rsc_0_1_q, twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_0_2_radr, twiddle_rsc_0_2_re, twiddle_rsc_0_2_q, twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_0_3_radr, twiddle_rsc_0_3_re, twiddle_rsc_0_3_q, twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_0_4_radr, twiddle_rsc_0_4_re, twiddle_rsc_0_4_q, twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_0_5_radr, twiddle_rsc_0_5_re, twiddle_rsc_0_5_q, twiddle_rsc_triosy_0_5_lz,
      twiddle_rsc_0_6_radr, twiddle_rsc_0_6_re, twiddle_rsc_0_6_q, twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_0_7_radr, twiddle_rsc_0_7_re, twiddle_rsc_0_7_q, twiddle_rsc_triosy_0_7_lz
);
  input clk;
  input rst;
  output [6:0] vec_rsc_0_0_radr;
  output vec_rsc_0_0_re;
  input [63:0] vec_rsc_0_0_q;
  output [6:0] vec_rsc_0_0_wadr;
  output [63:0] vec_rsc_0_0_d;
  output vec_rsc_0_0_we;
  output vec_rsc_triosy_0_0_lz;
  output [6:0] vec_rsc_0_1_radr;
  output vec_rsc_0_1_re;
  input [63:0] vec_rsc_0_1_q;
  output [6:0] vec_rsc_0_1_wadr;
  output [63:0] vec_rsc_0_1_d;
  output vec_rsc_0_1_we;
  output vec_rsc_triosy_0_1_lz;
  output [6:0] vec_rsc_0_2_radr;
  output vec_rsc_0_2_re;
  input [63:0] vec_rsc_0_2_q;
  output [6:0] vec_rsc_0_2_wadr;
  output [63:0] vec_rsc_0_2_d;
  output vec_rsc_0_2_we;
  output vec_rsc_triosy_0_2_lz;
  output [6:0] vec_rsc_0_3_radr;
  output vec_rsc_0_3_re;
  input [63:0] vec_rsc_0_3_q;
  output [6:0] vec_rsc_0_3_wadr;
  output [63:0] vec_rsc_0_3_d;
  output vec_rsc_0_3_we;
  output vec_rsc_triosy_0_3_lz;
  output [6:0] vec_rsc_0_4_radr;
  output vec_rsc_0_4_re;
  input [63:0] vec_rsc_0_4_q;
  output [6:0] vec_rsc_0_4_wadr;
  output [63:0] vec_rsc_0_4_d;
  output vec_rsc_0_4_we;
  output vec_rsc_triosy_0_4_lz;
  output [6:0] vec_rsc_0_5_radr;
  output vec_rsc_0_5_re;
  input [63:0] vec_rsc_0_5_q;
  output [6:0] vec_rsc_0_5_wadr;
  output [63:0] vec_rsc_0_5_d;
  output vec_rsc_0_5_we;
  output vec_rsc_triosy_0_5_lz;
  output [6:0] vec_rsc_0_6_radr;
  output vec_rsc_0_6_re;
  input [63:0] vec_rsc_0_6_q;
  output [6:0] vec_rsc_0_6_wadr;
  output [63:0] vec_rsc_0_6_d;
  output vec_rsc_0_6_we;
  output vec_rsc_triosy_0_6_lz;
  output [6:0] vec_rsc_0_7_radr;
  output vec_rsc_0_7_re;
  input [63:0] vec_rsc_0_7_q;
  output [6:0] vec_rsc_0_7_wadr;
  output [63:0] vec_rsc_0_7_d;
  output vec_rsc_0_7_we;
  output vec_rsc_triosy_0_7_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  output [6:0] twiddle_rsc_0_0_radr;
  output twiddle_rsc_0_0_re;
  input [63:0] twiddle_rsc_0_0_q;
  output twiddle_rsc_triosy_0_0_lz;
  output [6:0] twiddle_rsc_0_1_radr;
  output twiddle_rsc_0_1_re;
  input [63:0] twiddle_rsc_0_1_q;
  output twiddle_rsc_triosy_0_1_lz;
  output [6:0] twiddle_rsc_0_2_radr;
  output twiddle_rsc_0_2_re;
  input [63:0] twiddle_rsc_0_2_q;
  output twiddle_rsc_triosy_0_2_lz;
  output [6:0] twiddle_rsc_0_3_radr;
  output twiddle_rsc_0_3_re;
  input [63:0] twiddle_rsc_0_3_q;
  output twiddle_rsc_triosy_0_3_lz;
  output [6:0] twiddle_rsc_0_4_radr;
  output twiddle_rsc_0_4_re;
  input [63:0] twiddle_rsc_0_4_q;
  output twiddle_rsc_triosy_0_4_lz;
  output [6:0] twiddle_rsc_0_5_radr;
  output twiddle_rsc_0_5_re;
  input [63:0] twiddle_rsc_0_5_q;
  output twiddle_rsc_triosy_0_5_lz;
  output [6:0] twiddle_rsc_0_6_radr;
  output twiddle_rsc_0_6_re;
  input [63:0] twiddle_rsc_0_6_q;
  output twiddle_rsc_triosy_0_6_lz;
  output [6:0] twiddle_rsc_0_7_radr;
  output twiddle_rsc_0_7_re;
  input [63:0] twiddle_rsc_0_7_q;
  output twiddle_rsc_triosy_0_7_lz;


  // Interconnect Declarations
  wire [6:0] vec_rsc_0_0_i_radr_d;
  wire [63:0] vec_rsc_0_0_i_q_d;
  wire [6:0] vec_rsc_0_1_i_radr_d;
  wire [63:0] vec_rsc_0_1_i_q_d;
  wire [6:0] vec_rsc_0_2_i_radr_d;
  wire [63:0] vec_rsc_0_2_i_q_d;
  wire [6:0] vec_rsc_0_3_i_radr_d;
  wire [63:0] vec_rsc_0_3_i_q_d;
  wire [6:0] vec_rsc_0_4_i_radr_d;
  wire [63:0] vec_rsc_0_4_i_q_d;
  wire [6:0] vec_rsc_0_5_i_radr_d;
  wire [63:0] vec_rsc_0_5_i_q_d;
  wire [6:0] vec_rsc_0_6_i_radr_d;
  wire [63:0] vec_rsc_0_6_i_q_d;
  wire [6:0] vec_rsc_0_7_i_radr_d;
  wire [63:0] vec_rsc_0_7_i_q_d;
  wire [63:0] twiddle_rsc_0_0_i_q_d;
  wire [63:0] twiddle_rsc_0_1_i_q_d;
  wire [63:0] twiddle_rsc_0_2_i_q_d;
  wire [63:0] twiddle_rsc_0_3_i_q_d;
  wire [63:0] twiddle_rsc_0_4_i_q_d;
  wire [63:0] twiddle_rsc_0_5_i_q_d;
  wire [63:0] twiddle_rsc_0_6_i_q_d;
  wire [63:0] twiddle_rsc_0_7_i_q_d;
  wire [6:0] vec_rsc_0_0_i_wadr_d_iff;
  wire [63:0] vec_rsc_0_0_i_d_d_iff;
  wire vec_rsc_0_0_i_we_d_iff;
  wire vec_rsc_0_0_i_re_d_iff;
  wire [6:0] vec_rsc_0_1_i_wadr_d_iff;
  wire [63:0] vec_rsc_0_1_i_d_d_iff;
  wire vec_rsc_0_1_i_we_d_iff;
  wire vec_rsc_0_1_i_re_d_iff;
  wire vec_rsc_0_2_i_we_d_iff;
  wire vec_rsc_0_2_i_re_d_iff;
  wire vec_rsc_0_3_i_we_d_iff;
  wire vec_rsc_0_3_i_re_d_iff;
  wire vec_rsc_0_4_i_we_d_iff;
  wire vec_rsc_0_4_i_re_d_iff;
  wire vec_rsc_0_5_i_we_d_iff;
  wire vec_rsc_0_5_i_re_d_iff;
  wire vec_rsc_0_6_i_we_d_iff;
  wire vec_rsc_0_6_i_re_d_iff;
  wire vec_rsc_0_7_i_we_d_iff;
  wire vec_rsc_0_7_i_re_d_iff;
  wire [6:0] twiddle_rsc_0_0_i_radr_d_iff;
  wire twiddle_rsc_0_0_i_re_d_iff;
  wire twiddle_rsc_0_1_i_re_d_iff;
  wire twiddle_rsc_0_2_i_re_d_iff;
  wire twiddle_rsc_0_3_i_re_d_iff;
  wire twiddle_rsc_0_4_i_re_d_iff;
  wire twiddle_rsc_0_5_i_re_d_iff;
  wire twiddle_rsc_0_6_i_re_d_iff;
  wire twiddle_rsc_0_7_i_re_d_iff;


  // Interconnect Declarations for Component Instantiations 
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_9_64_7_128_128_64_5_gen vec_rsc_0_0_i
      (
      .we(vec_rsc_0_0_we),
      .d(vec_rsc_0_0_d),
      .wadr(vec_rsc_0_0_wadr),
      .q(vec_rsc_0_0_q),
      .re(vec_rsc_0_0_re),
      .radr(vec_rsc_0_0_radr),
      .radr_d(vec_rsc_0_0_i_radr_d),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .we_d(vec_rsc_0_0_i_we_d_iff),
      .re_d(vec_rsc_0_0_i_re_d_iff),
      .q_d(vec_rsc_0_0_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_we_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_10_64_7_128_128_64_5_gen vec_rsc_0_1_i
      (
      .we(vec_rsc_0_1_we),
      .d(vec_rsc_0_1_d),
      .wadr(vec_rsc_0_1_wadr),
      .q(vec_rsc_0_1_q),
      .re(vec_rsc_0_1_re),
      .radr(vec_rsc_0_1_radr),
      .radr_d(vec_rsc_0_1_i_radr_d),
      .wadr_d(vec_rsc_0_1_i_wadr_d_iff),
      .d_d(vec_rsc_0_1_i_d_d_iff),
      .we_d(vec_rsc_0_1_i_we_d_iff),
      .re_d(vec_rsc_0_1_i_re_d_iff),
      .q_d(vec_rsc_0_1_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_we_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_11_64_7_128_128_64_5_gen vec_rsc_0_2_i
      (
      .we(vec_rsc_0_2_we),
      .d(vec_rsc_0_2_d),
      .wadr(vec_rsc_0_2_wadr),
      .q(vec_rsc_0_2_q),
      .re(vec_rsc_0_2_re),
      .radr(vec_rsc_0_2_radr),
      .radr_d(vec_rsc_0_2_i_radr_d),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .we_d(vec_rsc_0_2_i_we_d_iff),
      .re_d(vec_rsc_0_2_i_re_d_iff),
      .q_d(vec_rsc_0_2_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_we_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_12_64_7_128_128_64_5_gen vec_rsc_0_3_i
      (
      .we(vec_rsc_0_3_we),
      .d(vec_rsc_0_3_d),
      .wadr(vec_rsc_0_3_wadr),
      .q(vec_rsc_0_3_q),
      .re(vec_rsc_0_3_re),
      .radr(vec_rsc_0_3_radr),
      .radr_d(vec_rsc_0_3_i_radr_d),
      .wadr_d(vec_rsc_0_1_i_wadr_d_iff),
      .d_d(vec_rsc_0_1_i_d_d_iff),
      .we_d(vec_rsc_0_3_i_we_d_iff),
      .re_d(vec_rsc_0_3_i_re_d_iff),
      .q_d(vec_rsc_0_3_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_we_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_13_64_7_128_128_64_5_gen vec_rsc_0_4_i
      (
      .we(vec_rsc_0_4_we),
      .d(vec_rsc_0_4_d),
      .wadr(vec_rsc_0_4_wadr),
      .q(vec_rsc_0_4_q),
      .re(vec_rsc_0_4_re),
      .radr(vec_rsc_0_4_radr),
      .radr_d(vec_rsc_0_4_i_radr_d),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .we_d(vec_rsc_0_4_i_we_d_iff),
      .re_d(vec_rsc_0_4_i_re_d_iff),
      .q_d(vec_rsc_0_4_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_we_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_14_64_7_128_128_64_5_gen vec_rsc_0_5_i
      (
      .we(vec_rsc_0_5_we),
      .d(vec_rsc_0_5_d),
      .wadr(vec_rsc_0_5_wadr),
      .q(vec_rsc_0_5_q),
      .re(vec_rsc_0_5_re),
      .radr(vec_rsc_0_5_radr),
      .radr_d(vec_rsc_0_5_i_radr_d),
      .wadr_d(vec_rsc_0_1_i_wadr_d_iff),
      .d_d(vec_rsc_0_1_i_d_d_iff),
      .we_d(vec_rsc_0_5_i_we_d_iff),
      .re_d(vec_rsc_0_5_i_re_d_iff),
      .q_d(vec_rsc_0_5_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_we_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_15_64_7_128_128_64_5_gen vec_rsc_0_6_i
      (
      .we(vec_rsc_0_6_we),
      .d(vec_rsc_0_6_d),
      .wadr(vec_rsc_0_6_wadr),
      .q(vec_rsc_0_6_q),
      .re(vec_rsc_0_6_re),
      .radr(vec_rsc_0_6_radr),
      .radr_d(vec_rsc_0_6_i_radr_d),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .we_d(vec_rsc_0_6_i_we_d_iff),
      .re_d(vec_rsc_0_6_i_re_d_iff),
      .q_d(vec_rsc_0_6_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_we_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_16_64_7_128_128_64_5_gen vec_rsc_0_7_i
      (
      .we(vec_rsc_0_7_we),
      .d(vec_rsc_0_7_d),
      .wadr(vec_rsc_0_7_wadr),
      .q(vec_rsc_0_7_q),
      .re(vec_rsc_0_7_re),
      .radr(vec_rsc_0_7_radr),
      .radr_d(vec_rsc_0_7_i_radr_d),
      .wadr_d(vec_rsc_0_1_i_wadr_d_iff),
      .d_d(vec_rsc_0_1_i_d_d_iff),
      .we_d(vec_rsc_0_7_i_we_d_iff),
      .re_d(vec_rsc_0_7_i_re_d_iff),
      .q_d(vec_rsc_0_7_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_we_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_17_64_7_128_128_64_5_gen twiddle_rsc_0_0_i
      (
      .q(twiddle_rsc_0_0_q),
      .re(twiddle_rsc_0_0_re),
      .radr(twiddle_rsc_0_0_radr),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .re_d(twiddle_rsc_0_0_i_re_d_iff),
      .q_d(twiddle_rsc_0_0_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_re_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_18_64_7_128_128_64_5_gen twiddle_rsc_0_1_i
      (
      .q(twiddle_rsc_0_1_q),
      .re(twiddle_rsc_0_1_re),
      .radr(twiddle_rsc_0_1_radr),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .re_d(twiddle_rsc_0_1_i_re_d_iff),
      .q_d(twiddle_rsc_0_1_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_re_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_19_64_7_128_128_64_5_gen twiddle_rsc_0_2_i
      (
      .q(twiddle_rsc_0_2_q),
      .re(twiddle_rsc_0_2_re),
      .radr(twiddle_rsc_0_2_radr),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .re_d(twiddle_rsc_0_2_i_re_d_iff),
      .q_d(twiddle_rsc_0_2_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_re_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_20_64_7_128_128_64_5_gen twiddle_rsc_0_3_i
      (
      .q(twiddle_rsc_0_3_q),
      .re(twiddle_rsc_0_3_re),
      .radr(twiddle_rsc_0_3_radr),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .re_d(twiddle_rsc_0_3_i_re_d_iff),
      .q_d(twiddle_rsc_0_3_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_re_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_21_64_7_128_128_64_5_gen twiddle_rsc_0_4_i
      (
      .q(twiddle_rsc_0_4_q),
      .re(twiddle_rsc_0_4_re),
      .radr(twiddle_rsc_0_4_radr),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .re_d(twiddle_rsc_0_4_i_re_d_iff),
      .q_d(twiddle_rsc_0_4_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_re_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_22_64_7_128_128_64_5_gen twiddle_rsc_0_5_i
      (
      .q(twiddle_rsc_0_5_q),
      .re(twiddle_rsc_0_5_re),
      .radr(twiddle_rsc_0_5_radr),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .re_d(twiddle_rsc_0_5_i_re_d_iff),
      .q_d(twiddle_rsc_0_5_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_re_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_23_64_7_128_128_64_5_gen twiddle_rsc_0_6_i
      (
      .q(twiddle_rsc_0_6_q),
      .re(twiddle_rsc_0_6_re),
      .radr(twiddle_rsc_0_6_radr),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .re_d(twiddle_rsc_0_6_i_re_d_iff),
      .q_d(twiddle_rsc_0_6_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_re_d_iff)
    );
  DIT_RELOOP_ccs_sample_mem_ccs_ram_sync_1R1W_rport_24_64_7_128_128_64_5_gen twiddle_rsc_0_7_i
      (
      .q(twiddle_rsc_0_7_q),
      .re(twiddle_rsc_0_7_re),
      .radr(twiddle_rsc_0_7_radr),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .re_d(twiddle_rsc_0_7_i_re_d_iff),
      .q_d(twiddle_rsc_0_7_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_re_d_iff)
    );
  DIT_RELOOP_core DIT_RELOOP_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .twiddle_rsc_triosy_0_0_lz(twiddle_rsc_triosy_0_0_lz),
      .twiddle_rsc_triosy_0_1_lz(twiddle_rsc_triosy_0_1_lz),
      .twiddle_rsc_triosy_0_2_lz(twiddle_rsc_triosy_0_2_lz),
      .twiddle_rsc_triosy_0_3_lz(twiddle_rsc_triosy_0_3_lz),
      .twiddle_rsc_triosy_0_4_lz(twiddle_rsc_triosy_0_4_lz),
      .twiddle_rsc_triosy_0_5_lz(twiddle_rsc_triosy_0_5_lz),
      .twiddle_rsc_triosy_0_6_lz(twiddle_rsc_triosy_0_6_lz),
      .twiddle_rsc_triosy_0_7_lz(twiddle_rsc_triosy_0_7_lz),
      .vec_rsc_0_0_i_radr_d(vec_rsc_0_0_i_radr_d),
      .vec_rsc_0_0_i_q_d(vec_rsc_0_0_i_q_d),
      .vec_rsc_0_1_i_radr_d(vec_rsc_0_1_i_radr_d),
      .vec_rsc_0_1_i_q_d(vec_rsc_0_1_i_q_d),
      .vec_rsc_0_2_i_radr_d(vec_rsc_0_2_i_radr_d),
      .vec_rsc_0_2_i_q_d(vec_rsc_0_2_i_q_d),
      .vec_rsc_0_3_i_radr_d(vec_rsc_0_3_i_radr_d),
      .vec_rsc_0_3_i_q_d(vec_rsc_0_3_i_q_d),
      .vec_rsc_0_4_i_radr_d(vec_rsc_0_4_i_radr_d),
      .vec_rsc_0_4_i_q_d(vec_rsc_0_4_i_q_d),
      .vec_rsc_0_5_i_radr_d(vec_rsc_0_5_i_radr_d),
      .vec_rsc_0_5_i_q_d(vec_rsc_0_5_i_q_d),
      .vec_rsc_0_6_i_radr_d(vec_rsc_0_6_i_radr_d),
      .vec_rsc_0_6_i_q_d(vec_rsc_0_6_i_q_d),
      .vec_rsc_0_7_i_radr_d(vec_rsc_0_7_i_radr_d),
      .vec_rsc_0_7_i_q_d(vec_rsc_0_7_i_q_d),
      .twiddle_rsc_0_0_i_q_d(twiddle_rsc_0_0_i_q_d),
      .twiddle_rsc_0_1_i_q_d(twiddle_rsc_0_1_i_q_d),
      .twiddle_rsc_0_2_i_q_d(twiddle_rsc_0_2_i_q_d),
      .twiddle_rsc_0_3_i_q_d(twiddle_rsc_0_3_i_q_d),
      .twiddle_rsc_0_4_i_q_d(twiddle_rsc_0_4_i_q_d),
      .twiddle_rsc_0_5_i_q_d(twiddle_rsc_0_5_i_q_d),
      .twiddle_rsc_0_6_i_q_d(twiddle_rsc_0_6_i_q_d),
      .twiddle_rsc_0_7_i_q_d(twiddle_rsc_0_7_i_q_d),
      .vec_rsc_0_0_i_wadr_d_pff(vec_rsc_0_0_i_wadr_d_iff),
      .vec_rsc_0_0_i_d_d_pff(vec_rsc_0_0_i_d_d_iff),
      .vec_rsc_0_0_i_we_d_pff(vec_rsc_0_0_i_we_d_iff),
      .vec_rsc_0_0_i_re_d_pff(vec_rsc_0_0_i_re_d_iff),
      .vec_rsc_0_1_i_wadr_d_pff(vec_rsc_0_1_i_wadr_d_iff),
      .vec_rsc_0_1_i_d_d_pff(vec_rsc_0_1_i_d_d_iff),
      .vec_rsc_0_1_i_we_d_pff(vec_rsc_0_1_i_we_d_iff),
      .vec_rsc_0_1_i_re_d_pff(vec_rsc_0_1_i_re_d_iff),
      .vec_rsc_0_2_i_we_d_pff(vec_rsc_0_2_i_we_d_iff),
      .vec_rsc_0_2_i_re_d_pff(vec_rsc_0_2_i_re_d_iff),
      .vec_rsc_0_3_i_we_d_pff(vec_rsc_0_3_i_we_d_iff),
      .vec_rsc_0_3_i_re_d_pff(vec_rsc_0_3_i_re_d_iff),
      .vec_rsc_0_4_i_we_d_pff(vec_rsc_0_4_i_we_d_iff),
      .vec_rsc_0_4_i_re_d_pff(vec_rsc_0_4_i_re_d_iff),
      .vec_rsc_0_5_i_we_d_pff(vec_rsc_0_5_i_we_d_iff),
      .vec_rsc_0_5_i_re_d_pff(vec_rsc_0_5_i_re_d_iff),
      .vec_rsc_0_6_i_we_d_pff(vec_rsc_0_6_i_we_d_iff),
      .vec_rsc_0_6_i_re_d_pff(vec_rsc_0_6_i_re_d_iff),
      .vec_rsc_0_7_i_we_d_pff(vec_rsc_0_7_i_we_d_iff),
      .vec_rsc_0_7_i_re_d_pff(vec_rsc_0_7_i_re_d_iff),
      .twiddle_rsc_0_0_i_radr_d_pff(twiddle_rsc_0_0_i_radr_d_iff),
      .twiddle_rsc_0_0_i_re_d_pff(twiddle_rsc_0_0_i_re_d_iff),
      .twiddle_rsc_0_1_i_re_d_pff(twiddle_rsc_0_1_i_re_d_iff),
      .twiddle_rsc_0_2_i_re_d_pff(twiddle_rsc_0_2_i_re_d_iff),
      .twiddle_rsc_0_3_i_re_d_pff(twiddle_rsc_0_3_i_re_d_iff),
      .twiddle_rsc_0_4_i_re_d_pff(twiddle_rsc_0_4_i_re_d_iff),
      .twiddle_rsc_0_5_i_re_d_pff(twiddle_rsc_0_5_i_re_d_iff),
      .twiddle_rsc_0_6_i_re_d_pff(twiddle_rsc_0_6_i_re_d_iff),
      .twiddle_rsc_0_7_i_re_d_pff(twiddle_rsc_0_7_i_re_d_iff)
    );
endmodule



