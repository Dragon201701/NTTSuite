
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v5.v 
module mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   ls5382@newnano.poly.edu
//  Generated date: Thu Sep 16 11:26:42 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_7_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_7_14_32_16384_16384_32_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output we;
  output [31:0] d;
  output [13:0] wadr;
  input [31:0] d_d;
  output [31:0] q_d;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_5_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_5_14_32_16384_16384_32_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output [31:0] q_d;
  input [13:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_4_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_4_14_32_16384_16384_32_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output [31:0] q_d;
  input [13:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_1_14_32_16384_16384_32_1_gen
// ------------------------------------------------------------------


module ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_1_14_32_16384_16384_32_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [13:0] radr;
  output [31:0] q_d;
  input [13:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module ntt_flat_core_core_fsm (
  clk, rst, fsm_output, for_C_0_tr0, INNER_LOOP_C_2_tr0, STAGE_LOOP_C_1_tr0
);
  input clk;
  input rst;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;
  input for_C_0_tr0;
  input INNER_LOOP_C_2_tr0;
  input STAGE_LOOP_C_1_tr0;


  // FSM State Type Declaration for ntt_flat_core_core_fsm_1
  parameter
    main_C_0 = 3'd0,
    for_C_0 = 3'd1,
    STAGE_LOOP_C_0 = 3'd2,
    INNER_LOOP_C_0 = 3'd3,
    INNER_LOOP_C_1 = 3'd4,
    INNER_LOOP_C_2 = 3'd5,
    STAGE_LOOP_C_1 = 3'd6,
    main_C_1 = 3'd7;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ntt_flat_core_core_fsm_1
    case (state_var)
      for_C_0 : begin
        fsm_output = 8'b00000010;
        if ( for_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      STAGE_LOOP_C_0 : begin
        fsm_output = 8'b00000100;
        state_var_NS = INNER_LOOP_C_0;
      end
      INNER_LOOP_C_0 : begin
        fsm_output = 8'b00001000;
        state_var_NS = INNER_LOOP_C_1;
      end
      INNER_LOOP_C_1 : begin
        fsm_output = 8'b00010000;
        state_var_NS = INNER_LOOP_C_2;
      end
      INNER_LOOP_C_2 : begin
        fsm_output = 8'b00100000;
        if ( INNER_LOOP_C_2_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_1;
        end
        else begin
          state_var_NS = INNER_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 8'b01000000;
        if ( STAGE_LOOP_C_1_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 8'b10000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 8'b00000001;
        state_var_NS = for_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_core_wait_dp
// ------------------------------------------------------------------


module ntt_flat_core_wait_dp (
  clk, mult_t_mul_cmp_z, mult_t_mul_cmp_z_oreg
);
  input clk;
  input [51:0] mult_t_mul_cmp_z;
  output [31:0] mult_t_mul_cmp_z_oreg;


  // Interconnect Declarations
  reg [31:0] mult_t_mul_cmp_z_oreg_pconst_51_20;


  // Interconnect Declarations for Component Instantiations 
  assign mult_t_mul_cmp_z_oreg = mult_t_mul_cmp_z_oreg_pconst_51_20;
  always @(posedge clk) begin
    mult_t_mul_cmp_z_oreg_pconst_51_20 <= mult_t_mul_cmp_z[51:20];
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat_core
// ------------------------------------------------------------------


module ntt_flat_core (
  clk, rst, vec_rsc_triosy_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_triosy_lz, twiddle_rsc_triosy_lz,
      twiddle_h_rsc_triosy_lz, result_rsc_triosy_0_0_lz, result_rsc_triosy_1_0_lz,
      result_rsc_triosy_2_0_lz, result_rsc_triosy_3_0_lz, result_rsc_triosy_4_0_lz,
      result_rsc_triosy_5_0_lz, result_rsc_triosy_6_0_lz, result_rsc_triosy_7_0_lz,
      result_rsc_triosy_8_0_lz, result_rsc_triosy_9_0_lz, result_rsc_triosy_10_0_lz,
      result_rsc_triosy_11_0_lz, result_rsc_triosy_12_0_lz, result_rsc_triosy_13_0_lz,
      result_rsc_triosy_14_0_lz, vec_rsci_q_d, vec_rsci_radr_d, vec_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsci_q_d, twiddle_h_rsci_q_d, result_rsc_0_0_i_d_d, result_rsc_0_0_i_q_d,
      result_rsc_0_0_i_wadr_d, result_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      result_rsc_1_0_i_q_d, result_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d, result_rsc_2_0_i_q_d,
      result_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d, result_rsc_3_0_i_q_d, result_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      result_rsc_4_0_i_q_d, result_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d, result_rsc_5_0_i_q_d,
      result_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d, result_rsc_6_0_i_q_d, result_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      result_rsc_7_0_i_q_d, result_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d, result_rsc_8_0_i_q_d,
      result_rsc_8_0_i_readA_r_ram_ir_internal_RMASK_B_d, result_rsc_9_0_i_q_d, result_rsc_9_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      result_rsc_10_0_i_q_d, result_rsc_10_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      result_rsc_11_0_i_q_d, result_rsc_11_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      result_rsc_12_0_i_q_d, result_rsc_12_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      result_rsc_13_0_i_q_d, result_rsc_13_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      result_rsc_14_0_i_q_d, result_rsc_14_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      mult_t_mul_cmp_a, mult_t_mul_cmp_b, mult_t_mul_cmp_z, twiddle_rsci_radr_d_pff,
      twiddle_rsci_readA_r_ram_ir_internal_RMASK_B_d_pff, result_rsc_0_0_i_radr_d_pff,
      result_rsc_0_0_i_we_d_pff, result_rsc_1_0_i_d_d_pff, result_rsc_1_0_i_we_d_pff,
      result_rsc_2_0_i_we_d_pff, result_rsc_3_0_i_we_d_pff, result_rsc_4_0_i_we_d_pff,
      result_rsc_5_0_i_we_d_pff, result_rsc_6_0_i_we_d_pff, result_rsc_7_0_i_we_d_pff,
      result_rsc_8_0_i_we_d_pff, result_rsc_9_0_i_we_d_pff, result_rsc_10_0_i_we_d_pff,
      result_rsc_11_0_i_we_d_pff, result_rsc_12_0_i_we_d_pff, result_rsc_13_0_i_we_d_pff,
      result_rsc_14_0_i_we_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_lz;
  input [31:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  output r_rsc_triosy_lz;
  output twiddle_rsc_triosy_lz;
  output twiddle_h_rsc_triosy_lz;
  output result_rsc_triosy_0_0_lz;
  output result_rsc_triosy_1_0_lz;
  output result_rsc_triosy_2_0_lz;
  output result_rsc_triosy_3_0_lz;
  output result_rsc_triosy_4_0_lz;
  output result_rsc_triosy_5_0_lz;
  output result_rsc_triosy_6_0_lz;
  output result_rsc_triosy_7_0_lz;
  output result_rsc_triosy_8_0_lz;
  output result_rsc_triosy_9_0_lz;
  output result_rsc_triosy_10_0_lz;
  output result_rsc_triosy_11_0_lz;
  output result_rsc_triosy_12_0_lz;
  output result_rsc_triosy_13_0_lz;
  output result_rsc_triosy_14_0_lz;
  input [31:0] vec_rsci_q_d;
  output [13:0] vec_rsci_radr_d;
  output vec_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] twiddle_rsci_q_d;
  input [31:0] twiddle_h_rsci_q_d;
  output [31:0] result_rsc_0_0_i_d_d;
  input [31:0] result_rsc_0_0_i_q_d;
  output [13:0] result_rsc_0_0_i_wadr_d;
  output result_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_1_0_i_q_d;
  output result_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_2_0_i_q_d;
  output result_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_3_0_i_q_d;
  output result_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_4_0_i_q_d;
  output result_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_5_0_i_q_d;
  output result_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_6_0_i_q_d;
  output result_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_7_0_i_q_d;
  output result_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_8_0_i_q_d;
  output result_rsc_8_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_9_0_i_q_d;
  output result_rsc_9_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_10_0_i_q_d;
  output result_rsc_10_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_11_0_i_q_d;
  output result_rsc_11_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_12_0_i_q_d;
  output result_rsc_12_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_13_0_i_q_d;
  output result_rsc_13_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] result_rsc_14_0_i_q_d;
  output result_rsc_14_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  output [31:0] mult_t_mul_cmp_a;
  reg [31:0] mult_t_mul_cmp_a;
  output [31:0] mult_t_mul_cmp_b;
  reg [31:0] mult_t_mul_cmp_b;
  input [51:0] mult_t_mul_cmp_z;
  output [13:0] twiddle_rsci_radr_d_pff;
  wire [28:0] nl_twiddle_rsci_radr_d_pff;
  output twiddle_rsci_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output [13:0] result_rsc_0_0_i_radr_d_pff;
  output result_rsc_0_0_i_we_d_pff;
  output [31:0] result_rsc_1_0_i_d_d_pff;
  output result_rsc_1_0_i_we_d_pff;
  output result_rsc_2_0_i_we_d_pff;
  output result_rsc_3_0_i_we_d_pff;
  output result_rsc_4_0_i_we_d_pff;
  output result_rsc_5_0_i_we_d_pff;
  output result_rsc_6_0_i_we_d_pff;
  output result_rsc_7_0_i_we_d_pff;
  output result_rsc_8_0_i_we_d_pff;
  output result_rsc_9_0_i_we_d_pff;
  output result_rsc_10_0_i_we_d_pff;
  output result_rsc_11_0_i_we_d_pff;
  output result_rsc_12_0_i_we_d_pff;
  output result_rsc_13_0_i_we_d_pff;
  output result_rsc_14_0_i_we_d_pff;


  // Interconnect Declarations
  wire [31:0] p_rsci_idat;
  wire [31:0] mult_t_mul_cmp_z_oreg;
  wire [7:0] fsm_output;
  wire [3:0] butterFly_f2_acc_1_tmp;
  wire [4:0] nl_butterFly_f2_acc_1_tmp;
  wire [3:0] butterFly_f1_acc_1_tmp;
  wire [4:0] nl_butterFly_f1_acc_1_tmp;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire and_dcpl_17;
  wire and_dcpl_19;
  wire and_dcpl_20;
  wire and_dcpl_21;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_25;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_31;
  wire and_dcpl_33;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_40;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire and_dcpl_45;
  wire and_dcpl_47;
  wire and_dcpl_50;
  wire and_dcpl_52;
  wire and_dcpl_54;
  wire and_dcpl_56;
  wire and_dcpl_58;
  wire and_dcpl_60;
  wire and_dcpl_62;
  wire and_dcpl_68;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_80;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_87;
  wire and_dcpl_101;
  wire and_dcpl_103;
  wire and_dcpl_105;
  wire or_dcpl_29;
  wire or_dcpl_30;
  wire [13:0] INNER_LOOP_j_13_0_sva_2;
  wire [14:0] nl_INNER_LOOP_j_13_0_sva_2;
  reg [3:0] butterFly_acc_4_itm_3;
  reg INNER_LOOP_stage_0;
  reg INNER_LOOP_stage_0_1;
  reg [3:0] butterFly_acc_4_itm_2;
  reg INNER_LOOP_stage_0_3;
  reg [3:0] butterFly_acc_itm_1;
  wire [4:0] nl_butterFly_acc_itm_1;
  reg [3:0] butterFly_acc_itm_2;
  reg [3:0] butterFly_acc_4_itm_1;
  wire [4:0] nl_butterFly_acc_4_itm_1;
  reg INNER_LOOP_stage_0_2;
  reg [31:0] p_sva;
  wire [31:0] modulo_add_base_sva_1;
  wire [32:0] nl_modulo_add_base_sva_1;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  wire [17:0] butterFly_idx2_17_0_sva_1;
  wire [18:0] nl_butterFly_idx2_17_0_sva_1;
  reg reg_vec_rsc_triosy_obj_ld_cse;
  wire INNER_LOOP_or_1_cse;
  wire nor_6_cse;
  wire butterFly_f2_nor_9_cse;
  reg [13:0] operator_33_true_return_13_0_sva;
  reg [17:0] INNER_LOOP_k_17_0_sva;
  wire [18:0] nl_INNER_LOOP_k_17_0_sva;
  reg [31:0] mult_res_lpi_3_dfm;
  reg [12:0] INNER_LOOP_idx1_acc_psp_sva_1_12_0;
  reg INNER_LOOP_k_17_0_sva_1_0;
  reg [13:0] butterFly_idx2_17_0_sva_3_13_0;
  wire [31:0] z_out;
  wire [31:0] z_out_1;
  wire [31:0] z_out_2;
  wire [31:0] z_out_3;
  wire [63:0] nl_z_out_3;
  wire [17:0] z_out_4;
  wire [13:0] z_out_5;
  wire [14:0] z_out_6;
  wire [15:0] nl_z_out_6;
  reg [3:0] operator_20_false_acc_psp_sva;
  wire [4:0] nl_operator_20_false_acc_psp_sva;
  reg [13:0] operator_20_false_rshift_psp_sva;
  reg [12:0] INNER_LOOP_g_rshift_psp_sva;
  reg [31:0] tmp_1_lpi_3_dfm;
  reg INNER_LOOP_stage_0_4;
  reg [16:0] INNER_LOOP_idx1_mul_itm;
  reg [31:0] mult_z_mul_itm;
  wire [63:0] nl_mult_z_mul_itm;
  reg [31:0] operator_96_false_operator_96_false_slc_mult_t_mul_51_20_itm;
  reg [3:0] butterFly_f2_acc_1_svs_1;
  reg [31:0] modulo_add_qr_lpi_3_dfm_1;
  reg butterFly_f1_butterFly_f1_nor_itm_1;
  reg butterFly_f1_nor_itm_1;
  reg butterFly_f1_nor_1_itm_1;
  reg butterFly_f1_butterFly_f1_and_2_itm_1;
  reg butterFly_f1_nor_3_itm_1;
  reg butterFly_f1_butterFly_f1_and_4_itm_1;
  reg butterFly_f1_butterFly_f1_and_5_itm_1;
  reg butterFly_f1_butterFly_f1_and_6_itm_1;
  reg butterFly_f1_nor_6_itm_1;
  reg butterFly_f1_butterFly_f1_and_8_itm_1;
  reg butterFly_f1_butterFly_f1_and_9_itm_1;
  reg butterFly_f1_butterFly_f1_and_10_itm_1;
  reg butterFly_f1_butterFly_f1_and_11_itm_1;
  reg butterFly_f1_butterFly_f1_and_12_itm_1;
  reg butterFly_f1_butterFly_f1_and_13_itm_1;
  reg butterFly_f2_butterFly_f2_nor_itm_1;
  reg butterFly_f2_nor_itm_1;
  reg butterFly_f2_nor_1_itm_1;
  reg butterFly_f2_butterFly_f2_and_2_itm_1;
  reg butterFly_f2_nor_3_itm_1;
  reg butterFly_f2_butterFly_f2_and_4_itm_1;
  reg butterFly_f2_butterFly_f2_and_5_itm_1;
  reg butterFly_f2_butterFly_f2_and_6_itm_1;
  reg butterFly_f2_nor_6_itm_1;
  reg butterFly_f2_butterFly_f2_and_8_itm_1;
  reg butterFly_f2_butterFly_f2_and_9_itm_1;
  reg butterFly_f2_butterFly_f2_and_10_itm_1;
  reg butterFly_f2_butterFly_f2_and_11_itm_1;
  reg butterFly_f2_butterFly_f2_and_12_itm_1;
  reg butterFly_f2_butterFly_f2_and_13_itm_1;
  reg [31:0] INNER_LOOP_tf_asn_itm_1;
  reg [31:0] INNER_LOOP_tf_asn_itm_2;
  reg [31:0] mult_z_mul_itm_1;
  reg [31:0] INNER_LOOP_tf_h_asn_itm_1;
  reg [31:0] mult_z_mul_itm_1_1;
  reg [12:0] INNER_LOOP_j_13_0_sva_12_0;
  reg INNER_LOOP_k_17_0_sva_2_0;
  reg [12:0] INNER_LOOP_idx1_acc_psp_sva_2_12_0;
  reg [13:0] butterFly_idx2_17_0_sva_1_13_0;
  reg [13:0] butterFly_idx2_17_0_sva_2_13_0;
  wire [16:0] INNER_LOOP_idx1_acc_psp_sva_1;
  wire [17:0] nl_INNER_LOOP_idx1_acc_psp_sva_1;
  reg [3:0] reg_butterFly_f1_acc_1_svs_st_1_cse;
  wire INNER_LOOP_j_or_cse;
  wire operator_20_false_acc_itm_4_1;
  wire z_out_7_32;

  wire[0:0] butterFly_mux_nl;
  wire[0:0] INNER_LOOP_INNER_LOOP_and_nl;
  wire[0:0] or_101_nl;
  wire[13:0] for_i_for_i_mux_nl;
  wire[0:0] INNER_LOOP_nor_nl;
  wire[31:0] modulo_add_qif_acc_nl;
  wire[32:0] nl_modulo_add_qif_acc_nl;
  wire[0:0] for_and_1_nl;
  wire[4:0] operator_20_false_acc_nl;
  wire[5:0] nl_operator_20_false_acc_nl;
  wire[32:0] acc_nl;
  wire[33:0] nl_acc_nl;
  wire[0:0] modulo_sub_qif_modulo_sub_qif_or_1_nl;
  wire[0:0] modulo_sub_qif_or_1_nl;
  wire[31:0] modulo_sub_qif_mux_2_nl;
  wire[32:0] acc_1_nl;
  wire[33:0] nl_acc_1_nl;
  wire[31:0] mult_res_mux_3_nl;
  wire[31:0] mult_z_mux_2_nl;
  wire[31:0] mult_z_mux_3_nl;
  wire[13:0] STAGE_LOOP_mux_1_nl;
  wire[33:0] acc_3_nl;
  wire[34:0] nl_acc_3_nl;
  wire[31:0] modulo_add_mux_3_nl;
  wire[31:0] modulo_add_mux_4_nl;
  wire[0:0] butterFly_f1_mux_32_nl;
  wire[0:0] butterFly_f1_mux_33_nl;
  wire[0:0] butterFly_f1_butterFly_f1_and_14_nl;
  wire[0:0] butterFly_f2_butterFly_f2_and_14_nl;
  wire[0:0] butterFly_f1_mux_34_nl;
  wire[0:0] butterFly_f1_butterFly_f1_and_15_nl;
  wire[0:0] butterFly_f2_butterFly_f2_and_15_nl;
  wire[0:0] butterFly_f1_mux_35_nl;
  wire[0:0] butterFly_f1_mux_36_nl;
  wire[0:0] butterFly_f1_butterFly_f1_and_16_nl;
  wire[0:0] butterFly_f2_butterFly_f2_and_16_nl;
  wire[0:0] butterFly_f1_mux_37_nl;
  wire[0:0] butterFly_f1_mux_38_nl;
  wire[0:0] butterFly_f1_mux_39_nl;
  wire[0:0] butterFly_f1_mux_40_nl;
  wire[0:0] butterFly_f1_butterFly_f1_and_17_nl;
  wire[0:0] butterFly_f2_butterFly_f2_and_17_nl;
  wire[0:0] butterFly_f1_mux_41_nl;
  wire[0:0] butterFly_f1_mux_42_nl;
  wire[0:0] butterFly_f1_mux_43_nl;
  wire[0:0] butterFly_f1_mux_44_nl;
  wire[0:0] butterFly_f1_mux_45_nl;
  wire[0:0] butterFly_f1_mux_46_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [12:0] nl_INNER_LOOP_k_lshift_rg_a;
  assign nl_INNER_LOOP_k_lshift_rg_a = MUX_v_13_2_2(13'b0000000000001, (z_out_5[12:0]),
      fsm_output[3]);
  wire[3:0] operator_20_false_1_acc_nl;
  wire[4:0] nl_operator_20_false_1_acc_nl;
  wire [3:0] nl_INNER_LOOP_k_lshift_rg_s;
  assign nl_operator_20_false_1_acc_nl = STAGE_LOOP_i_3_0_sva + 4'b1111;
  assign operator_20_false_1_acc_nl = nl_operator_20_false_1_acc_nl[3:0];
  assign nl_INNER_LOOP_k_lshift_rg_s = MUX_v_4_2_2(operator_20_false_1_acc_nl, operator_20_false_acc_psp_sva,
      fsm_output[3]);
  wire[12:0] operator_20_false_operator_20_false_and_nl;
  wire [14:0] nl_INNER_LOOP_g_rshift_rg_a;
  assign operator_20_false_operator_20_false_and_nl = MUX_v_13_2_2(13'b0000000000000,
      INNER_LOOP_j_13_0_sva_12_0, (fsm_output[3]));
  assign nl_INNER_LOOP_g_rshift_rg_a = {(~ (fsm_output[3])) , 1'b0 , operator_20_false_operator_20_false_and_nl};
  wire [3:0] nl_INNER_LOOP_g_rshift_rg_s;
  assign nl_INNER_LOOP_g_rshift_rg_s = MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, operator_20_false_acc_psp_sva,
      fsm_output[3]);
  wire [0:0] nl_ntt_flat_core_core_fsm_inst_INNER_LOOP_C_2_tr0;
  assign nl_ntt_flat_core_core_fsm_inst_INNER_LOOP_C_2_tr0 = (~(INNER_LOOP_stage_0_2
      | INNER_LOOP_stage_0_3)) & nor_6_cse;
  wire [0:0] nl_ntt_flat_core_core_fsm_inst_STAGE_LOOP_C_1_tr0;
  assign nl_ntt_flat_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 = operator_20_false_acc_itm_4_1;
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd32)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(vec_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(twiddle_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_14_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_14_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_13_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_13_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_12_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_12_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_11_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_11_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_10_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_10_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_9_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_9_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_8_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_8_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_7_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_7_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_6_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_6_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_5_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_5_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_4_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_4_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_3_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_3_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_2_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_2_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_1_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_1_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_obj_ld_cse),
      .lz(result_rsc_triosy_0_0_lz)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd18)) INNER_LOOP_k_lshift_rg (
      .a(nl_INNER_LOOP_k_lshift_rg_a[12:0]),
      .s(nl_INNER_LOOP_k_lshift_rg_s[3:0]),
      .z(z_out_4)
    );
  mgc_shift_r_v5 #(.width_a(32'sd15),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd14)) INNER_LOOP_g_rshift_rg (
      .a(nl_INNER_LOOP_g_rshift_rg_a[14:0]),
      .s(nl_INNER_LOOP_g_rshift_rg_s[3:0]),
      .z(z_out_5)
    );
  ntt_flat_core_wait_dp ntt_flat_core_wait_dp_inst (
      .clk(clk),
      .mult_t_mul_cmp_z(mult_t_mul_cmp_z),
      .mult_t_mul_cmp_z_oreg(mult_t_mul_cmp_z_oreg)
    );
  ntt_flat_core_core_fsm ntt_flat_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .for_C_0_tr0(nor_6_cse),
      .INNER_LOOP_C_2_tr0(nl_ntt_flat_core_core_fsm_inst_INNER_LOOP_C_2_tr0[0:0]),
      .STAGE_LOOP_C_1_tr0(nl_ntt_flat_core_core_fsm_inst_STAGE_LOOP_C_1_tr0[0:0])
    );
  assign nor_6_cse = ~(INNER_LOOP_stage_0_1 | INNER_LOOP_stage_0);
  assign butterFly_f2_nor_9_cse = ~((butterFly_f2_acc_1_tmp[1:0]!=2'b00));
  assign INNER_LOOP_j_or_cse = (fsm_output[5:3]!=3'b000);
  assign INNER_LOOP_or_1_cse = (fsm_output[2]) | (fsm_output[5]);
  assign nl_butterFly_f2_acc_1_tmp = (butterFly_idx2_17_0_sva_1[17:14]) + STAGE_LOOP_i_3_0_sva;
  assign butterFly_f2_acc_1_tmp = nl_butterFly_f2_acc_1_tmp[3:0];
  assign nl_butterFly_f1_acc_1_tmp = (INNER_LOOP_idx1_acc_psp_sva_1[16:13]) + STAGE_LOOP_i_3_0_sva;
  assign butterFly_f1_acc_1_tmp = nl_butterFly_f1_acc_1_tmp[3:0];
  assign nl_INNER_LOOP_j_13_0_sva_2 = conv_u2u_13_14(INNER_LOOP_j_13_0_sva_12_0)
      + 14'b00000000000001;
  assign INNER_LOOP_j_13_0_sva_2 = nl_INNER_LOOP_j_13_0_sva_2[13:0];
  assign nl_modulo_add_base_sva_1 = mult_z_mul_itm_1 + tmp_1_lpi_3_dfm;
  assign modulo_add_base_sva_1 = nl_modulo_add_base_sva_1[31:0];
  assign nl_butterFly_idx2_17_0_sva_1 = ({INNER_LOOP_idx1_acc_psp_sva_1 , (INNER_LOOP_k_17_0_sva[0])})
      + conv_u2u_14_18(operator_20_false_rshift_psp_sva);
  assign butterFly_idx2_17_0_sva_1 = nl_butterFly_idx2_17_0_sva_1[17:0];
  assign nl_INNER_LOOP_idx1_acc_psp_sva_1 = INNER_LOOP_idx1_mul_itm + (INNER_LOOP_k_17_0_sva[17:1]);
  assign INNER_LOOP_idx1_acc_psp_sva_1 = nl_INNER_LOOP_idx1_acc_psp_sva_1[16:0];
  assign nl_operator_20_false_acc_nl = ({1'b1 , (~ (z_out_6[3:0]))}) + 5'b01111;
  assign operator_20_false_acc_nl = nl_operator_20_false_acc_nl[4:0];
  assign operator_20_false_acc_itm_4_1 = readslicef_5_1_4(operator_20_false_acc_nl);
  assign and_dcpl_15 = ~((butterFly_acc_itm_2[2:1]!=2'b00));
  assign and_dcpl_16 = INNER_LOOP_stage_0_3 & (~ (butterFly_acc_itm_2[3]));
  assign and_dcpl_17 = and_dcpl_16 & (~ (butterFly_acc_itm_2[0]));
  assign and_dcpl_19 = ~((butterFly_acc_4_itm_3[3:2]!=2'b00));
  assign and_dcpl_20 = (~ (butterFly_acc_4_itm_3[1])) & INNER_LOOP_stage_0_4;
  assign and_dcpl_21 = and_dcpl_20 & (~ (butterFly_acc_4_itm_3[0]));
  assign and_dcpl_23 = ~((reg_butterFly_f1_acc_1_svs_st_1_cse[3:2]!=2'b00));
  assign and_dcpl_24 = INNER_LOOP_stage_0_2 & (~ (reg_butterFly_f1_acc_1_svs_st_1_cse[0]));
  assign and_dcpl_25 = and_dcpl_24 & (~ (reg_butterFly_f1_acc_1_svs_st_1_cse[1]));
  assign and_dcpl_28 = INNER_LOOP_stage_0_1 & (~ (butterFly_f2_acc_1_tmp[3]));
  assign and_dcpl_29 = and_dcpl_28 & (~ (butterFly_f2_acc_1_tmp[2]));
  assign and_dcpl_31 = and_dcpl_16 & (butterFly_acc_itm_2[0]);
  assign and_dcpl_33 = and_dcpl_20 & (butterFly_acc_4_itm_3[0]);
  assign and_dcpl_35 = INNER_LOOP_stage_0_2 & (reg_butterFly_f1_acc_1_svs_st_1_cse[0]);
  assign and_dcpl_36 = and_dcpl_35 & (~ (reg_butterFly_f1_acc_1_svs_st_1_cse[1]));
  assign and_dcpl_38 = (butterFly_f2_acc_1_tmp[1:0]==2'b01);
  assign and_dcpl_40 = (butterFly_acc_itm_2[2:1]==2'b01);
  assign and_dcpl_42 = (butterFly_acc_4_itm_3[1]) & INNER_LOOP_stage_0_4;
  assign and_dcpl_43 = and_dcpl_42 & (~ (butterFly_acc_4_itm_3[0]));
  assign and_dcpl_45 = and_dcpl_24 & (reg_butterFly_f1_acc_1_svs_st_1_cse[1]);
  assign and_dcpl_47 = (butterFly_f2_acc_1_tmp[1:0]==2'b10);
  assign and_dcpl_50 = and_dcpl_42 & (butterFly_acc_4_itm_3[0]);
  assign and_dcpl_52 = and_dcpl_35 & (reg_butterFly_f1_acc_1_svs_st_1_cse[1]);
  assign and_dcpl_54 = (butterFly_f2_acc_1_tmp[1:0]==2'b11);
  assign and_dcpl_56 = (butterFly_acc_itm_2[2:1]==2'b10);
  assign and_dcpl_58 = (butterFly_acc_4_itm_3[3:2]==2'b01);
  assign and_dcpl_60 = (reg_butterFly_f1_acc_1_svs_st_1_cse[3:2]==2'b01);
  assign and_dcpl_62 = and_dcpl_28 & (butterFly_f2_acc_1_tmp[2]);
  assign and_dcpl_68 = (butterFly_acc_itm_2[2:1]==2'b11);
  assign and_dcpl_77 = INNER_LOOP_stage_0_3 & (butterFly_acc_itm_2[3]);
  assign and_dcpl_78 = and_dcpl_77 & (~ (butterFly_acc_itm_2[0]));
  assign and_dcpl_80 = (butterFly_acc_4_itm_3[3:2]==2'b10);
  assign and_dcpl_82 = (reg_butterFly_f1_acc_1_svs_st_1_cse[3:2]==2'b10);
  assign and_dcpl_84 = INNER_LOOP_stage_0_1 & (butterFly_f2_acc_1_tmp[3]);
  assign and_dcpl_85 = and_dcpl_84 & (~ (butterFly_f2_acc_1_tmp[2]));
  assign and_dcpl_87 = and_dcpl_77 & (butterFly_acc_itm_2[0]);
  assign and_dcpl_101 = (butterFly_acc_4_itm_3[3:2]==2'b11);
  assign and_dcpl_103 = (reg_butterFly_f1_acc_1_svs_st_1_cse[3:2]==2'b11);
  assign and_dcpl_105 = and_dcpl_84 & (butterFly_f2_acc_1_tmp[2]);
  assign or_dcpl_29 = (fsm_output[0]) | (fsm_output[2]);
  assign or_dcpl_30 = (fsm_output[7:6]!=2'b00);
  assign vec_rsci_radr_d = butterFly_idx2_17_0_sva_2_13_0;
  assign vec_rsci_readA_r_ram_ir_internal_RMASK_B_d = INNER_LOOP_stage_0 & (fsm_output[1]);
  assign nl_twiddle_rsci_radr_d_pff = $signed(operator_33_true_return_13_0_sva) *
      $signed(conv_u2s_14_15(INNER_LOOP_k_17_0_sva[13:0]));
  assign twiddle_rsci_radr_d_pff = nl_twiddle_rsci_radr_d_pff[13:0];
  assign twiddle_rsci_readA_r_ram_ir_internal_RMASK_B_d_pff = INNER_LOOP_stage_0_1
      & (fsm_output[4]);
  assign result_rsc_0_0_i_d_d = MUX1HOT_v_32_3_2(vec_rsci_q_d, mult_res_lpi_3_dfm,
      modulo_add_qr_lpi_3_dfm_1, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign result_rsc_0_0_i_radr_d_pff = MUX_v_14_2_2(({INNER_LOOP_idx1_acc_psp_sva_1_12_0
      , INNER_LOOP_k_17_0_sva_1_0}), (butterFly_idx2_17_0_sva_1[13:0]), fsm_output[5]);
  assign result_rsc_0_0_i_wadr_d = MUX_v_14_2_2(butterFly_idx2_17_0_sva_3_13_0, ({INNER_LOOP_idx1_acc_psp_sva_2_12_0
      , INNER_LOOP_k_17_0_sva_2_0}), fsm_output[5]);
  assign result_rsc_0_0_i_we_d_pff = (and_dcpl_17 & and_dcpl_15 & (fsm_output[5]))
      | (INNER_LOOP_stage_0_1 & (fsm_output[1])) | (and_dcpl_21 & and_dcpl_19 & (fsm_output[4]));
  assign result_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_25 & and_dcpl_23
      & (fsm_output[3])) | (and_dcpl_29 & butterFly_f2_nor_9_cse & (fsm_output[5]));
  assign result_rsc_1_0_i_d_d_pff = MUX_v_32_2_2(mult_res_lpi_3_dfm, modulo_add_qr_lpi_3_dfm_1,
      fsm_output[5]);
  assign result_rsc_1_0_i_we_d_pff = (and_dcpl_31 & and_dcpl_15 & (fsm_output[5]))
      | (and_dcpl_33 & and_dcpl_19 & (fsm_output[4]));
  assign result_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_36 & and_dcpl_23
      & (fsm_output[3])) | (and_dcpl_29 & and_dcpl_38 & (fsm_output[5]));
  assign result_rsc_2_0_i_we_d_pff = (and_dcpl_17 & and_dcpl_40 & (fsm_output[5]))
      | (and_dcpl_43 & and_dcpl_19 & (fsm_output[4]));
  assign result_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_45 & and_dcpl_23
      & (fsm_output[3])) | (and_dcpl_29 & and_dcpl_47 & (fsm_output[5]));
  assign result_rsc_3_0_i_we_d_pff = (and_dcpl_31 & and_dcpl_40 & (fsm_output[5]))
      | (and_dcpl_50 & and_dcpl_19 & (fsm_output[4]));
  assign result_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_52 & and_dcpl_23
      & (fsm_output[3])) | (and_dcpl_29 & and_dcpl_54 & (fsm_output[5]));
  assign result_rsc_4_0_i_we_d_pff = (and_dcpl_17 & and_dcpl_56 & (fsm_output[5]))
      | (and_dcpl_21 & and_dcpl_58 & (fsm_output[4]));
  assign result_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_25 & and_dcpl_60
      & (fsm_output[3])) | (and_dcpl_62 & butterFly_f2_nor_9_cse & (fsm_output[5]));
  assign result_rsc_5_0_i_we_d_pff = (and_dcpl_31 & and_dcpl_56 & (fsm_output[5]))
      | (and_dcpl_33 & and_dcpl_58 & (fsm_output[4]));
  assign result_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_36 & and_dcpl_60
      & (fsm_output[3])) | (and_dcpl_62 & and_dcpl_38 & (fsm_output[5]));
  assign result_rsc_6_0_i_we_d_pff = (and_dcpl_17 & and_dcpl_68 & (fsm_output[5]))
      | (and_dcpl_43 & and_dcpl_58 & (fsm_output[4]));
  assign result_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_45 & and_dcpl_60
      & (fsm_output[3])) | (and_dcpl_62 & and_dcpl_47 & (fsm_output[5]));
  assign result_rsc_7_0_i_we_d_pff = (and_dcpl_31 & and_dcpl_68 & (fsm_output[5]))
      | (and_dcpl_50 & and_dcpl_58 & (fsm_output[4]));
  assign result_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_52 & and_dcpl_60
      & (fsm_output[3])) | (and_dcpl_62 & and_dcpl_54 & (fsm_output[5]));
  assign result_rsc_8_0_i_we_d_pff = (and_dcpl_78 & and_dcpl_15 & (fsm_output[5]))
      | (and_dcpl_21 & and_dcpl_80 & (fsm_output[4]));
  assign result_rsc_8_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_25 & and_dcpl_82
      & (fsm_output[3])) | (and_dcpl_85 & butterFly_f2_nor_9_cse & (fsm_output[5]));
  assign result_rsc_9_0_i_we_d_pff = (and_dcpl_87 & and_dcpl_15 & (fsm_output[5]))
      | (and_dcpl_33 & and_dcpl_80 & (fsm_output[4]));
  assign result_rsc_9_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_36 & and_dcpl_82
      & (fsm_output[3])) | (and_dcpl_85 & and_dcpl_38 & (fsm_output[5]));
  assign result_rsc_10_0_i_we_d_pff = (and_dcpl_78 & and_dcpl_40 & (fsm_output[5]))
      | (and_dcpl_43 & and_dcpl_80 & (fsm_output[4]));
  assign result_rsc_10_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_45 & and_dcpl_82
      & (fsm_output[3])) | (and_dcpl_85 & and_dcpl_47 & (fsm_output[5]));
  assign result_rsc_11_0_i_we_d_pff = (and_dcpl_87 & and_dcpl_40 & (fsm_output[5]))
      | (and_dcpl_50 & and_dcpl_80 & (fsm_output[4]));
  assign result_rsc_11_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_52 & and_dcpl_82
      & (fsm_output[3])) | (and_dcpl_85 & and_dcpl_54 & (fsm_output[5]));
  assign result_rsc_12_0_i_we_d_pff = (and_dcpl_78 & and_dcpl_56 & (fsm_output[5]))
      | (and_dcpl_21 & and_dcpl_101 & (fsm_output[4]));
  assign result_rsc_12_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_25 & and_dcpl_103
      & (fsm_output[3])) | (and_dcpl_105 & butterFly_f2_nor_9_cse & (fsm_output[5]));
  assign result_rsc_13_0_i_we_d_pff = (and_dcpl_87 & and_dcpl_56 & (fsm_output[5]))
      | (and_dcpl_33 & and_dcpl_101 & (fsm_output[4]));
  assign result_rsc_13_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_36 & and_dcpl_103
      & (fsm_output[3])) | (and_dcpl_105 & and_dcpl_38 & (fsm_output[5]));
  assign result_rsc_14_0_i_we_d_pff = (and_dcpl_78 & and_dcpl_68 & (fsm_output[5]))
      | (and_dcpl_43 & and_dcpl_101 & (fsm_output[4]));
  assign result_rsc_14_0_i_readA_r_ram_ir_internal_RMASK_B_d = (and_dcpl_45 & and_dcpl_103
      & (fsm_output[3])) | (and_dcpl_105 & and_dcpl_47 & (fsm_output[5]));
  always @(posedge clk) begin
    if ( (fsm_output[7]) | (fsm_output[0]) ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_obj_ld_cse <= 1'b0;
      INNER_LOOP_stage_0 <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_obj_ld_cse <= operator_20_false_acc_itm_4_1 & (fsm_output[6]);
      INNER_LOOP_stage_0 <= (butterFly_mux_nl & (~(or_dcpl_30 | (INNER_LOOP_stage_0_1
          & (INNER_LOOP_j_13_0_sva_2[13]) & (fsm_output[3]))))) | or_dcpl_29;
    end
  end
  always @(posedge clk) begin
    mult_t_mul_cmp_b <= INNER_LOOP_tf_h_asn_itm_1;
    mult_z_mul_itm_1 <= MUX_v_32_2_2(z_out_2, mult_z_mul_itm, fsm_output[5]);
    INNER_LOOP_tf_asn_itm_2 <= INNER_LOOP_tf_asn_itm_1;
  end
  always @(posedge clk) begin
    if ( INNER_LOOP_stage_0_2 ) begin
      mult_t_mul_cmp_a <= MUX_v_32_2_2(({1'b0 , (z_out_1[30:0])}), z_out, z_out_1[31]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      INNER_LOOP_stage_0_1 <= 1'b0;
    end
    else if ( (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[2])
        ) begin
      INNER_LOOP_stage_0_1 <= (INNER_LOOP_stage_0 & (~ (fsm_output[0]))) | (fsm_output[2]);
    end
  end
  always @(posedge clk) begin
    if ( (fsm_output[5]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[7]) |
        (fsm_output[0]) | (fsm_output[6]) ) begin
      butterFly_idx2_17_0_sva_2_13_0 <= MUX_v_14_2_2(14'b00000000000000, for_i_for_i_mux_nl,
          INNER_LOOP_nor_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ (fsm_output[3]) ) begin
      butterFly_idx2_17_0_sva_3_13_0 <= butterFly_idx2_17_0_sva_2_13_0;
    end
  end
  always @(posedge clk) begin
    if ( (fsm_output[6]) | (fsm_output[1]) ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, (z_out_6[3:0]), fsm_output[6]);
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP_stage_0_3 ) begin
      mult_z_mul_itm_1_1 <= z_out_3;
      operator_96_false_operator_96_false_slc_mult_t_mul_51_20_itm <= mult_t_mul_cmp_z_oreg;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      INNER_LOOP_idx1_acc_psp_sva_1_12_0 <= INNER_LOOP_idx1_acc_psp_sva_1[12:0];
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      INNER_LOOP_k_17_0_sva_1_0 <= INNER_LOOP_k_17_0_sva[0];
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP_stage_0_1 ) begin
      INNER_LOOP_g_rshift_psp_sva <= z_out_5[12:0];
      INNER_LOOP_idx1_mul_itm <= z_out_3[16:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f2_butterFly_f2_nor_itm_1 <= 1'b0;
      butterFly_f2_acc_1_svs_1 <= 4'b0000;
      butterFly_f2_nor_itm_1 <= 1'b0;
      butterFly_f2_nor_1_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_2_itm_1 <= 1'b0;
      butterFly_f2_nor_3_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_4_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_5_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_6_itm_1 <= 1'b0;
      butterFly_f2_nor_6_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_8_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_9_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_10_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_11_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_12_itm_1 <= 1'b0;
      butterFly_f2_butterFly_f2_and_13_itm_1 <= 1'b0;
    end
    else if ( INNER_LOOP_stage_0_1 ) begin
      butterFly_f2_butterFly_f2_nor_itm_1 <= ~((butterFly_f2_acc_1_tmp!=4'b0000));
      butterFly_f2_acc_1_svs_1 <= butterFly_f2_acc_1_tmp;
      butterFly_f2_nor_itm_1 <= ~((butterFly_f2_acc_1_tmp[3:1]!=3'b000));
      butterFly_f2_nor_1_itm_1 <= ~((butterFly_f2_acc_1_tmp[3]) | (butterFly_f2_acc_1_tmp[2])
          | (butterFly_f2_acc_1_tmp[0]));
      butterFly_f2_butterFly_f2_and_2_itm_1 <= (butterFly_f2_acc_1_tmp==4'b0011);
      butterFly_f2_nor_3_itm_1 <= ~((butterFly_f2_acc_1_tmp[3]) | (butterFly_f2_acc_1_tmp[1])
          | (butterFly_f2_acc_1_tmp[0]));
      butterFly_f2_butterFly_f2_and_4_itm_1 <= (butterFly_f2_acc_1_tmp==4'b0101);
      butterFly_f2_butterFly_f2_and_5_itm_1 <= (butterFly_f2_acc_1_tmp==4'b0110);
      butterFly_f2_butterFly_f2_and_6_itm_1 <= (butterFly_f2_acc_1_tmp==4'b0111);
      butterFly_f2_nor_6_itm_1 <= ~((butterFly_f2_acc_1_tmp[2:0]!=3'b000));
      butterFly_f2_butterFly_f2_and_8_itm_1 <= (butterFly_f2_acc_1_tmp==4'b1001);
      butterFly_f2_butterFly_f2_and_9_itm_1 <= (butterFly_f2_acc_1_tmp==4'b1010);
      butterFly_f2_butterFly_f2_and_10_itm_1 <= (butterFly_f2_acc_1_tmp==4'b1011);
      butterFly_f2_butterFly_f2_and_11_itm_1 <= (butterFly_f2_acc_1_tmp[3:2]==2'b11)
          & butterFly_f2_nor_9_cse;
      butterFly_f2_butterFly_f2_and_12_itm_1 <= (butterFly_f2_acc_1_tmp==4'b1101);
      butterFly_f2_butterFly_f2_and_13_itm_1 <= (butterFly_f2_acc_1_tmp==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_butterFly_f1_acc_1_svs_st_1_cse <= 4'b0000;
    end
    else if ( fsm_output[5] ) begin
      reg_butterFly_f1_acc_1_svs_st_1_cse <= butterFly_f1_acc_1_tmp;
    end
  end
  always @(posedge clk) begin
    if ( (INNER_LOOP_stage_0_1 | (~ (fsm_output[3]))) & (fsm_output[5:4]==2'b00)
        ) begin
      INNER_LOOP_j_13_0_sva_12_0 <= MUX_v_13_2_2(13'b0000000000000, (INNER_LOOP_j_13_0_sva_2[12:0]),
          INNER_LOOP_j_or_cse);
    end
  end
  always @(posedge clk) begin
    if ( ~ INNER_LOOP_j_or_cse ) begin
      operator_20_false_acc_psp_sva <= nl_operator_20_false_acc_psp_sva[3:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_acc_4_itm_3 <= 4'b0000;
    end
    else if ( fsm_output[5] ) begin
      butterFly_acc_4_itm_3 <= butterFly_acc_4_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_nor_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_nor_itm_1 <= ~((butterFly_f1_acc_1_tmp!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_nor_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_nor_itm_1 <= ~((butterFly_f1_acc_1_tmp[3:1]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_nor_1_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_nor_1_itm_1 <= ~((butterFly_f1_acc_1_tmp[3]) | (butterFly_f1_acc_1_tmp[2])
          | (butterFly_f1_acc_1_tmp[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_2_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_2_itm_1 <= (butterFly_f1_acc_1_tmp==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_nor_3_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_nor_3_itm_1 <= ~((butterFly_f1_acc_1_tmp[3]) | (butterFly_f1_acc_1_tmp[1])
          | (butterFly_f1_acc_1_tmp[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_4_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_4_itm_1 <= (butterFly_f1_acc_1_tmp==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_5_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_5_itm_1 <= (butterFly_f1_acc_1_tmp==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_6_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_6_itm_1 <= (butterFly_f1_acc_1_tmp==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_nor_6_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_nor_6_itm_1 <= ~((butterFly_f1_acc_1_tmp[2:0]!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_8_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_8_itm_1 <= (butterFly_f1_acc_1_tmp==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_9_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_9_itm_1 <= (butterFly_f1_acc_1_tmp==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_10_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_10_itm_1 <= (butterFly_f1_acc_1_tmp==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_11_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_11_itm_1 <= (butterFly_f1_acc_1_tmp==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_12_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_12_itm_1 <= (butterFly_f1_acc_1_tmp==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_f1_butterFly_f1_and_13_itm_1 <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      butterFly_f1_butterFly_f1_and_13_itm_1 <= (butterFly_f1_acc_1_tmp==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( ~ INNER_LOOP_j_or_cse ) begin
      operator_33_true_return_13_0_sva <= z_out_4[13:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ INNER_LOOP_j_or_cse ) begin
      operator_20_false_rshift_psp_sva <= z_out_5;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_acc_itm_2 <= 4'b0000;
    end
    else if ( fsm_output[5] ) begin
      butterFly_acc_itm_2 <= butterFly_acc_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      INNER_LOOP_stage_0_2 <= 1'b0;
      INNER_LOOP_stage_0_3 <= 1'b0;
      INNER_LOOP_stage_0_4 <= 1'b0;
    end
    else if ( INNER_LOOP_or_1_cse ) begin
      INNER_LOOP_stage_0_2 <= INNER_LOOP_stage_0_1 & (~ (fsm_output[2]));
      INNER_LOOP_stage_0_3 <= INNER_LOOP_stage_0_2 & (~ (fsm_output[2]));
      INNER_LOOP_stage_0_4 <= INNER_LOOP_stage_0_3 & (~ (fsm_output[2]));
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      modulo_add_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_sva_1, modulo_add_qif_acc_nl,
          for_and_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      INNER_LOOP_idx1_acc_psp_sva_2_12_0 <= INNER_LOOP_idx1_acc_psp_sva_1_12_0;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      INNER_LOOP_k_17_0_sva_2_0 <= INNER_LOOP_k_17_0_sva_1_0;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      INNER_LOOP_tf_h_asn_itm_1 <= twiddle_h_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_acc_4_itm_2 <= 4'b0000;
    end
    else if ( fsm_output[5] ) begin
      butterFly_acc_4_itm_2 <= butterFly_acc_4_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_acc_itm_1 <= 4'b0000;
    end
    else if ( fsm_output[5] ) begin
      butterFly_acc_itm_1 <= nl_butterFly_acc_itm_1[3:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly_acc_4_itm_1 <= 4'b0000;
    end
    else if ( fsm_output[5] ) begin
      butterFly_acc_4_itm_1 <= nl_butterFly_acc_4_itm_1[3:0];
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      INNER_LOOP_tf_asn_itm_1 <= twiddle_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( fsm_output[5] ) begin
      butterFly_idx2_17_0_sva_1_13_0 <= butterFly_idx2_17_0_sva_1[13:0];
    end
  end
  always @(posedge clk) begin
    if ( ((butterFly_acc_4_itm_3!=4'b1111)) & INNER_LOOP_stage_0_4 ) begin
      mult_res_lpi_3_dfm <= MUX_v_32_2_2(z_out, z_out_1, z_out_7_32);
    end
  end
  always @(posedge clk) begin
    if ( ~ (fsm_output[4]) ) begin
      tmp_1_lpi_3_dfm <= z_out_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ (fsm_output[4]) ) begin
      INNER_LOOP_k_17_0_sva <= nl_INNER_LOOP_k_17_0_sva[17:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ (fsm_output[4]) ) begin
      mult_z_mul_itm <= nl_mult_z_mul_itm[31:0];
    end
  end
  assign INNER_LOOP_INNER_LOOP_and_nl = INNER_LOOP_stage_0 & (~ (z_out_6[14]));
  assign or_101_nl = ((~(INNER_LOOP_stage_0_1 & (INNER_LOOP_j_13_0_sva_2[13]))) &
      (fsm_output[3])) | (fsm_output[5:4]!=2'b00);
  assign butterFly_mux_nl = MUX_s_1_2_2(INNER_LOOP_INNER_LOOP_and_nl, INNER_LOOP_stage_0,
      or_101_nl);
  assign for_i_for_i_mux_nl = MUX_v_14_2_2((z_out_6[13:0]), butterFly_idx2_17_0_sva_1_13_0,
      fsm_output[5]);
  assign INNER_LOOP_nor_nl = ~(or_dcpl_30 | or_dcpl_29);
  assign nl_operator_20_false_acc_psp_sva  = (~ STAGE_LOOP_i_3_0_sva) + 4'b1111;
  assign nl_modulo_add_qif_acc_nl = modulo_add_base_sva_1 - p_sva;
  assign modulo_add_qif_acc_nl = nl_modulo_add_qif_acc_nl[31:0];
  assign for_and_1_nl = z_out_7_32 & (fsm_output[5]);
  assign nl_butterFly_acc_itm_1  = (INNER_LOOP_idx1_acc_psp_sva_1[16:13]) + STAGE_LOOP_i_3_0_sva
      + 4'b0001;
  assign nl_butterFly_acc_4_itm_1  = (butterFly_idx2_17_0_sva_1[17:14]) + STAGE_LOOP_i_3_0_sva
      + 4'b0001;
  assign nl_INNER_LOOP_k_17_0_sva  = conv_u2u_13_18(INNER_LOOP_j_13_0_sva_12_0) -
      z_out_4;
  assign nl_mult_z_mul_itm  = mult_t_mul_cmp_a * INNER_LOOP_tf_asn_itm_2;
  assign modulo_sub_qif_modulo_sub_qif_or_1_nl = (z_out_1[31]) | (~ (fsm_output[3]));
  assign modulo_sub_qif_or_1_nl = (~ (fsm_output[5])) | (fsm_output[3]);
  assign modulo_sub_qif_mux_2_nl = MUX_v_32_2_2(p_sva, (~ p_sva), fsm_output[3]);
  assign nl_acc_nl = ({modulo_sub_qif_modulo_sub_qif_or_1_nl , (z_out_1[30:0]) ,
      modulo_sub_qif_or_1_nl}) + ({modulo_sub_qif_mux_2_nl , 1'b1});
  assign acc_nl = nl_acc_nl[32:0];
  assign z_out = readslicef_33_32_1(acc_nl);
  assign mult_res_mux_3_nl = MUX_v_32_2_2((~ mult_z_mul_itm_1_1), (~ tmp_1_lpi_3_dfm),
      fsm_output[5]);
  assign nl_acc_1_nl = ({mult_z_mul_itm_1 , 1'b1}) + ({mult_res_mux_3_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[32:0];
  assign z_out_1 = readslicef_33_32_1(acc_1_nl);
  assign mult_z_mux_2_nl = MUX_v_32_2_2(operator_96_false_operator_96_false_slc_mult_t_mul_51_20_itm,
      ({19'b0000000000000000000 , INNER_LOOP_g_rshift_psp_sva}), fsm_output[4]);
  assign mult_z_mux_3_nl = MUX_v_32_2_2(p_sva, ({18'b000000000000000000 , operator_20_false_rshift_psp_sva}),
      fsm_output[4]);
  assign nl_z_out_3 = mult_z_mux_2_nl * mult_z_mux_3_nl;
  assign z_out_3 = nl_z_out_3[31:0];
  assign STAGE_LOOP_mux_1_nl = MUX_v_14_2_2(({10'b0000000000 , STAGE_LOOP_i_3_0_sva}),
      butterFly_idx2_17_0_sva_2_13_0, fsm_output[1]);
  assign nl_z_out_6 = conv_u2u_14_15(STAGE_LOOP_mux_1_nl) + 15'b000000000000001;
  assign z_out_6 = nl_z_out_6[14:0];
  assign modulo_add_mux_3_nl = MUX_v_32_2_2(p_sva, z_out_1, fsm_output[3]);
  assign modulo_add_mux_4_nl = MUX_v_32_2_2((~ modulo_add_base_sva_1), (~ p_sva),
      fsm_output[3]);
  assign nl_acc_3_nl = ({1'b1 , modulo_add_mux_3_nl , 1'b1}) + conv_u2u_33_34({modulo_add_mux_4_nl
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[33:0];
  assign z_out_7_32 = readslicef_34_1_33(acc_3_nl);
  assign butterFly_f1_mux_32_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_nor_itm_1,
      butterFly_f2_butterFly_f2_nor_itm_1, fsm_output[3]);
  assign butterFly_f1_butterFly_f1_and_14_nl = (reg_butterFly_f1_acc_1_svs_st_1_cse[0])
      & butterFly_f1_nor_itm_1;
  assign butterFly_f2_butterFly_f2_and_14_nl = (butterFly_f2_acc_1_svs_1[0]) & butterFly_f2_nor_itm_1;
  assign butterFly_f1_mux_33_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_14_nl,
      butterFly_f2_butterFly_f2_and_14_nl, fsm_output[3]);
  assign butterFly_f1_butterFly_f1_and_15_nl = (reg_butterFly_f1_acc_1_svs_st_1_cse[1])
      & butterFly_f1_nor_1_itm_1;
  assign butterFly_f2_butterFly_f2_and_15_nl = (butterFly_f2_acc_1_svs_1[1]) & butterFly_f2_nor_1_itm_1;
  assign butterFly_f1_mux_34_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_15_nl,
      butterFly_f2_butterFly_f2_and_15_nl, fsm_output[3]);
  assign butterFly_f1_mux_35_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_2_itm_1,
      butterFly_f2_butterFly_f2_and_2_itm_1, fsm_output[3]);
  assign butterFly_f1_butterFly_f1_and_16_nl = (reg_butterFly_f1_acc_1_svs_st_1_cse[2])
      & butterFly_f1_nor_3_itm_1;
  assign butterFly_f2_butterFly_f2_and_16_nl = (butterFly_f2_acc_1_svs_1[2]) & butterFly_f2_nor_3_itm_1;
  assign butterFly_f1_mux_36_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_16_nl,
      butterFly_f2_butterFly_f2_and_16_nl, fsm_output[3]);
  assign butterFly_f1_mux_37_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_4_itm_1,
      butterFly_f2_butterFly_f2_and_4_itm_1, fsm_output[3]);
  assign butterFly_f1_mux_38_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_5_itm_1,
      butterFly_f2_butterFly_f2_and_5_itm_1, fsm_output[3]);
  assign butterFly_f1_mux_39_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_6_itm_1,
      butterFly_f2_butterFly_f2_and_6_itm_1, fsm_output[3]);
  assign butterFly_f1_butterFly_f1_and_17_nl = (reg_butterFly_f1_acc_1_svs_st_1_cse[3])
      & butterFly_f1_nor_6_itm_1;
  assign butterFly_f2_butterFly_f2_and_17_nl = (butterFly_f2_acc_1_svs_1[3]) & butterFly_f2_nor_6_itm_1;
  assign butterFly_f1_mux_40_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_17_nl,
      butterFly_f2_butterFly_f2_and_17_nl, fsm_output[3]);
  assign butterFly_f1_mux_41_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_8_itm_1,
      butterFly_f2_butterFly_f2_and_8_itm_1, fsm_output[3]);
  assign butterFly_f1_mux_42_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_9_itm_1,
      butterFly_f2_butterFly_f2_and_9_itm_1, fsm_output[3]);
  assign butterFly_f1_mux_43_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_10_itm_1,
      butterFly_f2_butterFly_f2_and_10_itm_1, fsm_output[3]);
  assign butterFly_f1_mux_44_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_11_itm_1,
      butterFly_f2_butterFly_f2_and_11_itm_1, fsm_output[3]);
  assign butterFly_f1_mux_45_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_12_itm_1,
      butterFly_f2_butterFly_f2_and_12_itm_1, fsm_output[3]);
  assign butterFly_f1_mux_46_nl = MUX_s_1_2_2(butterFly_f1_butterFly_f1_and_13_itm_1,
      butterFly_f2_butterFly_f2_and_13_itm_1, fsm_output[3]);
  assign z_out_2 = MUX1HOT_v_32_15_2(result_rsc_0_0_i_q_d, result_rsc_1_0_i_q_d,
      result_rsc_2_0_i_q_d, result_rsc_3_0_i_q_d, result_rsc_4_0_i_q_d, result_rsc_5_0_i_q_d,
      result_rsc_6_0_i_q_d, result_rsc_7_0_i_q_d, result_rsc_8_0_i_q_d, result_rsc_9_0_i_q_d,
      result_rsc_10_0_i_q_d, result_rsc_11_0_i_q_d, result_rsc_12_0_i_q_d, result_rsc_13_0_i_q_d,
      result_rsc_14_0_i_q_d, {butterFly_f1_mux_32_nl , butterFly_f1_mux_33_nl , butterFly_f1_mux_34_nl
      , butterFly_f1_mux_35_nl , butterFly_f1_mux_36_nl , butterFly_f1_mux_37_nl
      , butterFly_f1_mux_38_nl , butterFly_f1_mux_39_nl , butterFly_f1_mux_40_nl
      , butterFly_f1_mux_41_nl , butterFly_f1_mux_42_nl , butterFly_f1_mux_43_nl
      , butterFly_f1_mux_44_nl , butterFly_f1_mux_45_nl , butterFly_f1_mux_46_nl});

  function automatic [31:0] MUX1HOT_v_32_15_2;
    input [31:0] input_14;
    input [31:0] input_13;
    input [31:0] input_12;
    input [31:0] input_11;
    input [31:0] input_10;
    input [31:0] input_9;
    input [31:0] input_8;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [14:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    result = result | ( input_8 & {32{sel[8]}});
    result = result | ( input_9 & {32{sel[9]}});
    result = result | ( input_10 & {32{sel[10]}});
    result = result | ( input_11 & {32{sel[11]}});
    result = result | ( input_12 & {32{sel[12]}});
    result = result | ( input_13 & {32{sel[13]}});
    result = result | ( input_14 & {32{sel[14]}});
    MUX1HOT_v_32_15_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input [0:0] sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input [0:0] sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [31:0] readslicef_33_32_1;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_33_32_1 = tmp[31:0];
  end
  endfunction


  function automatic [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [14:0] conv_u2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2s_14_15 =  {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_13_18 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_18 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [14:0] conv_u2u_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_15 = {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_14_18 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_18 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ntt_flat
// ------------------------------------------------------------------


module ntt_flat (
  clk, rst, vec_rsc_radr, vec_rsc_q, vec_rsc_triosy_lz, p_rsc_dat, p_rsc_triosy_lz,
      r_rsc_dat, r_rsc_triosy_lz, twiddle_rsc_radr, twiddle_rsc_q, twiddle_rsc_triosy_lz,
      twiddle_h_rsc_radr, twiddle_h_rsc_q, twiddle_h_rsc_triosy_lz, result_rsc_0_0_wadr,
      result_rsc_0_0_d, result_rsc_0_0_we, result_rsc_0_0_radr, result_rsc_0_0_q,
      result_rsc_triosy_0_0_lz, result_rsc_1_0_wadr, result_rsc_1_0_d, result_rsc_1_0_we,
      result_rsc_1_0_radr, result_rsc_1_0_q, result_rsc_triosy_1_0_lz, result_rsc_2_0_wadr,
      result_rsc_2_0_d, result_rsc_2_0_we, result_rsc_2_0_radr, result_rsc_2_0_q,
      result_rsc_triosy_2_0_lz, result_rsc_3_0_wadr, result_rsc_3_0_d, result_rsc_3_0_we,
      result_rsc_3_0_radr, result_rsc_3_0_q, result_rsc_triosy_3_0_lz, result_rsc_4_0_wadr,
      result_rsc_4_0_d, result_rsc_4_0_we, result_rsc_4_0_radr, result_rsc_4_0_q,
      result_rsc_triosy_4_0_lz, result_rsc_5_0_wadr, result_rsc_5_0_d, result_rsc_5_0_we,
      result_rsc_5_0_radr, result_rsc_5_0_q, result_rsc_triosy_5_0_lz, result_rsc_6_0_wadr,
      result_rsc_6_0_d, result_rsc_6_0_we, result_rsc_6_0_radr, result_rsc_6_0_q,
      result_rsc_triosy_6_0_lz, result_rsc_7_0_wadr, result_rsc_7_0_d, result_rsc_7_0_we,
      result_rsc_7_0_radr, result_rsc_7_0_q, result_rsc_triosy_7_0_lz, result_rsc_8_0_wadr,
      result_rsc_8_0_d, result_rsc_8_0_we, result_rsc_8_0_radr, result_rsc_8_0_q,
      result_rsc_triosy_8_0_lz, result_rsc_9_0_wadr, result_rsc_9_0_d, result_rsc_9_0_we,
      result_rsc_9_0_radr, result_rsc_9_0_q, result_rsc_triosy_9_0_lz, result_rsc_10_0_wadr,
      result_rsc_10_0_d, result_rsc_10_0_we, result_rsc_10_0_radr, result_rsc_10_0_q,
      result_rsc_triosy_10_0_lz, result_rsc_11_0_wadr, result_rsc_11_0_d, result_rsc_11_0_we,
      result_rsc_11_0_radr, result_rsc_11_0_q, result_rsc_triosy_11_0_lz, result_rsc_12_0_wadr,
      result_rsc_12_0_d, result_rsc_12_0_we, result_rsc_12_0_radr, result_rsc_12_0_q,
      result_rsc_triosy_12_0_lz, result_rsc_13_0_wadr, result_rsc_13_0_d, result_rsc_13_0_we,
      result_rsc_13_0_radr, result_rsc_13_0_q, result_rsc_triosy_13_0_lz, result_rsc_14_0_wadr,
      result_rsc_14_0_d, result_rsc_14_0_we, result_rsc_14_0_radr, result_rsc_14_0_q,
      result_rsc_triosy_14_0_lz
);
  input clk;
  input rst;
  output [13:0] vec_rsc_radr;
  input [31:0] vec_rsc_q;
  output vec_rsc_triosy_lz;
  input [31:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [31:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  output [13:0] twiddle_rsc_radr;
  input [31:0] twiddle_rsc_q;
  output twiddle_rsc_triosy_lz;
  output [13:0] twiddle_h_rsc_radr;
  input [31:0] twiddle_h_rsc_q;
  output twiddle_h_rsc_triosy_lz;
  output [13:0] result_rsc_0_0_wadr;
  output [31:0] result_rsc_0_0_d;
  output result_rsc_0_0_we;
  output [13:0] result_rsc_0_0_radr;
  input [31:0] result_rsc_0_0_q;
  output result_rsc_triosy_0_0_lz;
  output [13:0] result_rsc_1_0_wadr;
  output [31:0] result_rsc_1_0_d;
  output result_rsc_1_0_we;
  output [13:0] result_rsc_1_0_radr;
  input [31:0] result_rsc_1_0_q;
  output result_rsc_triosy_1_0_lz;
  output [13:0] result_rsc_2_0_wadr;
  output [31:0] result_rsc_2_0_d;
  output result_rsc_2_0_we;
  output [13:0] result_rsc_2_0_radr;
  input [31:0] result_rsc_2_0_q;
  output result_rsc_triosy_2_0_lz;
  output [13:0] result_rsc_3_0_wadr;
  output [31:0] result_rsc_3_0_d;
  output result_rsc_3_0_we;
  output [13:0] result_rsc_3_0_radr;
  input [31:0] result_rsc_3_0_q;
  output result_rsc_triosy_3_0_lz;
  output [13:0] result_rsc_4_0_wadr;
  output [31:0] result_rsc_4_0_d;
  output result_rsc_4_0_we;
  output [13:0] result_rsc_4_0_radr;
  input [31:0] result_rsc_4_0_q;
  output result_rsc_triosy_4_0_lz;
  output [13:0] result_rsc_5_0_wadr;
  output [31:0] result_rsc_5_0_d;
  output result_rsc_5_0_we;
  output [13:0] result_rsc_5_0_radr;
  input [31:0] result_rsc_5_0_q;
  output result_rsc_triosy_5_0_lz;
  output [13:0] result_rsc_6_0_wadr;
  output [31:0] result_rsc_6_0_d;
  output result_rsc_6_0_we;
  output [13:0] result_rsc_6_0_radr;
  input [31:0] result_rsc_6_0_q;
  output result_rsc_triosy_6_0_lz;
  output [13:0] result_rsc_7_0_wadr;
  output [31:0] result_rsc_7_0_d;
  output result_rsc_7_0_we;
  output [13:0] result_rsc_7_0_radr;
  input [31:0] result_rsc_7_0_q;
  output result_rsc_triosy_7_0_lz;
  output [13:0] result_rsc_8_0_wadr;
  output [31:0] result_rsc_8_0_d;
  output result_rsc_8_0_we;
  output [13:0] result_rsc_8_0_radr;
  input [31:0] result_rsc_8_0_q;
  output result_rsc_triosy_8_0_lz;
  output [13:0] result_rsc_9_0_wadr;
  output [31:0] result_rsc_9_0_d;
  output result_rsc_9_0_we;
  output [13:0] result_rsc_9_0_radr;
  input [31:0] result_rsc_9_0_q;
  output result_rsc_triosy_9_0_lz;
  output [13:0] result_rsc_10_0_wadr;
  output [31:0] result_rsc_10_0_d;
  output result_rsc_10_0_we;
  output [13:0] result_rsc_10_0_radr;
  input [31:0] result_rsc_10_0_q;
  output result_rsc_triosy_10_0_lz;
  output [13:0] result_rsc_11_0_wadr;
  output [31:0] result_rsc_11_0_d;
  output result_rsc_11_0_we;
  output [13:0] result_rsc_11_0_radr;
  input [31:0] result_rsc_11_0_q;
  output result_rsc_triosy_11_0_lz;
  output [13:0] result_rsc_12_0_wadr;
  output [31:0] result_rsc_12_0_d;
  output result_rsc_12_0_we;
  output [13:0] result_rsc_12_0_radr;
  input [31:0] result_rsc_12_0_q;
  output result_rsc_triosy_12_0_lz;
  output [13:0] result_rsc_13_0_wadr;
  output [31:0] result_rsc_13_0_d;
  output result_rsc_13_0_we;
  output [13:0] result_rsc_13_0_radr;
  input [31:0] result_rsc_13_0_q;
  output result_rsc_triosy_13_0_lz;
  output [13:0] result_rsc_14_0_wadr;
  output [31:0] result_rsc_14_0_d;
  output result_rsc_14_0_we;
  output [13:0] result_rsc_14_0_radr;
  input [31:0] result_rsc_14_0_q;
  output result_rsc_triosy_14_0_lz;


  // Interconnect Declarations
  wire [31:0] vec_rsci_q_d;
  wire [13:0] vec_rsci_radr_d;
  wire vec_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] twiddle_rsci_q_d;
  wire [31:0] twiddle_h_rsci_q_d;
  wire [31:0] result_rsc_0_0_i_d_d;
  wire [31:0] result_rsc_0_0_i_q_d;
  wire [13:0] result_rsc_0_0_i_wadr_d;
  wire result_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_1_0_i_q_d;
  wire result_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_2_0_i_q_d;
  wire result_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_3_0_i_q_d;
  wire result_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_4_0_i_q_d;
  wire result_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_5_0_i_q_d;
  wire result_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_6_0_i_q_d;
  wire result_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_7_0_i_q_d;
  wire result_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_8_0_i_q_d;
  wire result_rsc_8_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_9_0_i_q_d;
  wire result_rsc_9_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_10_0_i_q_d;
  wire result_rsc_10_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_11_0_i_q_d;
  wire result_rsc_11_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_12_0_i_q_d;
  wire result_rsc_12_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_13_0_i_q_d;
  wire result_rsc_13_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] result_rsc_14_0_i_q_d;
  wire result_rsc_14_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] mult_t_mul_cmp_a;
  wire [31:0] mult_t_mul_cmp_b;
  wire [13:0] twiddle_rsci_radr_d_iff;
  wire twiddle_rsci_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire [13:0] result_rsc_0_0_i_radr_d_iff;
  wire result_rsc_0_0_i_we_d_iff;
  wire [31:0] result_rsc_1_0_i_d_d_iff;
  wire result_rsc_1_0_i_we_d_iff;
  wire result_rsc_2_0_i_we_d_iff;
  wire result_rsc_3_0_i_we_d_iff;
  wire result_rsc_4_0_i_we_d_iff;
  wire result_rsc_5_0_i_we_d_iff;
  wire result_rsc_6_0_i_we_d_iff;
  wire result_rsc_7_0_i_we_d_iff;
  wire result_rsc_8_0_i_we_d_iff;
  wire result_rsc_9_0_i_we_d_iff;
  wire result_rsc_10_0_i_we_d_iff;
  wire result_rsc_11_0_i_we_d_iff;
  wire result_rsc_12_0_i_we_d_iff;
  wire result_rsc_13_0_i_we_d_iff;
  wire result_rsc_14_0_i_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [51:0] nl_ntt_flat_core_inst_mult_t_mul_cmp_z;
  assign nl_ntt_flat_core_inst_mult_t_mul_cmp_z = conv_u2u_64_52(mult_t_mul_cmp_a
      * mult_t_mul_cmp_b);
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_1_14_32_16384_16384_32_1_gen vec_rsci
      (
      .q(vec_rsc_q),
      .radr(vec_rsc_radr),
      .q_d(vec_rsci_q_d),
      .radr_d(vec_rsci_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_4_14_32_16384_16384_32_1_gen twiddle_rsci
      (
      .q(twiddle_rsc_q),
      .radr(twiddle_rsc_radr),
      .q_d(twiddle_rsci_q_d),
      .radr_d(twiddle_rsci_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsci_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_5_14_32_16384_16384_32_1_gen twiddle_h_rsci
      (
      .q(twiddle_h_rsc_q),
      .radr(twiddle_h_rsc_radr),
      .q_d(twiddle_h_rsci_q_d),
      .radr_d(twiddle_rsci_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsci_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_7_14_32_16384_16384_32_1_gen result_rsc_0_0_i
      (
      .q(result_rsc_0_0_q),
      .radr(result_rsc_0_0_radr),
      .we(result_rsc_0_0_we),
      .d(result_rsc_0_0_d),
      .wadr(result_rsc_0_0_wadr),
      .d_d(result_rsc_0_0_i_d_d),
      .q_d(result_rsc_0_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_14_32_16384_16384_32_1_gen result_rsc_1_0_i
      (
      .q(result_rsc_1_0_q),
      .radr(result_rsc_1_0_radr),
      .we(result_rsc_1_0_we),
      .d(result_rsc_1_0_d),
      .wadr(result_rsc_1_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_1_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_14_32_16384_16384_32_1_gen result_rsc_2_0_i
      (
      .q(result_rsc_2_0_q),
      .radr(result_rsc_2_0_radr),
      .we(result_rsc_2_0_we),
      .d(result_rsc_2_0_d),
      .wadr(result_rsc_2_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_2_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_14_32_16384_16384_32_1_gen result_rsc_3_0_i
      (
      .q(result_rsc_3_0_q),
      .radr(result_rsc_3_0_radr),
      .we(result_rsc_3_0_we),
      .d(result_rsc_3_0_d),
      .wadr(result_rsc_3_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_3_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_14_32_16384_16384_32_1_gen result_rsc_4_0_i
      (
      .q(result_rsc_4_0_q),
      .radr(result_rsc_4_0_radr),
      .we(result_rsc_4_0_we),
      .d(result_rsc_4_0_d),
      .wadr(result_rsc_4_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_4_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_14_32_16384_16384_32_1_gen result_rsc_5_0_i
      (
      .q(result_rsc_5_0_q),
      .radr(result_rsc_5_0_radr),
      .we(result_rsc_5_0_we),
      .d(result_rsc_5_0_d),
      .wadr(result_rsc_5_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_5_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_14_32_16384_16384_32_1_gen result_rsc_6_0_i
      (
      .q(result_rsc_6_0_q),
      .radr(result_rsc_6_0_radr),
      .we(result_rsc_6_0_we),
      .d(result_rsc_6_0_d),
      .wadr(result_rsc_6_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_6_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_14_32_16384_16384_32_1_gen result_rsc_7_0_i
      (
      .q(result_rsc_7_0_q),
      .radr(result_rsc_7_0_radr),
      .we(result_rsc_7_0_we),
      .d(result_rsc_7_0_d),
      .wadr(result_rsc_7_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_7_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_14_32_16384_16384_32_1_gen result_rsc_8_0_i
      (
      .q(result_rsc_8_0_q),
      .radr(result_rsc_8_0_radr),
      .we(result_rsc_8_0_we),
      .d(result_rsc_8_0_d),
      .wadr(result_rsc_8_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_8_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_8_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_8_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_8_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_14_32_16384_16384_32_1_gen result_rsc_9_0_i
      (
      .q(result_rsc_9_0_q),
      .radr(result_rsc_9_0_radr),
      .we(result_rsc_9_0_we),
      .d(result_rsc_9_0_d),
      .wadr(result_rsc_9_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_9_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_9_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_9_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_9_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_14_32_16384_16384_32_1_gen result_rsc_10_0_i
      (
      .q(result_rsc_10_0_q),
      .radr(result_rsc_10_0_radr),
      .we(result_rsc_10_0_we),
      .d(result_rsc_10_0_d),
      .wadr(result_rsc_10_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_10_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_10_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_10_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_10_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_14_32_16384_16384_32_1_gen result_rsc_11_0_i
      (
      .q(result_rsc_11_0_q),
      .radr(result_rsc_11_0_radr),
      .we(result_rsc_11_0_we),
      .d(result_rsc_11_0_d),
      .wadr(result_rsc_11_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_11_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_11_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_11_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_11_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_14_32_16384_16384_32_1_gen result_rsc_12_0_i
      (
      .q(result_rsc_12_0_q),
      .radr(result_rsc_12_0_radr),
      .we(result_rsc_12_0_we),
      .d(result_rsc_12_0_d),
      .wadr(result_rsc_12_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_12_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_12_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_12_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_12_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_14_32_16384_16384_32_1_gen result_rsc_13_0_i
      (
      .q(result_rsc_13_0_q),
      .radr(result_rsc_13_0_radr),
      .we(result_rsc_13_0_we),
      .d(result_rsc_13_0_d),
      .wadr(result_rsc_13_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_13_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_13_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_13_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_13_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_14_32_16384_16384_32_1_gen result_rsc_14_0_i
      (
      .q(result_rsc_14_0_q),
      .radr(result_rsc_14_0_radr),
      .we(result_rsc_14_0_we),
      .d(result_rsc_14_0_d),
      .wadr(result_rsc_14_0_wadr),
      .d_d(result_rsc_1_0_i_d_d_iff),
      .q_d(result_rsc_14_0_i_q_d),
      .radr_d(result_rsc_0_0_i_radr_d_iff),
      .wadr_d(result_rsc_0_0_i_wadr_d),
      .we_d(result_rsc_14_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(result_rsc_14_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(result_rsc_14_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  ntt_flat_core ntt_flat_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_lz(vec_rsc_triosy_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .twiddle_rsc_triosy_lz(twiddle_rsc_triosy_lz),
      .twiddle_h_rsc_triosy_lz(twiddle_h_rsc_triosy_lz),
      .result_rsc_triosy_0_0_lz(result_rsc_triosy_0_0_lz),
      .result_rsc_triosy_1_0_lz(result_rsc_triosy_1_0_lz),
      .result_rsc_triosy_2_0_lz(result_rsc_triosy_2_0_lz),
      .result_rsc_triosy_3_0_lz(result_rsc_triosy_3_0_lz),
      .result_rsc_triosy_4_0_lz(result_rsc_triosy_4_0_lz),
      .result_rsc_triosy_5_0_lz(result_rsc_triosy_5_0_lz),
      .result_rsc_triosy_6_0_lz(result_rsc_triosy_6_0_lz),
      .result_rsc_triosy_7_0_lz(result_rsc_triosy_7_0_lz),
      .result_rsc_triosy_8_0_lz(result_rsc_triosy_8_0_lz),
      .result_rsc_triosy_9_0_lz(result_rsc_triosy_9_0_lz),
      .result_rsc_triosy_10_0_lz(result_rsc_triosy_10_0_lz),
      .result_rsc_triosy_11_0_lz(result_rsc_triosy_11_0_lz),
      .result_rsc_triosy_12_0_lz(result_rsc_triosy_12_0_lz),
      .result_rsc_triosy_13_0_lz(result_rsc_triosy_13_0_lz),
      .result_rsc_triosy_14_0_lz(result_rsc_triosy_14_0_lz),
      .vec_rsci_q_d(vec_rsci_q_d),
      .vec_rsci_radr_d(vec_rsci_radr_d),
      .vec_rsci_readA_r_ram_ir_internal_RMASK_B_d(vec_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsci_q_d(twiddle_rsci_q_d),
      .twiddle_h_rsci_q_d(twiddle_h_rsci_q_d),
      .result_rsc_0_0_i_d_d(result_rsc_0_0_i_d_d),
      .result_rsc_0_0_i_q_d(result_rsc_0_0_i_q_d),
      .result_rsc_0_0_i_wadr_d(result_rsc_0_0_i_wadr_d),
      .result_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_1_0_i_q_d(result_rsc_1_0_i_q_d),
      .result_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_2_0_i_q_d(result_rsc_2_0_i_q_d),
      .result_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_3_0_i_q_d(result_rsc_3_0_i_q_d),
      .result_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_4_0_i_q_d(result_rsc_4_0_i_q_d),
      .result_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_5_0_i_q_d(result_rsc_5_0_i_q_d),
      .result_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_6_0_i_q_d(result_rsc_6_0_i_q_d),
      .result_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_7_0_i_q_d(result_rsc_7_0_i_q_d),
      .result_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_8_0_i_q_d(result_rsc_8_0_i_q_d),
      .result_rsc_8_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_8_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_9_0_i_q_d(result_rsc_9_0_i_q_d),
      .result_rsc_9_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_9_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_10_0_i_q_d(result_rsc_10_0_i_q_d),
      .result_rsc_10_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_10_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_11_0_i_q_d(result_rsc_11_0_i_q_d),
      .result_rsc_11_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_11_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_12_0_i_q_d(result_rsc_12_0_i_q_d),
      .result_rsc_12_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_12_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_13_0_i_q_d(result_rsc_13_0_i_q_d),
      .result_rsc_13_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_13_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .result_rsc_14_0_i_q_d(result_rsc_14_0_i_q_d),
      .result_rsc_14_0_i_readA_r_ram_ir_internal_RMASK_B_d(result_rsc_14_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .mult_t_mul_cmp_a(mult_t_mul_cmp_a),
      .mult_t_mul_cmp_b(mult_t_mul_cmp_b),
      .mult_t_mul_cmp_z(nl_ntt_flat_core_inst_mult_t_mul_cmp_z[51:0]),
      .twiddle_rsci_radr_d_pff(twiddle_rsci_radr_d_iff),
      .twiddle_rsci_readA_r_ram_ir_internal_RMASK_B_d_pff(twiddle_rsci_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .result_rsc_0_0_i_radr_d_pff(result_rsc_0_0_i_radr_d_iff),
      .result_rsc_0_0_i_we_d_pff(result_rsc_0_0_i_we_d_iff),
      .result_rsc_1_0_i_d_d_pff(result_rsc_1_0_i_d_d_iff),
      .result_rsc_1_0_i_we_d_pff(result_rsc_1_0_i_we_d_iff),
      .result_rsc_2_0_i_we_d_pff(result_rsc_2_0_i_we_d_iff),
      .result_rsc_3_0_i_we_d_pff(result_rsc_3_0_i_we_d_iff),
      .result_rsc_4_0_i_we_d_pff(result_rsc_4_0_i_we_d_iff),
      .result_rsc_5_0_i_we_d_pff(result_rsc_5_0_i_we_d_iff),
      .result_rsc_6_0_i_we_d_pff(result_rsc_6_0_i_we_d_iff),
      .result_rsc_7_0_i_we_d_pff(result_rsc_7_0_i_we_d_iff),
      .result_rsc_8_0_i_we_d_pff(result_rsc_8_0_i_we_d_iff),
      .result_rsc_9_0_i_we_d_pff(result_rsc_9_0_i_we_d_iff),
      .result_rsc_10_0_i_we_d_pff(result_rsc_10_0_i_we_d_iff),
      .result_rsc_11_0_i_we_d_pff(result_rsc_11_0_i_we_d_iff),
      .result_rsc_12_0_i_we_d_pff(result_rsc_12_0_i_we_d_iff),
      .result_rsc_13_0_i_we_d_pff(result_rsc_13_0_i_we_d_iff),
      .result_rsc_14_0_i_we_d_pff(result_rsc_14_0_i_we_d_iff)
    );

  function automatic [51:0] conv_u2u_64_52 ;
    input [63:0]  vector ;
  begin
    conv_u2u_64_52 = vector[51:0];
  end
  endfunction

endmodule



