
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_out_dreg_pkg_v2 IS

COMPONENT mgc_out_dreg_v2
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_out_dreg_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_out_dreg_v2 IS
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END mgc_out_dreg_v2;

ARCHITECTURE beh OF mgc_out_dreg_v2 IS
BEGIN

  z <= d;

END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_rem IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END mgc_rem;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_rem IS
BEGIN
  z <= std_logic_vector(unsigned(a) rem unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) rem   signed(b));
END beh;

--------> ../td_ccore_solutions/modulo_dev_d3e65941ee7586d7daaa2e36d0d005555a5b_0/rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Thu Aug 26 01:37:25 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    modulo_dev_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_dev_core IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_dev_core;

ARCHITECTURE v1 OF modulo_dev_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL base_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat : STD_LOGIC;
  SIGNAL result_rem_12_cmp_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_result_acc_tmp : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_dcpl_1 : STD_LOGIC;
  SIGNAL and_dcpl_2 : STD_LOGIC;
  SIGNAL and_dcpl_3 : STD_LOGIC;
  SIGNAL and_dcpl_4 : STD_LOGIC;
  SIGNAL and_dcpl_6 : STD_LOGIC;
  SIGNAL and_dcpl_8 : STD_LOGIC;
  SIGNAL and_dcpl_9 : STD_LOGIC;
  SIGNAL and_dcpl_11 : STD_LOGIC;
  SIGNAL and_dcpl_13 : STD_LOGIC;
  SIGNAL and_dcpl_18 : STD_LOGIC;
  SIGNAL and_dcpl_26 : STD_LOGIC;
  SIGNAL and_dcpl_27 : STD_LOGIC;
  SIGNAL and_dcpl_28 : STD_LOGIC;
  SIGNAL and_dcpl_29 : STD_LOGIC;
  SIGNAL and_dcpl_30 : STD_LOGIC;
  SIGNAL and_dcpl_31 : STD_LOGIC;
  SIGNAL and_dcpl_32 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_34 : STD_LOGIC;
  SIGNAL and_dcpl_35 : STD_LOGIC;
  SIGNAL and_dcpl_36 : STD_LOGIC;
  SIGNAL and_dcpl_37 : STD_LOGIC;
  SIGNAL and_dcpl_38 : STD_LOGIC;
  SIGNAL and_dcpl_39 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_41 : STD_LOGIC;
  SIGNAL and_dcpl_42 : STD_LOGIC;
  SIGNAL and_dcpl_43 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_47 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL and_dcpl_51 : STD_LOGIC;
  SIGNAL and_dcpl_52 : STD_LOGIC;
  SIGNAL and_dcpl_53 : STD_LOGIC;
  SIGNAL and_dcpl_54 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_56 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_59 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_dcpl_68 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_73 : STD_LOGIC;
  SIGNAL and_dcpl_74 : STD_LOGIC;
  SIGNAL and_dcpl_75 : STD_LOGIC;
  SIGNAL and_dcpl_76 : STD_LOGIC;
  SIGNAL and_dcpl_77 : STD_LOGIC;
  SIGNAL and_dcpl_78 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL and_dcpl_80 : STD_LOGIC;
  SIGNAL and_dcpl_81 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_86 : STD_LOGIC;
  SIGNAL and_dcpl_88 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_96 : STD_LOGIC;
  SIGNAL and_dcpl_98 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_100 : STD_LOGIC;
  SIGNAL and_dcpl_101 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_105 : STD_LOGIC;
  SIGNAL and_dcpl_106 : STD_LOGIC;
  SIGNAL and_dcpl_107 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_113 : STD_LOGIC;
  SIGNAL and_dcpl_114 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_116 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_118 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL and_dcpl_120 : STD_LOGIC;
  SIGNAL and_dcpl_122 : STD_LOGIC;
  SIGNAL and_dcpl_125 : STD_LOGIC;
  SIGNAL and_dcpl_127 : STD_LOGIC;
  SIGNAL and_dcpl_128 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL and_dcpl_130 : STD_LOGIC;
  SIGNAL and_dcpl_131 : STD_LOGIC;
  SIGNAL and_dcpl_132 : STD_LOGIC;
  SIGNAL and_dcpl_133 : STD_LOGIC;
  SIGNAL and_dcpl_134 : STD_LOGIC;
  SIGNAL and_dcpl_135 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_137 : STD_LOGIC;
  SIGNAL and_dcpl_139 : STD_LOGIC;
  SIGNAL and_dcpl_140 : STD_LOGIC;
  SIGNAL and_dcpl_142 : STD_LOGIC;
  SIGNAL and_dcpl_143 : STD_LOGIC;
  SIGNAL and_dcpl_145 : STD_LOGIC;
  SIGNAL and_dcpl_147 : STD_LOGIC;
  SIGNAL and_dcpl_149 : STD_LOGIC;
  SIGNAL and_dcpl_150 : STD_LOGIC;
  SIGNAL and_dcpl_151 : STD_LOGIC;
  SIGNAL and_dcpl_152 : STD_LOGIC;
  SIGNAL and_dcpl_153 : STD_LOGIC;
  SIGNAL and_dcpl_154 : STD_LOGIC;
  SIGNAL and_dcpl_155 : STD_LOGIC;
  SIGNAL and_dcpl_156 : STD_LOGIC;
  SIGNAL and_dcpl_157 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_159 : STD_LOGIC;
  SIGNAL and_dcpl_160 : STD_LOGIC;
  SIGNAL and_dcpl_161 : STD_LOGIC;
  SIGNAL and_dcpl_162 : STD_LOGIC;
  SIGNAL and_dcpl_163 : STD_LOGIC;
  SIGNAL and_dcpl_165 : STD_LOGIC;
  SIGNAL and_dcpl_166 : STD_LOGIC;
  SIGNAL and_dcpl_168 : STD_LOGIC;
  SIGNAL and_dcpl_170 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_176 : STD_LOGIC;
  SIGNAL and_dcpl_177 : STD_LOGIC;
  SIGNAL and_dcpl_178 : STD_LOGIC;
  SIGNAL and_dcpl_179 : STD_LOGIC;
  SIGNAL and_dcpl_180 : STD_LOGIC;
  SIGNAL and_dcpl_181 : STD_LOGIC;
  SIGNAL and_dcpl_182 : STD_LOGIC;
  SIGNAL and_dcpl_183 : STD_LOGIC;
  SIGNAL and_dcpl_184 : STD_LOGIC;
  SIGNAL and_dcpl_185 : STD_LOGIC;
  SIGNAL and_dcpl_186 : STD_LOGIC;
  SIGNAL and_dcpl_187 : STD_LOGIC;
  SIGNAL and_dcpl_188 : STD_LOGIC;
  SIGNAL and_dcpl_189 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_194 : STD_LOGIC;
  SIGNAL and_dcpl_196 : STD_LOGIC;
  SIGNAL and_dcpl_197 : STD_LOGIC;
  SIGNAL and_dcpl_199 : STD_LOGIC;
  SIGNAL and_dcpl_201 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_203 : STD_LOGIC;
  SIGNAL and_dcpl_204 : STD_LOGIC;
  SIGNAL and_dcpl_205 : STD_LOGIC;
  SIGNAL and_dcpl_206 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL and_dcpl_208 : STD_LOGIC;
  SIGNAL and_dcpl_209 : STD_LOGIC;
  SIGNAL and_dcpl_211 : STD_LOGIC;
  SIGNAL and_dcpl_212 : STD_LOGIC;
  SIGNAL and_dcpl_214 : STD_LOGIC;
  SIGNAL and_dcpl_218 : STD_LOGIC;
  SIGNAL and_dcpl_221 : STD_LOGIC;
  SIGNAL and_dcpl_228 : STD_LOGIC;
  SIGNAL and_dcpl_232 : STD_LOGIC;
  SIGNAL and_dcpl_233 : STD_LOGIC;
  SIGNAL and_dcpl_234 : STD_LOGIC;
  SIGNAL and_dcpl_235 : STD_LOGIC;
  SIGNAL and_dcpl_237 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_240 : STD_LOGIC;
  SIGNAL and_dcpl_244 : STD_LOGIC;
  SIGNAL and_dcpl_249 : STD_LOGIC;
  SIGNAL and_dcpl_254 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL and_dcpl_261 : STD_LOGIC;
  SIGNAL and_dcpl_262 : STD_LOGIC;
  SIGNAL and_dcpl_263 : STD_LOGIC;
  SIGNAL or_tmp_2 : STD_LOGIC;
  SIGNAL and_dcpl_269 : STD_LOGIC;
  SIGNAL mux_tmp_1 : STD_LOGIC;
  SIGNAL and_dcpl_275 : STD_LOGIC;
  SIGNAL mux_tmp_3 : STD_LOGIC;
  SIGNAL mux_tmp_4 : STD_LOGIC;
  SIGNAL and_dcpl_281 : STD_LOGIC;
  SIGNAL mux_tmp_6 : STD_LOGIC;
  SIGNAL mux_tmp_7 : STD_LOGIC;
  SIGNAL mux_tmp_8 : STD_LOGIC;
  SIGNAL and_dcpl_287 : STD_LOGIC;
  SIGNAL mux_tmp_10 : STD_LOGIC;
  SIGNAL mux_tmp_11 : STD_LOGIC;
  SIGNAL mux_tmp_12 : STD_LOGIC;
  SIGNAL mux_tmp_13 : STD_LOGIC;
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL mux_tmp_15 : STD_LOGIC;
  SIGNAL mux_tmp_16 : STD_LOGIC;
  SIGNAL mux_tmp_17 : STD_LOGIC;
  SIGNAL mux_tmp_18 : STD_LOGIC;
  SIGNAL mux_tmp_19 : STD_LOGIC;
  SIGNAL and_dcpl_299 : STD_LOGIC;
  SIGNAL mux_tmp_21 : STD_LOGIC;
  SIGNAL mux_tmp_22 : STD_LOGIC;
  SIGNAL mux_tmp_23 : STD_LOGIC;
  SIGNAL mux_tmp_24 : STD_LOGIC;
  SIGNAL mux_tmp_25 : STD_LOGIC;
  SIGNAL mux_tmp_26 : STD_LOGIC;
  SIGNAL and_dcpl_305 : STD_LOGIC;
  SIGNAL mux_tmp_28 : STD_LOGIC;
  SIGNAL mux_tmp_29 : STD_LOGIC;
  SIGNAL mux_tmp_30 : STD_LOGIC;
  SIGNAL mux_tmp_31 : STD_LOGIC;
  SIGNAL mux_tmp_32 : STD_LOGIC;
  SIGNAL mux_tmp_33 : STD_LOGIC;
  SIGNAL mux_tmp_34 : STD_LOGIC;
  SIGNAL and_dcpl_311 : STD_LOGIC;
  SIGNAL and_tmp_6 : STD_LOGIC;
  SIGNAL mux_tmp_36 : STD_LOGIC;
  SIGNAL mux_tmp_37 : STD_LOGIC;
  SIGNAL and_dcpl_318 : STD_LOGIC;
  SIGNAL and_dcpl_319 : STD_LOGIC;
  SIGNAL or_tmp_102 : STD_LOGIC;
  SIGNAL and_dcpl_322 : STD_LOGIC;
  SIGNAL mux_tmp_39 : STD_LOGIC;
  SIGNAL and_dcpl_325 : STD_LOGIC;
  SIGNAL mux_tmp_41 : STD_LOGIC;
  SIGNAL mux_tmp_42 : STD_LOGIC;
  SIGNAL and_dcpl_329 : STD_LOGIC;
  SIGNAL mux_tmp_44 : STD_LOGIC;
  SIGNAL mux_tmp_45 : STD_LOGIC;
  SIGNAL mux_tmp_46 : STD_LOGIC;
  SIGNAL and_dcpl_333 : STD_LOGIC;
  SIGNAL mux_tmp_48 : STD_LOGIC;
  SIGNAL mux_tmp_49 : STD_LOGIC;
  SIGNAL mux_tmp_50 : STD_LOGIC;
  SIGNAL mux_tmp_51 : STD_LOGIC;
  SIGNAL and_dcpl_337 : STD_LOGIC;
  SIGNAL mux_tmp_53 : STD_LOGIC;
  SIGNAL mux_tmp_54 : STD_LOGIC;
  SIGNAL mux_tmp_55 : STD_LOGIC;
  SIGNAL mux_tmp_56 : STD_LOGIC;
  SIGNAL mux_tmp_57 : STD_LOGIC;
  SIGNAL and_dcpl_341 : STD_LOGIC;
  SIGNAL mux_tmp_59 : STD_LOGIC;
  SIGNAL mux_tmp_60 : STD_LOGIC;
  SIGNAL mux_tmp_61 : STD_LOGIC;
  SIGNAL mux_tmp_62 : STD_LOGIC;
  SIGNAL mux_tmp_63 : STD_LOGIC;
  SIGNAL mux_tmp_64 : STD_LOGIC;
  SIGNAL and_dcpl_344 : STD_LOGIC;
  SIGNAL mux_tmp_66 : STD_LOGIC;
  SIGNAL mux_tmp_67 : STD_LOGIC;
  SIGNAL mux_tmp_68 : STD_LOGIC;
  SIGNAL mux_tmp_69 : STD_LOGIC;
  SIGNAL mux_tmp_70 : STD_LOGIC;
  SIGNAL mux_tmp_71 : STD_LOGIC;
  SIGNAL mux_tmp_72 : STD_LOGIC;
  SIGNAL and_dcpl_347 : STD_LOGIC;
  SIGNAL and_tmp_13 : STD_LOGIC;
  SIGNAL mux_tmp_74 : STD_LOGIC;
  SIGNAL mux_tmp_75 : STD_LOGIC;
  SIGNAL and_dcpl_352 : STD_LOGIC;
  SIGNAL and_dcpl_353 : STD_LOGIC;
  SIGNAL or_tmp_202 : STD_LOGIC;
  SIGNAL and_dcpl_357 : STD_LOGIC;
  SIGNAL mux_tmp_77 : STD_LOGIC;
  SIGNAL and_dcpl_361 : STD_LOGIC;
  SIGNAL mux_tmp_79 : STD_LOGIC;
  SIGNAL mux_tmp_80 : STD_LOGIC;
  SIGNAL and_dcpl_364 : STD_LOGIC;
  SIGNAL mux_tmp_82 : STD_LOGIC;
  SIGNAL mux_tmp_83 : STD_LOGIC;
  SIGNAL mux_tmp_84 : STD_LOGIC;
  SIGNAL and_dcpl_367 : STD_LOGIC;
  SIGNAL mux_tmp_86 : STD_LOGIC;
  SIGNAL mux_tmp_87 : STD_LOGIC;
  SIGNAL mux_tmp_88 : STD_LOGIC;
  SIGNAL mux_tmp_89 : STD_LOGIC;
  SIGNAL and_dcpl_370 : STD_LOGIC;
  SIGNAL mux_tmp_91 : STD_LOGIC;
  SIGNAL mux_tmp_92 : STD_LOGIC;
  SIGNAL mux_tmp_93 : STD_LOGIC;
  SIGNAL mux_tmp_94 : STD_LOGIC;
  SIGNAL mux_tmp_95 : STD_LOGIC;
  SIGNAL and_dcpl_373 : STD_LOGIC;
  SIGNAL mux_tmp_97 : STD_LOGIC;
  SIGNAL mux_tmp_98 : STD_LOGIC;
  SIGNAL mux_tmp_99 : STD_LOGIC;
  SIGNAL mux_tmp_100 : STD_LOGIC;
  SIGNAL mux_tmp_101 : STD_LOGIC;
  SIGNAL mux_tmp_102 : STD_LOGIC;
  SIGNAL and_dcpl_377 : STD_LOGIC;
  SIGNAL mux_tmp_104 : STD_LOGIC;
  SIGNAL mux_tmp_105 : STD_LOGIC;
  SIGNAL mux_tmp_106 : STD_LOGIC;
  SIGNAL mux_tmp_107 : STD_LOGIC;
  SIGNAL mux_tmp_108 : STD_LOGIC;
  SIGNAL mux_tmp_109 : STD_LOGIC;
  SIGNAL mux_tmp_110 : STD_LOGIC;
  SIGNAL and_dcpl_381 : STD_LOGIC;
  SIGNAL and_tmp_20 : STD_LOGIC;
  SIGNAL mux_tmp_112 : STD_LOGIC;
  SIGNAL mux_tmp_113 : STD_LOGIC;
  SIGNAL and_dcpl_386 : STD_LOGIC;
  SIGNAL and_dcpl_387 : STD_LOGIC;
  SIGNAL or_tmp_302 : STD_LOGIC;
  SIGNAL and_dcpl_390 : STD_LOGIC;
  SIGNAL mux_tmp_115 : STD_LOGIC;
  SIGNAL and_dcpl_393 : STD_LOGIC;
  SIGNAL mux_tmp_117 : STD_LOGIC;
  SIGNAL mux_tmp_118 : STD_LOGIC;
  SIGNAL and_dcpl_396 : STD_LOGIC;
  SIGNAL mux_tmp_120 : STD_LOGIC;
  SIGNAL mux_tmp_121 : STD_LOGIC;
  SIGNAL mux_tmp_122 : STD_LOGIC;
  SIGNAL and_dcpl_399 : STD_LOGIC;
  SIGNAL mux_tmp_124 : STD_LOGIC;
  SIGNAL mux_tmp_125 : STD_LOGIC;
  SIGNAL mux_tmp_126 : STD_LOGIC;
  SIGNAL mux_tmp_127 : STD_LOGIC;
  SIGNAL and_dcpl_402 : STD_LOGIC;
  SIGNAL mux_tmp_129 : STD_LOGIC;
  SIGNAL mux_tmp_130 : STD_LOGIC;
  SIGNAL mux_tmp_131 : STD_LOGIC;
  SIGNAL mux_tmp_132 : STD_LOGIC;
  SIGNAL mux_tmp_133 : STD_LOGIC;
  SIGNAL and_dcpl_405 : STD_LOGIC;
  SIGNAL mux_tmp_135 : STD_LOGIC;
  SIGNAL mux_tmp_136 : STD_LOGIC;
  SIGNAL mux_tmp_137 : STD_LOGIC;
  SIGNAL mux_tmp_138 : STD_LOGIC;
  SIGNAL mux_tmp_139 : STD_LOGIC;
  SIGNAL mux_tmp_140 : STD_LOGIC;
  SIGNAL and_dcpl_408 : STD_LOGIC;
  SIGNAL mux_tmp_142 : STD_LOGIC;
  SIGNAL mux_tmp_143 : STD_LOGIC;
  SIGNAL mux_tmp_144 : STD_LOGIC;
  SIGNAL mux_tmp_145 : STD_LOGIC;
  SIGNAL mux_tmp_146 : STD_LOGIC;
  SIGNAL mux_tmp_147 : STD_LOGIC;
  SIGNAL mux_tmp_148 : STD_LOGIC;
  SIGNAL and_dcpl_411 : STD_LOGIC;
  SIGNAL and_tmp_27 : STD_LOGIC;
  SIGNAL mux_tmp_150 : STD_LOGIC;
  SIGNAL mux_tmp_151 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL and_dcpl_418 : STD_LOGIC;
  SIGNAL or_tmp_402 : STD_LOGIC;
  SIGNAL and_dcpl_422 : STD_LOGIC;
  SIGNAL mux_tmp_153 : STD_LOGIC;
  SIGNAL and_dcpl_426 : STD_LOGIC;
  SIGNAL mux_tmp_155 : STD_LOGIC;
  SIGNAL mux_tmp_156 : STD_LOGIC;
  SIGNAL and_dcpl_430 : STD_LOGIC;
  SIGNAL mux_tmp_158 : STD_LOGIC;
  SIGNAL mux_tmp_159 : STD_LOGIC;
  SIGNAL mux_tmp_160 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL mux_tmp_162 : STD_LOGIC;
  SIGNAL mux_tmp_163 : STD_LOGIC;
  SIGNAL mux_tmp_164 : STD_LOGIC;
  SIGNAL mux_tmp_165 : STD_LOGIC;
  SIGNAL and_dcpl_437 : STD_LOGIC;
  SIGNAL mux_tmp_167 : STD_LOGIC;
  SIGNAL mux_tmp_168 : STD_LOGIC;
  SIGNAL mux_tmp_169 : STD_LOGIC;
  SIGNAL mux_tmp_170 : STD_LOGIC;
  SIGNAL mux_tmp_171 : STD_LOGIC;
  SIGNAL and_dcpl_441 : STD_LOGIC;
  SIGNAL mux_tmp_173 : STD_LOGIC;
  SIGNAL mux_tmp_174 : STD_LOGIC;
  SIGNAL mux_tmp_175 : STD_LOGIC;
  SIGNAL mux_tmp_176 : STD_LOGIC;
  SIGNAL mux_tmp_177 : STD_LOGIC;
  SIGNAL mux_tmp_178 : STD_LOGIC;
  SIGNAL and_dcpl_444 : STD_LOGIC;
  SIGNAL mux_tmp_180 : STD_LOGIC;
  SIGNAL mux_tmp_181 : STD_LOGIC;
  SIGNAL mux_tmp_182 : STD_LOGIC;
  SIGNAL mux_tmp_183 : STD_LOGIC;
  SIGNAL mux_tmp_184 : STD_LOGIC;
  SIGNAL mux_tmp_185 : STD_LOGIC;
  SIGNAL mux_tmp_186 : STD_LOGIC;
  SIGNAL and_dcpl_447 : STD_LOGIC;
  SIGNAL and_tmp_34 : STD_LOGIC;
  SIGNAL mux_tmp_188 : STD_LOGIC;
  SIGNAL mux_tmp_189 : STD_LOGIC;
  SIGNAL and_dcpl_452 : STD_LOGIC;
  SIGNAL or_tmp_502 : STD_LOGIC;
  SIGNAL and_dcpl_455 : STD_LOGIC;
  SIGNAL mux_tmp_191 : STD_LOGIC;
  SIGNAL and_dcpl_458 : STD_LOGIC;
  SIGNAL mux_tmp_193 : STD_LOGIC;
  SIGNAL mux_tmp_194 : STD_LOGIC;
  SIGNAL and_dcpl_462 : STD_LOGIC;
  SIGNAL mux_tmp_196 : STD_LOGIC;
  SIGNAL mux_tmp_197 : STD_LOGIC;
  SIGNAL mux_tmp_198 : STD_LOGIC;
  SIGNAL and_dcpl_464 : STD_LOGIC;
  SIGNAL mux_tmp_200 : STD_LOGIC;
  SIGNAL mux_tmp_201 : STD_LOGIC;
  SIGNAL mux_tmp_202 : STD_LOGIC;
  SIGNAL mux_tmp_203 : STD_LOGIC;
  SIGNAL and_dcpl_468 : STD_LOGIC;
  SIGNAL mux_tmp_205 : STD_LOGIC;
  SIGNAL mux_tmp_206 : STD_LOGIC;
  SIGNAL mux_tmp_207 : STD_LOGIC;
  SIGNAL mux_tmp_208 : STD_LOGIC;
  SIGNAL mux_tmp_209 : STD_LOGIC;
  SIGNAL and_dcpl_472 : STD_LOGIC;
  SIGNAL mux_tmp_211 : STD_LOGIC;
  SIGNAL mux_tmp_212 : STD_LOGIC;
  SIGNAL mux_tmp_213 : STD_LOGIC;
  SIGNAL mux_tmp_214 : STD_LOGIC;
  SIGNAL mux_tmp_215 : STD_LOGIC;
  SIGNAL mux_tmp_216 : STD_LOGIC;
  SIGNAL and_dcpl_474 : STD_LOGIC;
  SIGNAL mux_tmp_218 : STD_LOGIC;
  SIGNAL mux_tmp_219 : STD_LOGIC;
  SIGNAL mux_tmp_220 : STD_LOGIC;
  SIGNAL mux_tmp_221 : STD_LOGIC;
  SIGNAL mux_tmp_222 : STD_LOGIC;
  SIGNAL mux_tmp_223 : STD_LOGIC;
  SIGNAL mux_tmp_224 : STD_LOGIC;
  SIGNAL and_dcpl_476 : STD_LOGIC;
  SIGNAL and_tmp_41 : STD_LOGIC;
  SIGNAL mux_tmp_226 : STD_LOGIC;
  SIGNAL mux_tmp_227 : STD_LOGIC;
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL or_tmp_602 : STD_LOGIC;
  SIGNAL and_dcpl_484 : STD_LOGIC;
  SIGNAL mux_tmp_229 : STD_LOGIC;
  SIGNAL and_dcpl_488 : STD_LOGIC;
  SIGNAL mux_tmp_231 : STD_LOGIC;
  SIGNAL mux_tmp_232 : STD_LOGIC;
  SIGNAL and_dcpl_491 : STD_LOGIC;
  SIGNAL mux_tmp_234 : STD_LOGIC;
  SIGNAL mux_tmp_235 : STD_LOGIC;
  SIGNAL mux_tmp_236 : STD_LOGIC;
  SIGNAL and_dcpl_493 : STD_LOGIC;
  SIGNAL mux_tmp_238 : STD_LOGIC;
  SIGNAL mux_tmp_239 : STD_LOGIC;
  SIGNAL mux_tmp_240 : STD_LOGIC;
  SIGNAL mux_tmp_241 : STD_LOGIC;
  SIGNAL and_dcpl_496 : STD_LOGIC;
  SIGNAL mux_tmp_243 : STD_LOGIC;
  SIGNAL mux_tmp_244 : STD_LOGIC;
  SIGNAL mux_tmp_245 : STD_LOGIC;
  SIGNAL mux_tmp_246 : STD_LOGIC;
  SIGNAL mux_tmp_247 : STD_LOGIC;
  SIGNAL and_dcpl_499 : STD_LOGIC;
  SIGNAL mux_tmp_249 : STD_LOGIC;
  SIGNAL mux_tmp_250 : STD_LOGIC;
  SIGNAL mux_tmp_251 : STD_LOGIC;
  SIGNAL mux_tmp_252 : STD_LOGIC;
  SIGNAL mux_tmp_253 : STD_LOGIC;
  SIGNAL mux_tmp_254 : STD_LOGIC;
  SIGNAL and_dcpl_501 : STD_LOGIC;
  SIGNAL mux_tmp_256 : STD_LOGIC;
  SIGNAL mux_tmp_257 : STD_LOGIC;
  SIGNAL mux_tmp_258 : STD_LOGIC;
  SIGNAL mux_tmp_259 : STD_LOGIC;
  SIGNAL mux_tmp_260 : STD_LOGIC;
  SIGNAL mux_tmp_261 : STD_LOGIC;
  SIGNAL mux_tmp_262 : STD_LOGIC;
  SIGNAL and_dcpl_503 : STD_LOGIC;
  SIGNAL and_tmp_48 : STD_LOGIC;
  SIGNAL mux_tmp_264 : STD_LOGIC;
  SIGNAL mux_tmp_265 : STD_LOGIC;
  SIGNAL and_dcpl_507 : STD_LOGIC;
  SIGNAL or_tmp_702 : STD_LOGIC;
  SIGNAL and_dcpl_510 : STD_LOGIC;
  SIGNAL mux_tmp_267 : STD_LOGIC;
  SIGNAL and_dcpl_513 : STD_LOGIC;
  SIGNAL mux_tmp_269 : STD_LOGIC;
  SIGNAL mux_tmp_270 : STD_LOGIC;
  SIGNAL and_dcpl_516 : STD_LOGIC;
  SIGNAL mux_tmp_272 : STD_LOGIC;
  SIGNAL mux_tmp_273 : STD_LOGIC;
  SIGNAL mux_tmp_274 : STD_LOGIC;
  SIGNAL and_dcpl_518 : STD_LOGIC;
  SIGNAL mux_tmp_276 : STD_LOGIC;
  SIGNAL mux_tmp_277 : STD_LOGIC;
  SIGNAL mux_tmp_278 : STD_LOGIC;
  SIGNAL mux_tmp_279 : STD_LOGIC;
  SIGNAL and_dcpl_521 : STD_LOGIC;
  SIGNAL mux_tmp_281 : STD_LOGIC;
  SIGNAL mux_tmp_282 : STD_LOGIC;
  SIGNAL mux_tmp_283 : STD_LOGIC;
  SIGNAL mux_tmp_284 : STD_LOGIC;
  SIGNAL mux_tmp_285 : STD_LOGIC;
  SIGNAL and_dcpl_524 : STD_LOGIC;
  SIGNAL mux_tmp_287 : STD_LOGIC;
  SIGNAL mux_tmp_288 : STD_LOGIC;
  SIGNAL mux_tmp_289 : STD_LOGIC;
  SIGNAL mux_tmp_290 : STD_LOGIC;
  SIGNAL mux_tmp_291 : STD_LOGIC;
  SIGNAL mux_tmp_292 : STD_LOGIC;
  SIGNAL and_dcpl_526 : STD_LOGIC;
  SIGNAL mux_tmp_294 : STD_LOGIC;
  SIGNAL mux_tmp_295 : STD_LOGIC;
  SIGNAL mux_tmp_296 : STD_LOGIC;
  SIGNAL mux_tmp_297 : STD_LOGIC;
  SIGNAL mux_tmp_298 : STD_LOGIC;
  SIGNAL mux_tmp_299 : STD_LOGIC;
  SIGNAL mux_tmp_300 : STD_LOGIC;
  SIGNAL and_dcpl_528 : STD_LOGIC;
  SIGNAL and_tmp_55 : STD_LOGIC;
  SIGNAL mux_tmp_302 : STD_LOGIC;
  SIGNAL mux_tmp_303 : STD_LOGIC;
  SIGNAL and_dcpl_532 : STD_LOGIC;
  SIGNAL and_dcpl_533 : STD_LOGIC;
  SIGNAL not_tmp_645 : STD_LOGIC;
  SIGNAL or_tmp_801 : STD_LOGIC;
  SIGNAL and_dcpl_536 : STD_LOGIC;
  SIGNAL mux_tmp_305 : STD_LOGIC;
  SIGNAL and_dcpl_539 : STD_LOGIC;
  SIGNAL mux_tmp_307 : STD_LOGIC;
  SIGNAL mux_tmp_308 : STD_LOGIC;
  SIGNAL and_dcpl_542 : STD_LOGIC;
  SIGNAL mux_tmp_310 : STD_LOGIC;
  SIGNAL mux_tmp_311 : STD_LOGIC;
  SIGNAL mux_tmp_312 : STD_LOGIC;
  SIGNAL and_dcpl_546 : STD_LOGIC;
  SIGNAL mux_tmp_314 : STD_LOGIC;
  SIGNAL mux_tmp_315 : STD_LOGIC;
  SIGNAL mux_tmp_316 : STD_LOGIC;
  SIGNAL mux_tmp_317 : STD_LOGIC;
  SIGNAL and_dcpl_549 : STD_LOGIC;
  SIGNAL mux_tmp_319 : STD_LOGIC;
  SIGNAL mux_tmp_320 : STD_LOGIC;
  SIGNAL mux_tmp_321 : STD_LOGIC;
  SIGNAL mux_tmp_322 : STD_LOGIC;
  SIGNAL mux_tmp_323 : STD_LOGIC;
  SIGNAL and_dcpl_552 : STD_LOGIC;
  SIGNAL mux_tmp_325 : STD_LOGIC;
  SIGNAL mux_tmp_326 : STD_LOGIC;
  SIGNAL mux_tmp_327 : STD_LOGIC;
  SIGNAL mux_tmp_328 : STD_LOGIC;
  SIGNAL mux_tmp_329 : STD_LOGIC;
  SIGNAL mux_tmp_330 : STD_LOGIC;
  SIGNAL and_dcpl_556 : STD_LOGIC;
  SIGNAL mux_tmp_332 : STD_LOGIC;
  SIGNAL mux_tmp_333 : STD_LOGIC;
  SIGNAL mux_tmp_334 : STD_LOGIC;
  SIGNAL mux_tmp_335 : STD_LOGIC;
  SIGNAL mux_tmp_336 : STD_LOGIC;
  SIGNAL mux_tmp_337 : STD_LOGIC;
  SIGNAL mux_tmp_338 : STD_LOGIC;
  SIGNAL and_dcpl_560 : STD_LOGIC;
  SIGNAL or_tmp_897 : STD_LOGIC;
  SIGNAL mux_tmp_340 : STD_LOGIC;
  SIGNAL mux_tmp_341 : STD_LOGIC;
  SIGNAL mux_tmp_342 : STD_LOGIC;
  SIGNAL mux_tmp_343 : STD_LOGIC;
  SIGNAL mux_tmp_344 : STD_LOGIC;
  SIGNAL mux_tmp_345 : STD_LOGIC;
  SIGNAL mux_tmp_346 : STD_LOGIC;
  SIGNAL mux_tmp_347 : STD_LOGIC;
  SIGNAL mux_tmp_348 : STD_LOGIC;
  SIGNAL and_dcpl_566 : STD_LOGIC;
  SIGNAL or_tmp_909 : STD_LOGIC;
  SIGNAL and_dcpl_568 : STD_LOGIC;
  SIGNAL mux_tmp_350 : STD_LOGIC;
  SIGNAL and_dcpl_570 : STD_LOGIC;
  SIGNAL mux_tmp_352 : STD_LOGIC;
  SIGNAL mux_tmp_353 : STD_LOGIC;
  SIGNAL and_dcpl_572 : STD_LOGIC;
  SIGNAL mux_tmp_355 : STD_LOGIC;
  SIGNAL mux_tmp_356 : STD_LOGIC;
  SIGNAL mux_tmp_357 : STD_LOGIC;
  SIGNAL and_dcpl_576 : STD_LOGIC;
  SIGNAL mux_tmp_359 : STD_LOGIC;
  SIGNAL mux_tmp_360 : STD_LOGIC;
  SIGNAL mux_tmp_361 : STD_LOGIC;
  SIGNAL mux_tmp_362 : STD_LOGIC;
  SIGNAL and_dcpl_578 : STD_LOGIC;
  SIGNAL mux_tmp_364 : STD_LOGIC;
  SIGNAL mux_tmp_365 : STD_LOGIC;
  SIGNAL mux_tmp_366 : STD_LOGIC;
  SIGNAL mux_tmp_367 : STD_LOGIC;
  SIGNAL mux_tmp_368 : STD_LOGIC;
  SIGNAL and_dcpl_580 : STD_LOGIC;
  SIGNAL mux_tmp_370 : STD_LOGIC;
  SIGNAL mux_tmp_371 : STD_LOGIC;
  SIGNAL mux_tmp_372 : STD_LOGIC;
  SIGNAL mux_tmp_373 : STD_LOGIC;
  SIGNAL mux_tmp_374 : STD_LOGIC;
  SIGNAL mux_tmp_375 : STD_LOGIC;
  SIGNAL and_dcpl_583 : STD_LOGIC;
  SIGNAL mux_tmp_377 : STD_LOGIC;
  SIGNAL mux_tmp_378 : STD_LOGIC;
  SIGNAL mux_tmp_379 : STD_LOGIC;
  SIGNAL mux_tmp_380 : STD_LOGIC;
  SIGNAL mux_tmp_381 : STD_LOGIC;
  SIGNAL mux_tmp_382 : STD_LOGIC;
  SIGNAL mux_tmp_383 : STD_LOGIC;
  SIGNAL and_dcpl_586 : STD_LOGIC;
  SIGNAL or_tmp_1005 : STD_LOGIC;
  SIGNAL mux_tmp_385 : STD_LOGIC;
  SIGNAL mux_tmp_386 : STD_LOGIC;
  SIGNAL mux_tmp_387 : STD_LOGIC;
  SIGNAL mux_tmp_388 : STD_LOGIC;
  SIGNAL mux_tmp_389 : STD_LOGIC;
  SIGNAL mux_tmp_390 : STD_LOGIC;
  SIGNAL mux_tmp_391 : STD_LOGIC;
  SIGNAL mux_tmp_392 : STD_LOGIC;
  SIGNAL mux_tmp_393 : STD_LOGIC;
  SIGNAL and_dcpl_590 : STD_LOGIC;
  SIGNAL or_tmp_1017 : STD_LOGIC;
  SIGNAL and_dcpl_592 : STD_LOGIC;
  SIGNAL mux_tmp_395 : STD_LOGIC;
  SIGNAL and_dcpl_594 : STD_LOGIC;
  SIGNAL mux_tmp_397 : STD_LOGIC;
  SIGNAL mux_tmp_398 : STD_LOGIC;
  SIGNAL and_dcpl_596 : STD_LOGIC;
  SIGNAL mux_tmp_400 : STD_LOGIC;
  SIGNAL mux_tmp_401 : STD_LOGIC;
  SIGNAL mux_tmp_402 : STD_LOGIC;
  SIGNAL and_dcpl_599 : STD_LOGIC;
  SIGNAL mux_tmp_404 : STD_LOGIC;
  SIGNAL mux_tmp_405 : STD_LOGIC;
  SIGNAL mux_tmp_406 : STD_LOGIC;
  SIGNAL mux_tmp_407 : STD_LOGIC;
  SIGNAL and_dcpl_601 : STD_LOGIC;
  SIGNAL mux_tmp_409 : STD_LOGIC;
  SIGNAL mux_tmp_410 : STD_LOGIC;
  SIGNAL mux_tmp_411 : STD_LOGIC;
  SIGNAL mux_tmp_412 : STD_LOGIC;
  SIGNAL mux_tmp_413 : STD_LOGIC;
  SIGNAL and_dcpl_603 : STD_LOGIC;
  SIGNAL mux_tmp_415 : STD_LOGIC;
  SIGNAL mux_tmp_416 : STD_LOGIC;
  SIGNAL mux_tmp_417 : STD_LOGIC;
  SIGNAL mux_tmp_418 : STD_LOGIC;
  SIGNAL mux_tmp_419 : STD_LOGIC;
  SIGNAL mux_tmp_420 : STD_LOGIC;
  SIGNAL and_dcpl_607 : STD_LOGIC;
  SIGNAL mux_tmp_422 : STD_LOGIC;
  SIGNAL mux_tmp_423 : STD_LOGIC;
  SIGNAL mux_tmp_424 : STD_LOGIC;
  SIGNAL mux_tmp_425 : STD_LOGIC;
  SIGNAL mux_tmp_426 : STD_LOGIC;
  SIGNAL mux_tmp_427 : STD_LOGIC;
  SIGNAL mux_tmp_428 : STD_LOGIC;
  SIGNAL and_dcpl_611 : STD_LOGIC;
  SIGNAL or_tmp_1113 : STD_LOGIC;
  SIGNAL mux_tmp_430 : STD_LOGIC;
  SIGNAL mux_tmp_431 : STD_LOGIC;
  SIGNAL mux_tmp_432 : STD_LOGIC;
  SIGNAL mux_tmp_433 : STD_LOGIC;
  SIGNAL mux_tmp_434 : STD_LOGIC;
  SIGNAL mux_tmp_435 : STD_LOGIC;
  SIGNAL mux_tmp_436 : STD_LOGIC;
  SIGNAL mux_tmp_437 : STD_LOGIC;
  SIGNAL mux_tmp_438 : STD_LOGIC;
  SIGNAL main_stage_0_11 : STD_LOGIC;
  SIGNAL asn_itm_10 : STD_LOGIC;
  SIGNAL result_rem_11cyc_st_9 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_8 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_7 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_6 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_5 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_4 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_3 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_2 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_11 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL asn_itm_11 : STD_LOGIC;
  SIGNAL main_stage_0_12 : STD_LOGIC;
  SIGNAL main_stage_0_3 : STD_LOGIC;
  SIGNAL asn_itm_2 : STD_LOGIC;
  SIGNAL main_stage_0_4 : STD_LOGIC;
  SIGNAL asn_itm_3 : STD_LOGIC;
  SIGNAL main_stage_0_5 : STD_LOGIC;
  SIGNAL asn_itm_4 : STD_LOGIC;
  SIGNAL main_stage_0_6 : STD_LOGIC;
  SIGNAL asn_itm_5 : STD_LOGIC;
  SIGNAL main_stage_0_7 : STD_LOGIC;
  SIGNAL asn_itm_6 : STD_LOGIC;
  SIGNAL main_stage_0_8 : STD_LOGIC;
  SIGNAL asn_itm_7 : STD_LOGIC;
  SIGNAL main_stage_0_9 : STD_LOGIC;
  SIGNAL asn_itm_8 : STD_LOGIC;
  SIGNAL main_stage_0_10 : STD_LOGIC;
  SIGNAL asn_itm_9 : STD_LOGIC;
  SIGNAL main_stage_0_2 : STD_LOGIC;
  SIGNAL asn_itm_1 : STD_LOGIC;
  SIGNAL result_and_1_cse : STD_LOGIC;
  SIGNAL result_and_3_cse : STD_LOGIC;
  SIGNAL result_and_5_cse : STD_LOGIC;
  SIGNAL result_and_7_cse : STD_LOGIC;
  SIGNAL result_and_9_cse : STD_LOGIC;
  SIGNAL result_and_11_cse : STD_LOGIC;
  SIGNAL result_and_13_cse : STD_LOGIC;
  SIGNAL result_and_15_cse : STD_LOGIC;
  SIGNAL result_and_17_cse : STD_LOGIC;
  SIGNAL result_and_19_cse : STD_LOGIC;
  SIGNAL result_and_21_cse : STD_LOGIC;
  SIGNAL or_3_cse : STD_LOGIC;
  SIGNAL or_8_cse : STD_LOGIC;
  SIGNAL or_15_cse : STD_LOGIC;
  SIGNAL or_24_cse : STD_LOGIC;
  SIGNAL or_35_cse : STD_LOGIC;
  SIGNAL or_48_cse : STD_LOGIC;
  SIGNAL or_63_cse : STD_LOGIC;
  SIGNAL or_107_cse : STD_LOGIC;
  SIGNAL or_112_cse : STD_LOGIC;
  SIGNAL or_119_cse : STD_LOGIC;
  SIGNAL or_128_cse : STD_LOGIC;
  SIGNAL or_139_cse : STD_LOGIC;
  SIGNAL or_152_cse : STD_LOGIC;
  SIGNAL or_167_cse : STD_LOGIC;
  SIGNAL or_209_cse : STD_LOGIC;
  SIGNAL or_214_cse : STD_LOGIC;
  SIGNAL or_221_cse : STD_LOGIC;
  SIGNAL or_230_cse : STD_LOGIC;
  SIGNAL or_241_cse : STD_LOGIC;
  SIGNAL or_254_cse : STD_LOGIC;
  SIGNAL or_269_cse : STD_LOGIC;
  SIGNAL or_311_cse : STD_LOGIC;
  SIGNAL or_316_cse : STD_LOGIC;
  SIGNAL or_323_cse : STD_LOGIC;
  SIGNAL or_332_cse : STD_LOGIC;
  SIGNAL or_343_cse : STD_LOGIC;
  SIGNAL or_356_cse : STD_LOGIC;
  SIGNAL or_371_cse : STD_LOGIC;
  SIGNAL nand_144_cse : STD_LOGIC;
  SIGNAL or_413_cse : STD_LOGIC;
  SIGNAL or_418_cse : STD_LOGIC;
  SIGNAL or_425_cse : STD_LOGIC;
  SIGNAL or_434_cse : STD_LOGIC;
  SIGNAL or_445_cse : STD_LOGIC;
  SIGNAL or_458_cse : STD_LOGIC;
  SIGNAL or_473_cse : STD_LOGIC;
  SIGNAL nand_138_cse : STD_LOGIC;
  SIGNAL or_516_cse : STD_LOGIC;
  SIGNAL or_521_cse : STD_LOGIC;
  SIGNAL or_528_cse : STD_LOGIC;
  SIGNAL or_537_cse : STD_LOGIC;
  SIGNAL and_790_cse : STD_LOGIC;
  SIGNAL or_548_cse : STD_LOGIC;
  SIGNAL or_561_cse : STD_LOGIC;
  SIGNAL or_576_cse : STD_LOGIC;
  SIGNAL nand_146_cse : STD_LOGIC;
  SIGNAL or_617_cse : STD_LOGIC;
  SIGNAL or_622_cse : STD_LOGIC;
  SIGNAL or_629_cse : STD_LOGIC;
  SIGNAL or_638_cse : STD_LOGIC;
  SIGNAL or_649_cse : STD_LOGIC;
  SIGNAL or_662_cse : STD_LOGIC;
  SIGNAL or_677_cse : STD_LOGIC;
  SIGNAL or_718_cse : STD_LOGIC;
  SIGNAL nand_112_cse : STD_LOGIC;
  SIGNAL nand_108_cse : STD_LOGIC;
  SIGNAL nand_103_cse : STD_LOGIC;
  SIGNAL nand_97_cse : STD_LOGIC;
  SIGNAL or_763_cse : STD_LOGIC;
  SIGNAL nand_83_cse : STD_LOGIC;
  SIGNAL or_818_cse : STD_LOGIC;
  SIGNAL or_823_cse : STD_LOGIC;
  SIGNAL or_830_cse : STD_LOGIC;
  SIGNAL or_839_cse : STD_LOGIC;
  SIGNAL nand_58_cse : STD_LOGIC;
  SIGNAL or_850_cse : STD_LOGIC;
  SIGNAL nand_55_cse : STD_LOGIC;
  SIGNAL or_863_cse : STD_LOGIC;
  SIGNAL nand_51_cse : STD_LOGIC;
  SIGNAL or_878_cse : STD_LOGIC;
  SIGNAL and_749_cse : STD_LOGIC;
  SIGNAL or_928_cse : STD_LOGIC;
  SIGNAL and_747_cse : STD_LOGIC;
  SIGNAL or_933_cse : STD_LOGIC;
  SIGNAL and_744_cse : STD_LOGIC;
  SIGNAL or_940_cse : STD_LOGIC;
  SIGNAL and_740_cse : STD_LOGIC;
  SIGNAL or_949_cse : STD_LOGIC;
  SIGNAL or_960_cse : STD_LOGIC;
  SIGNAL and_731_cse : STD_LOGIC;
  SIGNAL or_973_cse : STD_LOGIC;
  SIGNAL and_725_cse : STD_LOGIC;
  SIGNAL nand_42_cse : STD_LOGIC;
  SIGNAL or_988_cse : STD_LOGIC;
  SIGNAL or_1037_cse : STD_LOGIC;
  SIGNAL or_1042_cse : STD_LOGIC;
  SIGNAL or_1049_cse : STD_LOGIC;
  SIGNAL or_1058_cse : STD_LOGIC;
  SIGNAL or_1069_cse : STD_LOGIC;
  SIGNAL or_1082_cse : STD_LOGIC;
  SIGNAL or_1097_cse : STD_LOGIC;
  SIGNAL base_buf_sva_mut_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_10 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL return_rsci_d_mx0c0 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c1 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c2 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c3 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c4 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c5 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c6 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c7 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c8 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c9 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c10 : STD_LOGIC;
  SIGNAL result_acc_imod_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_acc_idiv_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL m_and_cse : STD_LOGIC;
  SIGNAL m_and_1_cse : STD_LOGIC;
  SIGNAL m_and_2_cse : STD_LOGIC;
  SIGNAL m_and_3_cse : STD_LOGIC;
  SIGNAL m_and_4_cse : STD_LOGIC;
  SIGNAL m_and_5_cse : STD_LOGIC;
  SIGNAL m_and_6_cse : STD_LOGIC;
  SIGNAL m_and_7_cse : STD_LOGIC;
  SIGNAL m_and_8_cse : STD_LOGIC;
  SIGNAL m_and_9_cse : STD_LOGIC;
  SIGNAL m_and_10_cse : STD_LOGIC;
  SIGNAL m_and_11_cse : STD_LOGIC;
  SIGNAL m_and_12_cse : STD_LOGIC;
  SIGNAL m_and_13_cse : STD_LOGIC;
  SIGNAL m_and_14_cse : STD_LOGIC;
  SIGNAL m_and_15_cse : STD_LOGIC;
  SIGNAL m_and_16_cse : STD_LOGIC;
  SIGNAL m_and_17_cse : STD_LOGIC;
  SIGNAL m_and_18_cse : STD_LOGIC;
  SIGNAL m_and_19_cse : STD_LOGIC;
  SIGNAL m_and_20_cse : STD_LOGIC;
  SIGNAL m_and_21_cse : STD_LOGIC;
  SIGNAL m_and_22_cse : STD_LOGIC;
  SIGNAL m_and_23_cse : STD_LOGIC;
  SIGNAL m_and_24_cse : STD_LOGIC;
  SIGNAL m_and_25_cse : STD_LOGIC;
  SIGNAL m_and_26_cse : STD_LOGIC;
  SIGNAL m_and_27_cse : STD_LOGIC;
  SIGNAL m_and_28_cse : STD_LOGIC;
  SIGNAL m_and_29_cse : STD_LOGIC;
  SIGNAL m_and_30_cse : STD_LOGIC;
  SIGNAL m_and_31_cse : STD_LOGIC;
  SIGNAL m_and_32_cse : STD_LOGIC;
  SIGNAL m_and_33_cse : STD_LOGIC;
  SIGNAL m_and_34_cse : STD_LOGIC;
  SIGNAL m_and_35_cse : STD_LOGIC;
  SIGNAL m_and_36_cse : STD_LOGIC;
  SIGNAL m_and_37_cse : STD_LOGIC;
  SIGNAL m_and_38_cse : STD_LOGIC;
  SIGNAL m_and_39_cse : STD_LOGIC;
  SIGNAL m_and_40_cse : STD_LOGIC;
  SIGNAL m_and_41_cse : STD_LOGIC;
  SIGNAL m_and_42_cse : STD_LOGIC;
  SIGNAL m_and_43_cse : STD_LOGIC;
  SIGNAL m_and_44_cse : STD_LOGIC;
  SIGNAL m_and_45_cse : STD_LOGIC;
  SIGNAL m_and_46_cse : STD_LOGIC;
  SIGNAL m_and_47_cse : STD_LOGIC;
  SIGNAL m_and_48_cse : STD_LOGIC;
  SIGNAL m_and_49_cse : STD_LOGIC;
  SIGNAL m_and_50_cse : STD_LOGIC;
  SIGNAL m_and_51_cse : STD_LOGIC;
  SIGNAL m_and_52_cse : STD_LOGIC;
  SIGNAL m_and_53_cse : STD_LOGIC;
  SIGNAL m_and_54_cse : STD_LOGIC;
  SIGNAL m_and_55_cse : STD_LOGIC;
  SIGNAL m_and_56_cse : STD_LOGIC;
  SIGNAL m_and_57_cse : STD_LOGIC;
  SIGNAL m_and_58_cse : STD_LOGIC;
  SIGNAL m_and_59_cse : STD_LOGIC;
  SIGNAL m_and_60_cse : STD_LOGIC;
  SIGNAL m_and_61_cse : STD_LOGIC;
  SIGNAL m_and_62_cse : STD_LOGIC;
  SIGNAL m_and_63_cse : STD_LOGIC;
  SIGNAL m_and_64_cse : STD_LOGIC;
  SIGNAL m_and_65_cse : STD_LOGIC;
  SIGNAL m_and_66_cse : STD_LOGIC;
  SIGNAL m_and_67_cse : STD_LOGIC;
  SIGNAL m_and_68_cse : STD_LOGIC;
  SIGNAL m_and_69_cse : STD_LOGIC;
  SIGNAL m_and_70_cse : STD_LOGIC;
  SIGNAL m_and_71_cse : STD_LOGIC;
  SIGNAL m_and_72_cse : STD_LOGIC;
  SIGNAL m_and_73_cse : STD_LOGIC;
  SIGNAL m_and_74_cse : STD_LOGIC;
  SIGNAL m_and_75_cse : STD_LOGIC;
  SIGNAL m_and_76_cse : STD_LOGIC;
  SIGNAL m_and_77_cse : STD_LOGIC;
  SIGNAL m_and_78_cse : STD_LOGIC;
  SIGNAL m_and_79_cse : STD_LOGIC;
  SIGNAL m_and_80_cse : STD_LOGIC;
  SIGNAL m_and_81_cse : STD_LOGIC;
  SIGNAL m_and_82_cse : STD_LOGIC;
  SIGNAL m_and_83_cse : STD_LOGIC;
  SIGNAL m_and_84_cse : STD_LOGIC;
  SIGNAL m_and_85_cse : STD_LOGIC;
  SIGNAL m_and_86_cse : STD_LOGIC;
  SIGNAL m_and_87_cse : STD_LOGIC;
  SIGNAL m_and_88_cse : STD_LOGIC;
  SIGNAL m_and_89_cse : STD_LOGIC;
  SIGNAL m_and_90_cse : STD_LOGIC;
  SIGNAL m_and_91_cse : STD_LOGIC;
  SIGNAL m_and_92_cse : STD_LOGIC;
  SIGNAL m_and_93_cse : STD_LOGIC;
  SIGNAL m_and_94_cse : STD_LOGIC;
  SIGNAL m_and_95_cse : STD_LOGIC;
  SIGNAL m_and_96_cse : STD_LOGIC;
  SIGNAL m_and_97_cse : STD_LOGIC;
  SIGNAL m_and_98_cse : STD_LOGIC;

  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL nor_691_nl : STD_LOGIC;
  SIGNAL nor_690_nl : STD_LOGIC;
  SIGNAL or_10_nl : STD_LOGIC;
  SIGNAL mux_2_nl : STD_LOGIC;
  SIGNAL nor_689_nl : STD_LOGIC;
  SIGNAL nor_687_nl : STD_LOGIC;
  SIGNAL or_17_nl : STD_LOGIC;
  SIGNAL nor_688_nl : STD_LOGIC;
  SIGNAL mux_5_nl : STD_LOGIC;
  SIGNAL nor_686_nl : STD_LOGIC;
  SIGNAL nor_683_nl : STD_LOGIC;
  SIGNAL or_26_nl : STD_LOGIC;
  SIGNAL nor_684_nl : STD_LOGIC;
  SIGNAL nor_685_nl : STD_LOGIC;
  SIGNAL mux_9_nl : STD_LOGIC;
  SIGNAL nor_682_nl : STD_LOGIC;
  SIGNAL nor_678_nl : STD_LOGIC;
  SIGNAL or_37_nl : STD_LOGIC;
  SIGNAL nor_679_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL mux_14_nl : STD_LOGIC;
  SIGNAL nor_677_nl : STD_LOGIC;
  SIGNAL nor_672_nl : STD_LOGIC;
  SIGNAL or_50_nl : STD_LOGIC;
  SIGNAL nor_673_nl : STD_LOGIC;
  SIGNAL nor_674_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL nor_676_nl : STD_LOGIC;
  SIGNAL mux_20_nl : STD_LOGIC;
  SIGNAL nor_671_nl : STD_LOGIC;
  SIGNAL nor_665_nl : STD_LOGIC;
  SIGNAL or_65_nl : STD_LOGIC;
  SIGNAL nor_666_nl : STD_LOGIC;
  SIGNAL nor_667_nl : STD_LOGIC;
  SIGNAL nor_668_nl : STD_LOGIC;
  SIGNAL nor_669_nl : STD_LOGIC;
  SIGNAL nor_670_nl : STD_LOGIC;
  SIGNAL mux_27_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL nor_656_nl : STD_LOGIC;
  SIGNAL or_82_nl : STD_LOGIC;
  SIGNAL or_80_nl : STD_LOGIC;
  SIGNAL nor_657_nl : STD_LOGIC;
  SIGNAL nor_658_nl : STD_LOGIC;
  SIGNAL nor_659_nl : STD_LOGIC;
  SIGNAL nor_660_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL nor_662_nl : STD_LOGIC;
  SIGNAL mux_35_nl : STD_LOGIC;
  SIGNAL nor_663_nl : STD_LOGIC;
  SIGNAL nor_654_nl : STD_LOGIC;
  SIGNAL nor_655_nl : STD_LOGIC;
  SIGNAL mux_38_nl : STD_LOGIC;
  SIGNAL nor_653_nl : STD_LOGIC;
  SIGNAL nor_652_nl : STD_LOGIC;
  SIGNAL or_114_nl : STD_LOGIC;
  SIGNAL mux_40_nl : STD_LOGIC;
  SIGNAL nor_651_nl : STD_LOGIC;
  SIGNAL nor_649_nl : STD_LOGIC;
  SIGNAL or_121_nl : STD_LOGIC;
  SIGNAL nor_650_nl : STD_LOGIC;
  SIGNAL mux_43_nl : STD_LOGIC;
  SIGNAL nor_648_nl : STD_LOGIC;
  SIGNAL nor_645_nl : STD_LOGIC;
  SIGNAL or_130_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL nor_647_nl : STD_LOGIC;
  SIGNAL mux_47_nl : STD_LOGIC;
  SIGNAL nor_644_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL or_141_nl : STD_LOGIC;
  SIGNAL nor_641_nl : STD_LOGIC;
  SIGNAL nor_642_nl : STD_LOGIC;
  SIGNAL nor_643_nl : STD_LOGIC;
  SIGNAL mux_52_nl : STD_LOGIC;
  SIGNAL nor_639_nl : STD_LOGIC;
  SIGNAL nor_634_nl : STD_LOGIC;
  SIGNAL or_154_nl : STD_LOGIC;
  SIGNAL nor_635_nl : STD_LOGIC;
  SIGNAL nor_636_nl : STD_LOGIC;
  SIGNAL nor_637_nl : STD_LOGIC;
  SIGNAL nor_638_nl : STD_LOGIC;
  SIGNAL mux_58_nl : STD_LOGIC;
  SIGNAL nor_633_nl : STD_LOGIC;
  SIGNAL nor_627_nl : STD_LOGIC;
  SIGNAL or_169_nl : STD_LOGIC;
  SIGNAL nor_628_nl : STD_LOGIC;
  SIGNAL nor_629_nl : STD_LOGIC;
  SIGNAL nor_630_nl : STD_LOGIC;
  SIGNAL nor_631_nl : STD_LOGIC;
  SIGNAL nor_632_nl : STD_LOGIC;
  SIGNAL mux_65_nl : STD_LOGIC;
  SIGNAL nor_626_nl : STD_LOGIC;
  SIGNAL nor_618_nl : STD_LOGIC;
  SIGNAL or_186_nl : STD_LOGIC;
  SIGNAL or_184_nl : STD_LOGIC;
  SIGNAL nor_619_nl : STD_LOGIC;
  SIGNAL nor_620_nl : STD_LOGIC;
  SIGNAL nor_621_nl : STD_LOGIC;
  SIGNAL nor_622_nl : STD_LOGIC;
  SIGNAL nor_623_nl : STD_LOGIC;
  SIGNAL nor_624_nl : STD_LOGIC;
  SIGNAL mux_73_nl : STD_LOGIC;
  SIGNAL nor_625_nl : STD_LOGIC;
  SIGNAL nor_617_nl : STD_LOGIC;
  SIGNAL and_797_nl : STD_LOGIC;
  SIGNAL or_195_nl : STD_LOGIC;
  SIGNAL mux_76_nl : STD_LOGIC;
  SIGNAL nor_616_nl : STD_LOGIC;
  SIGNAL nor_615_nl : STD_LOGIC;
  SIGNAL or_216_nl : STD_LOGIC;
  SIGNAL mux_78_nl : STD_LOGIC;
  SIGNAL nor_614_nl : STD_LOGIC;
  SIGNAL nor_612_nl : STD_LOGIC;
  SIGNAL or_223_nl : STD_LOGIC;
  SIGNAL nor_613_nl : STD_LOGIC;
  SIGNAL mux_81_nl : STD_LOGIC;
  SIGNAL nor_611_nl : STD_LOGIC;
  SIGNAL nor_608_nl : STD_LOGIC;
  SIGNAL or_232_nl : STD_LOGIC;
  SIGNAL nor_609_nl : STD_LOGIC;
  SIGNAL nor_610_nl : STD_LOGIC;
  SIGNAL mux_85_nl : STD_LOGIC;
  SIGNAL nor_607_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL or_243_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL nor_605_nl : STD_LOGIC;
  SIGNAL nor_606_nl : STD_LOGIC;
  SIGNAL mux_90_nl : STD_LOGIC;
  SIGNAL nor_602_nl : STD_LOGIC;
  SIGNAL nor_597_nl : STD_LOGIC;
  SIGNAL or_256_nl : STD_LOGIC;
  SIGNAL nor_598_nl : STD_LOGIC;
  SIGNAL nor_599_nl : STD_LOGIC;
  SIGNAL nor_600_nl : STD_LOGIC;
  SIGNAL nor_601_nl : STD_LOGIC;
  SIGNAL mux_96_nl : STD_LOGIC;
  SIGNAL nor_596_nl : STD_LOGIC;
  SIGNAL nor_590_nl : STD_LOGIC;
  SIGNAL or_271_nl : STD_LOGIC;
  SIGNAL nor_591_nl : STD_LOGIC;
  SIGNAL nor_592_nl : STD_LOGIC;
  SIGNAL nor_593_nl : STD_LOGIC;
  SIGNAL nor_594_nl : STD_LOGIC;
  SIGNAL nor_595_nl : STD_LOGIC;
  SIGNAL mux_103_nl : STD_LOGIC;
  SIGNAL nor_589_nl : STD_LOGIC;
  SIGNAL nor_581_nl : STD_LOGIC;
  SIGNAL or_288_nl : STD_LOGIC;
  SIGNAL or_286_nl : STD_LOGIC;
  SIGNAL nor_582_nl : STD_LOGIC;
  SIGNAL nor_583_nl : STD_LOGIC;
  SIGNAL nor_584_nl : STD_LOGIC;
  SIGNAL nor_585_nl : STD_LOGIC;
  SIGNAL nor_586_nl : STD_LOGIC;
  SIGNAL nor_587_nl : STD_LOGIC;
  SIGNAL mux_111_nl : STD_LOGIC;
  SIGNAL nor_588_nl : STD_LOGIC;
  SIGNAL nor_579_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL mux_114_nl : STD_LOGIC;
  SIGNAL nor_578_nl : STD_LOGIC;
  SIGNAL nor_577_nl : STD_LOGIC;
  SIGNAL or_318_nl : STD_LOGIC;
  SIGNAL mux_116_nl : STD_LOGIC;
  SIGNAL nor_576_nl : STD_LOGIC;
  SIGNAL nor_574_nl : STD_LOGIC;
  SIGNAL or_325_nl : STD_LOGIC;
  SIGNAL nor_575_nl : STD_LOGIC;
  SIGNAL mux_119_nl : STD_LOGIC;
  SIGNAL nor_573_nl : STD_LOGIC;
  SIGNAL nor_570_nl : STD_LOGIC;
  SIGNAL or_334_nl : STD_LOGIC;
  SIGNAL nor_571_nl : STD_LOGIC;
  SIGNAL nor_572_nl : STD_LOGIC;
  SIGNAL mux_123_nl : STD_LOGIC;
  SIGNAL nor_569_nl : STD_LOGIC;
  SIGNAL nor_565_nl : STD_LOGIC;
  SIGNAL or_345_nl : STD_LOGIC;
  SIGNAL nor_566_nl : STD_LOGIC;
  SIGNAL nor_567_nl : STD_LOGIC;
  SIGNAL nor_568_nl : STD_LOGIC;
  SIGNAL mux_128_nl : STD_LOGIC;
  SIGNAL nor_564_nl : STD_LOGIC;
  SIGNAL nor_559_nl : STD_LOGIC;
  SIGNAL or_358_nl : STD_LOGIC;
  SIGNAL nor_560_nl : STD_LOGIC;
  SIGNAL nor_561_nl : STD_LOGIC;
  SIGNAL nor_562_nl : STD_LOGIC;
  SIGNAL nor_563_nl : STD_LOGIC;
  SIGNAL mux_134_nl : STD_LOGIC;
  SIGNAL nor_558_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL or_373_nl : STD_LOGIC;
  SIGNAL nor_553_nl : STD_LOGIC;
  SIGNAL nor_554_nl : STD_LOGIC;
  SIGNAL nor_555_nl : STD_LOGIC;
  SIGNAL nor_556_nl : STD_LOGIC;
  SIGNAL nor_557_nl : STD_LOGIC;
  SIGNAL mux_141_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL nor_543_nl : STD_LOGIC;
  SIGNAL or_390_nl : STD_LOGIC;
  SIGNAL or_388_nl : STD_LOGIC;
  SIGNAL nor_544_nl : STD_LOGIC;
  SIGNAL nor_545_nl : STD_LOGIC;
  SIGNAL nor_546_nl : STD_LOGIC;
  SIGNAL nor_547_nl : STD_LOGIC;
  SIGNAL nor_548_nl : STD_LOGIC;
  SIGNAL nor_549_nl : STD_LOGIC;
  SIGNAL mux_149_nl : STD_LOGIC;
  SIGNAL nor_550_nl : STD_LOGIC;
  SIGNAL nor_542_nl : STD_LOGIC;
  SIGNAL and_796_nl : STD_LOGIC;
  SIGNAL or_399_nl : STD_LOGIC;
  SIGNAL mux_152_nl : STD_LOGIC;
  SIGNAL and_795_nl : STD_LOGIC;
  SIGNAL nor_541_nl : STD_LOGIC;
  SIGNAL or_420_nl : STD_LOGIC;
  SIGNAL mux_154_nl : STD_LOGIC;
  SIGNAL and_794_nl : STD_LOGIC;
  SIGNAL nor_539_nl : STD_LOGIC;
  SIGNAL or_427_nl : STD_LOGIC;
  SIGNAL nor_540_nl : STD_LOGIC;
  SIGNAL mux_157_nl : STD_LOGIC;
  SIGNAL and_793_nl : STD_LOGIC;
  SIGNAL nor_536_nl : STD_LOGIC;
  SIGNAL or_436_nl : STD_LOGIC;
  SIGNAL nor_537_nl : STD_LOGIC;
  SIGNAL nor_538_nl : STD_LOGIC;
  SIGNAL mux_161_nl : STD_LOGIC;
  SIGNAL and_792_nl : STD_LOGIC;
  SIGNAL nor_532_nl : STD_LOGIC;
  SIGNAL or_447_nl : STD_LOGIC;
  SIGNAL nor_533_nl : STD_LOGIC;
  SIGNAL nor_534_nl : STD_LOGIC;
  SIGNAL nor_535_nl : STD_LOGIC;
  SIGNAL mux_166_nl : STD_LOGIC;
  SIGNAL and_791_nl : STD_LOGIC;
  SIGNAL nor_527_nl : STD_LOGIC;
  SIGNAL or_460_nl : STD_LOGIC;
  SIGNAL nor_528_nl : STD_LOGIC;
  SIGNAL nor_529_nl : STD_LOGIC;
  SIGNAL nor_530_nl : STD_LOGIC;
  SIGNAL nor_531_nl : STD_LOGIC;
  SIGNAL mux_172_nl : STD_LOGIC;
  SIGNAL and_789_nl : STD_LOGIC;
  SIGNAL nor_522_nl : STD_LOGIC;
  SIGNAL or_475_nl : STD_LOGIC;
  SIGNAL and_788_nl : STD_LOGIC;
  SIGNAL nor_523_nl : STD_LOGIC;
  SIGNAL nor_524_nl : STD_LOGIC;
  SIGNAL nor_525_nl : STD_LOGIC;
  SIGNAL nor_526_nl : STD_LOGIC;
  SIGNAL mux_179_nl : STD_LOGIC;
  SIGNAL and_787_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL or_492_nl : STD_LOGIC;
  SIGNAL or_490_nl : STD_LOGIC;
  SIGNAL nor_517_nl : STD_LOGIC;
  SIGNAL and_785_nl : STD_LOGIC;
  SIGNAL nor_518_nl : STD_LOGIC;
  SIGNAL nor_519_nl : STD_LOGIC;
  SIGNAL nor_520_nl : STD_LOGIC;
  SIGNAL nor_521_nl : STD_LOGIC;
  SIGNAL mux_187_nl : STD_LOGIC;
  SIGNAL and_786_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL or_501_nl : STD_LOGIC;
  SIGNAL mux_190_nl : STD_LOGIC;
  SIGNAL and_784_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL or_523_nl : STD_LOGIC;
  SIGNAL mux_192_nl : STD_LOGIC;
  SIGNAL and_783_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL or_530_nl : STD_LOGIC;
  SIGNAL nor_512_nl : STD_LOGIC;
  SIGNAL mux_195_nl : STD_LOGIC;
  SIGNAL and_782_nl : STD_LOGIC;
  SIGNAL nor_508_nl : STD_LOGIC;
  SIGNAL or_539_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL mux_199_nl : STD_LOGIC;
  SIGNAL and_781_nl : STD_LOGIC;
  SIGNAL nor_504_nl : STD_LOGIC;
  SIGNAL or_550_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL nor_506_nl : STD_LOGIC;
  SIGNAL nor_507_nl : STD_LOGIC;
  SIGNAL mux_204_nl : STD_LOGIC;
  SIGNAL and_780_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL or_563_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL nor_501_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL nor_503_nl : STD_LOGIC;
  SIGNAL mux_210_nl : STD_LOGIC;
  SIGNAL and_778_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL or_578_nl : STD_LOGIC;
  SIGNAL and_777_nl : STD_LOGIC;
  SIGNAL nor_495_nl : STD_LOGIC;
  SIGNAL nor_496_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL mux_217_nl : STD_LOGIC;
  SIGNAL and_776_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL or_595_nl : STD_LOGIC;
  SIGNAL or_593_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL and_774_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL nor_491_nl : STD_LOGIC;
  SIGNAL nor_492_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL mux_225_nl : STD_LOGIC;
  SIGNAL and_775_nl : STD_LOGIC;
  SIGNAL nor_487_nl : STD_LOGIC;
  SIGNAL and_773_nl : STD_LOGIC;
  SIGNAL or_604_nl : STD_LOGIC;
  SIGNAL mux_228_nl : STD_LOGIC;
  SIGNAL and_772_nl : STD_LOGIC;
  SIGNAL nor_486_nl : STD_LOGIC;
  SIGNAL or_624_nl : STD_LOGIC;
  SIGNAL mux_230_nl : STD_LOGIC;
  SIGNAL and_771_nl : STD_LOGIC;
  SIGNAL nor_484_nl : STD_LOGIC;
  SIGNAL or_631_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL mux_233_nl : STD_LOGIC;
  SIGNAL and_770_nl : STD_LOGIC;
  SIGNAL nor_481_nl : STD_LOGIC;
  SIGNAL or_640_nl : STD_LOGIC;
  SIGNAL nor_482_nl : STD_LOGIC;
  SIGNAL nor_483_nl : STD_LOGIC;
  SIGNAL mux_237_nl : STD_LOGIC;
  SIGNAL and_769_nl : STD_LOGIC;
  SIGNAL nor_477_nl : STD_LOGIC;
  SIGNAL or_651_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL nor_479_nl : STD_LOGIC;
  SIGNAL nor_480_nl : STD_LOGIC;
  SIGNAL mux_242_nl : STD_LOGIC;
  SIGNAL and_768_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL or_664_nl : STD_LOGIC;
  SIGNAL nor_473_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL nor_476_nl : STD_LOGIC;
  SIGNAL mux_248_nl : STD_LOGIC;
  SIGNAL and_766_nl : STD_LOGIC;
  SIGNAL nor_467_nl : STD_LOGIC;
  SIGNAL or_679_nl : STD_LOGIC;
  SIGNAL and_765_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL nor_471_nl : STD_LOGIC;
  SIGNAL mux_255_nl : STD_LOGIC;
  SIGNAL and_764_nl : STD_LOGIC;
  SIGNAL nor_461_nl : STD_LOGIC;
  SIGNAL or_696_nl : STD_LOGIC;
  SIGNAL or_694_nl : STD_LOGIC;
  SIGNAL nor_462_nl : STD_LOGIC;
  SIGNAL and_762_nl : STD_LOGIC;
  SIGNAL nor_463_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL nor_465_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL mux_263_nl : STD_LOGIC;
  SIGNAL and_763_nl : STD_LOGIC;
  SIGNAL nor_459_nl : STD_LOGIC;
  SIGNAL nor_460_nl : STD_LOGIC;
  SIGNAL or_705_nl : STD_LOGIC;
  SIGNAL mux_266_nl : STD_LOGIC;
  SIGNAL and_761_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL nand_153_nl : STD_LOGIC;
  SIGNAL mux_268_nl : STD_LOGIC;
  SIGNAL and_760_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL nand_152_nl : STD_LOGIC;
  SIGNAL nor_457_nl : STD_LOGIC;
  SIGNAL mux_271_nl : STD_LOGIC;
  SIGNAL and_759_nl : STD_LOGIC;
  SIGNAL nor_453_nl : STD_LOGIC;
  SIGNAL nand_151_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL mux_275_nl : STD_LOGIC;
  SIGNAL and_758_nl : STD_LOGIC;
  SIGNAL nor_449_nl : STD_LOGIC;
  SIGNAL nand_96_nl : STD_LOGIC;
  SIGNAL nor_450_nl : STD_LOGIC;
  SIGNAL nor_451_nl : STD_LOGIC;
  SIGNAL nor_452_nl : STD_LOGIC;
  SIGNAL mux_280_nl : STD_LOGIC;
  SIGNAL and_757_nl : STD_LOGIC;
  SIGNAL nor_444_nl : STD_LOGIC;
  SIGNAL nand_150_nl : STD_LOGIC;
  SIGNAL nor_445_nl : STD_LOGIC;
  SIGNAL nor_446_nl : STD_LOGIC;
  SIGNAL nor_447_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL mux_286_nl : STD_LOGIC;
  SIGNAL and_755_nl : STD_LOGIC;
  SIGNAL nor_439_nl : STD_LOGIC;
  SIGNAL nand_149_nl : STD_LOGIC;
  SIGNAL and_754_nl : STD_LOGIC;
  SIGNAL nor_440_nl : STD_LOGIC;
  SIGNAL nor_441_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL nor_443_nl : STD_LOGIC;
  SIGNAL mux_293_nl : STD_LOGIC;
  SIGNAL and_753_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL nand_72_nl : STD_LOGIC;
  SIGNAL nand_73_nl : STD_LOGIC;
  SIGNAL nor_434_nl : STD_LOGIC;
  SIGNAL and_751_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL nor_436_nl : STD_LOGIC;
  SIGNAL nor_437_nl : STD_LOGIC;
  SIGNAL nor_438_nl : STD_LOGIC;
  SIGNAL mux_301_nl : STD_LOGIC;
  SIGNAL and_752_nl : STD_LOGIC;
  SIGNAL nor_432_nl : STD_LOGIC;
  SIGNAL and_750_nl : STD_LOGIC;
  SIGNAL mux_304_nl : STD_LOGIC;
  SIGNAL nor_431_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL or_825_nl : STD_LOGIC;
  SIGNAL mux_306_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL nor_428_nl : STD_LOGIC;
  SIGNAL or_832_nl : STD_LOGIC;
  SIGNAL and_748_nl : STD_LOGIC;
  SIGNAL mux_309_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL nor_426_nl : STD_LOGIC;
  SIGNAL or_841_nl : STD_LOGIC;
  SIGNAL and_745_nl : STD_LOGIC;
  SIGNAL and_746_nl : STD_LOGIC;
  SIGNAL mux_313_nl : STD_LOGIC;
  SIGNAL nor_425_nl : STD_LOGIC;
  SIGNAL nor_424_nl : STD_LOGIC;
  SIGNAL or_852_nl : STD_LOGIC;
  SIGNAL and_741_nl : STD_LOGIC;
  SIGNAL and_742_nl : STD_LOGIC;
  SIGNAL and_743_nl : STD_LOGIC;
  SIGNAL mux_318_nl : STD_LOGIC;
  SIGNAL nor_423_nl : STD_LOGIC;
  SIGNAL nor_422_nl : STD_LOGIC;
  SIGNAL or_865_nl : STD_LOGIC;
  SIGNAL and_736_nl : STD_LOGIC;
  SIGNAL and_737_nl : STD_LOGIC;
  SIGNAL and_738_nl : STD_LOGIC;
  SIGNAL and_739_nl : STD_LOGIC;
  SIGNAL mux_324_nl : STD_LOGIC;
  SIGNAL nor_421_nl : STD_LOGIC;
  SIGNAL nor_419_nl : STD_LOGIC;
  SIGNAL or_880_nl : STD_LOGIC;
  SIGNAL nor_420_nl : STD_LOGIC;
  SIGNAL and_732_nl : STD_LOGIC;
  SIGNAL and_733_nl : STD_LOGIC;
  SIGNAL and_734_nl : STD_LOGIC;
  SIGNAL and_735_nl : STD_LOGIC;
  SIGNAL mux_331_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL nor_415_nl : STD_LOGIC;
  SIGNAL or_897_nl : STD_LOGIC;
  SIGNAL or_895_nl : STD_LOGIC;
  SIGNAL and_726_nl : STD_LOGIC;
  SIGNAL nor_416_nl : STD_LOGIC;
  SIGNAL and_727_nl : STD_LOGIC;
  SIGNAL and_728_nl : STD_LOGIC;
  SIGNAL and_729_nl : STD_LOGIC;
  SIGNAL and_730_nl : STD_LOGIC;
  SIGNAL mux_339_nl : STD_LOGIC;
  SIGNAL nor_417_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL or_914_nl : STD_LOGIC;
  SIGNAL nor_408_nl : STD_LOGIC;
  SIGNAL or_913_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL or_912_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL or_911_nl : STD_LOGIC;
  SIGNAL nor_411_nl : STD_LOGIC;
  SIGNAL or_910_nl : STD_LOGIC;
  SIGNAL nor_412_nl : STD_LOGIC;
  SIGNAL or_909_nl : STD_LOGIC;
  SIGNAL nor_413_nl : STD_LOGIC;
  SIGNAL or_908_nl : STD_LOGIC;
  SIGNAL and_724_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL mux_349_nl : STD_LOGIC;
  SIGNAL nor_406_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL or_935_nl : STD_LOGIC;
  SIGNAL mux_351_nl : STD_LOGIC;
  SIGNAL nor_404_nl : STD_LOGIC;
  SIGNAL nor_403_nl : STD_LOGIC;
  SIGNAL or_942_nl : STD_LOGIC;
  SIGNAL and_722_nl : STD_LOGIC;
  SIGNAL mux_354_nl : STD_LOGIC;
  SIGNAL nor_402_nl : STD_LOGIC;
  SIGNAL nor_401_nl : STD_LOGIC;
  SIGNAL or_951_nl : STD_LOGIC;
  SIGNAL and_719_nl : STD_LOGIC;
  SIGNAL and_720_nl : STD_LOGIC;
  SIGNAL mux_358_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL nor_399_nl : STD_LOGIC;
  SIGNAL or_962_nl : STD_LOGIC;
  SIGNAL and_715_nl : STD_LOGIC;
  SIGNAL and_716_nl : STD_LOGIC;
  SIGNAL and_717_nl : STD_LOGIC;
  SIGNAL mux_363_nl : STD_LOGIC;
  SIGNAL nor_398_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL or_975_nl : STD_LOGIC;
  SIGNAL and_710_nl : STD_LOGIC;
  SIGNAL and_711_nl : STD_LOGIC;
  SIGNAL and_712_nl : STD_LOGIC;
  SIGNAL and_713_nl : STD_LOGIC;
  SIGNAL mux_369_nl : STD_LOGIC;
  SIGNAL nor_396_nl : STD_LOGIC;
  SIGNAL nor_394_nl : STD_LOGIC;
  SIGNAL or_990_nl : STD_LOGIC;
  SIGNAL nor_395_nl : STD_LOGIC;
  SIGNAL and_706_nl : STD_LOGIC;
  SIGNAL and_707_nl : STD_LOGIC;
  SIGNAL and_708_nl : STD_LOGIC;
  SIGNAL and_709_nl : STD_LOGIC;
  SIGNAL mux_376_nl : STD_LOGIC;
  SIGNAL nor_393_nl : STD_LOGIC;
  SIGNAL nor_390_nl : STD_LOGIC;
  SIGNAL or_1007_nl : STD_LOGIC;
  SIGNAL or_1005_nl : STD_LOGIC;
  SIGNAL and_700_nl : STD_LOGIC;
  SIGNAL nor_391_nl : STD_LOGIC;
  SIGNAL and_701_nl : STD_LOGIC;
  SIGNAL and_702_nl : STD_LOGIC;
  SIGNAL and_703_nl : STD_LOGIC;
  SIGNAL and_704_nl : STD_LOGIC;
  SIGNAL mux_384_nl : STD_LOGIC;
  SIGNAL nor_392_nl : STD_LOGIC;
  SIGNAL nor_383_nl : STD_LOGIC;
  SIGNAL or_1024_nl : STD_LOGIC;
  SIGNAL nor_384_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL nor_385_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL or_1021_nl : STD_LOGIC;
  SIGNAL nor_387_nl : STD_LOGIC;
  SIGNAL or_1020_nl : STD_LOGIC;
  SIGNAL nor_388_nl : STD_LOGIC;
  SIGNAL or_1019_nl : STD_LOGIC;
  SIGNAL nor_389_nl : STD_LOGIC;
  SIGNAL or_1018_nl : STD_LOGIC;
  SIGNAL and_697_nl : STD_LOGIC;
  SIGNAL and_698_nl : STD_LOGIC;
  SIGNAL or_1016_nl : STD_LOGIC;
  SIGNAL mux_394_nl : STD_LOGIC;
  SIGNAL nor_382_nl : STD_LOGIC;
  SIGNAL nor_381_nl : STD_LOGIC;
  SIGNAL or_1044_nl : STD_LOGIC;
  SIGNAL mux_396_nl : STD_LOGIC;
  SIGNAL nor_380_nl : STD_LOGIC;
  SIGNAL nor_379_nl : STD_LOGIC;
  SIGNAL or_1051_nl : STD_LOGIC;
  SIGNAL and_695_nl : STD_LOGIC;
  SIGNAL mux_399_nl : STD_LOGIC;
  SIGNAL nor_378_nl : STD_LOGIC;
  SIGNAL nor_377_nl : STD_LOGIC;
  SIGNAL or_1060_nl : STD_LOGIC;
  SIGNAL and_692_nl : STD_LOGIC;
  SIGNAL and_693_nl : STD_LOGIC;
  SIGNAL mux_403_nl : STD_LOGIC;
  SIGNAL nor_376_nl : STD_LOGIC;
  SIGNAL nor_375_nl : STD_LOGIC;
  SIGNAL or_1071_nl : STD_LOGIC;
  SIGNAL and_688_nl : STD_LOGIC;
  SIGNAL and_689_nl : STD_LOGIC;
  SIGNAL and_690_nl : STD_LOGIC;
  SIGNAL mux_408_nl : STD_LOGIC;
  SIGNAL nor_374_nl : STD_LOGIC;
  SIGNAL nor_373_nl : STD_LOGIC;
  SIGNAL or_1084_nl : STD_LOGIC;
  SIGNAL and_683_nl : STD_LOGIC;
  SIGNAL and_684_nl : STD_LOGIC;
  SIGNAL and_685_nl : STD_LOGIC;
  SIGNAL and_686_nl : STD_LOGIC;
  SIGNAL mux_414_nl : STD_LOGIC;
  SIGNAL nor_372_nl : STD_LOGIC;
  SIGNAL nor_370_nl : STD_LOGIC;
  SIGNAL or_1099_nl : STD_LOGIC;
  SIGNAL nor_371_nl : STD_LOGIC;
  SIGNAL and_679_nl : STD_LOGIC;
  SIGNAL and_680_nl : STD_LOGIC;
  SIGNAL and_681_nl : STD_LOGIC;
  SIGNAL and_682_nl : STD_LOGIC;
  SIGNAL mux_421_nl : STD_LOGIC;
  SIGNAL nor_369_nl : STD_LOGIC;
  SIGNAL nor_366_nl : STD_LOGIC;
  SIGNAL or_1116_nl : STD_LOGIC;
  SIGNAL or_1114_nl : STD_LOGIC;
  SIGNAL and_673_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL and_674_nl : STD_LOGIC;
  SIGNAL and_675_nl : STD_LOGIC;
  SIGNAL and_676_nl : STD_LOGIC;
  SIGNAL and_677_nl : STD_LOGIC;
  SIGNAL mux_429_nl : STD_LOGIC;
  SIGNAL nor_368_nl : STD_LOGIC;
  SIGNAL nor_358_nl : STD_LOGIC;
  SIGNAL or_1133_nl : STD_LOGIC;
  SIGNAL nor_359_nl : STD_LOGIC;
  SIGNAL or_1132_nl : STD_LOGIC;
  SIGNAL nor_360_nl : STD_LOGIC;
  SIGNAL or_1131_nl : STD_LOGIC;
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL or_1130_nl : STD_LOGIC;
  SIGNAL nor_362_nl : STD_LOGIC;
  SIGNAL or_1129_nl : STD_LOGIC;
  SIGNAL nor_363_nl : STD_LOGIC;
  SIGNAL or_1128_nl : STD_LOGIC;
  SIGNAL nor_364_nl : STD_LOGIC;
  SIGNAL or_1127_nl : STD_LOGIC;
  SIGNAL and_671_nl : STD_LOGIC;
  SIGNAL nor_365_nl : STD_LOGIC;
  SIGNAL base_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL m_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL return_rsci_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL ccs_ccore_start_rsci_dat : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat_1 : STD_LOGIC_VECTOR (0 DOWNTO 0);

  SIGNAL result_rem_12_cmp_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_1_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_2_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_3_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_4_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_5_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_6_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_7_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_8_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_9_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_10_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_v_64_10_2(input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(9 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_11_2(input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  base_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 1,
      width => 64
      )
    PORT MAP(
      dat => base_rsci_dat,
      idat => base_rsci_idat_1
    );
  base_rsci_dat <= base_rsc_dat;
  base_rsci_idat <= base_rsci_idat_1;

  m_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => m_rsci_dat,
      idat => m_rsci_idat_1
    );
  m_rsci_dat <= m_rsc_dat;
  m_rsci_idat <= m_rsci_idat_1;

  return_rsci : work.mgc_out_dreg_pkg_v2.mgc_out_dreg_v2
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      d => return_rsci_d_1,
      z => return_rsci_z
    );
  return_rsci_d_1 <= return_rsci_d;
  return_rsc_z <= return_rsci_z;

  ccs_ccore_start_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 8,
      width => 1
      )
    PORT MAP(
      dat => ccs_ccore_start_rsci_dat,
      idat => ccs_ccore_start_rsci_idat_1
    );
  ccs_ccore_start_rsci_dat(0) <= ccs_ccore_start_rsc_dat;
  ccs_ccore_start_rsci_idat <= ccs_ccore_start_rsci_idat_1(0);

  result_rem_12_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_a_1,
      b => result_rem_12_cmp_b_1,
      z => result_rem_12_cmp_z_1
    );
  result_rem_12_cmp_a_1 <= result_rem_12_cmp_a;
  result_rem_12_cmp_b_1 <= result_rem_12_cmp_b;
  result_rem_12_cmp_z <= result_rem_12_cmp_z_1;

  result_rem_12_cmp_1 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_1_a_1,
      b => result_rem_12_cmp_1_b_1,
      z => result_rem_12_cmp_1_z_1
    );
  result_rem_12_cmp_1_a_1 <= result_rem_12_cmp_1_a;
  result_rem_12_cmp_1_b_1 <= result_rem_12_cmp_1_b;
  result_rem_12_cmp_1_z <= result_rem_12_cmp_1_z_1;

  result_rem_12_cmp_2 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_2_a_1,
      b => result_rem_12_cmp_2_b_1,
      z => result_rem_12_cmp_2_z_1
    );
  result_rem_12_cmp_2_a_1 <= result_rem_12_cmp_2_a;
  result_rem_12_cmp_2_b_1 <= result_rem_12_cmp_2_b;
  result_rem_12_cmp_2_z <= result_rem_12_cmp_2_z_1;

  result_rem_12_cmp_3 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_3_a_1,
      b => result_rem_12_cmp_3_b_1,
      z => result_rem_12_cmp_3_z_1
    );
  result_rem_12_cmp_3_a_1 <= result_rem_12_cmp_3_a;
  result_rem_12_cmp_3_b_1 <= result_rem_12_cmp_3_b;
  result_rem_12_cmp_3_z <= result_rem_12_cmp_3_z_1;

  result_rem_12_cmp_4 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_4_a_1,
      b => result_rem_12_cmp_4_b_1,
      z => result_rem_12_cmp_4_z_1
    );
  result_rem_12_cmp_4_a_1 <= result_rem_12_cmp_4_a;
  result_rem_12_cmp_4_b_1 <= result_rem_12_cmp_4_b;
  result_rem_12_cmp_4_z <= result_rem_12_cmp_4_z_1;

  result_rem_12_cmp_5 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_5_a_1,
      b => result_rem_12_cmp_5_b_1,
      z => result_rem_12_cmp_5_z_1
    );
  result_rem_12_cmp_5_a_1 <= result_rem_12_cmp_5_a;
  result_rem_12_cmp_5_b_1 <= result_rem_12_cmp_5_b;
  result_rem_12_cmp_5_z <= result_rem_12_cmp_5_z_1;

  result_rem_12_cmp_6 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_6_a_1,
      b => result_rem_12_cmp_6_b_1,
      z => result_rem_12_cmp_6_z_1
    );
  result_rem_12_cmp_6_a_1 <= result_rem_12_cmp_6_a;
  result_rem_12_cmp_6_b_1 <= result_rem_12_cmp_6_b;
  result_rem_12_cmp_6_z <= result_rem_12_cmp_6_z_1;

  result_rem_12_cmp_7 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_7_a_1,
      b => result_rem_12_cmp_7_b_1,
      z => result_rem_12_cmp_7_z_1
    );
  result_rem_12_cmp_7_a_1 <= result_rem_12_cmp_7_a;
  result_rem_12_cmp_7_b_1 <= result_rem_12_cmp_7_b;
  result_rem_12_cmp_7_z <= result_rem_12_cmp_7_z_1;

  result_rem_12_cmp_8 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_8_a_1,
      b => result_rem_12_cmp_8_b_1,
      z => result_rem_12_cmp_8_z_1
    );
  result_rem_12_cmp_8_a_1 <= result_rem_12_cmp_8_a;
  result_rem_12_cmp_8_b_1 <= result_rem_12_cmp_8_b;
  result_rem_12_cmp_8_z <= result_rem_12_cmp_8_z_1;

  result_rem_12_cmp_9 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_9_a_1,
      b => result_rem_12_cmp_9_b_1,
      z => result_rem_12_cmp_9_z_1
    );
  result_rem_12_cmp_9_a_1 <= result_rem_12_cmp_9_a;
  result_rem_12_cmp_9_b_1 <= result_rem_12_cmp_9_b;
  result_rem_12_cmp_9_z <= result_rem_12_cmp_9_z_1;

  result_rem_12_cmp_10 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_10_a_1,
      b => result_rem_12_cmp_10_b_1,
      z => result_rem_12_cmp_10_z_1
    );
  result_rem_12_cmp_10_a_1 <= result_rem_12_cmp_10_a;
  result_rem_12_cmp_10_b_1 <= result_rem_12_cmp_10_b;
  result_rem_12_cmp_10_z <= result_rem_12_cmp_10_z_1;

  result_and_1_cse <= ccs_ccore_en AND (and_dcpl_263 OR and_dcpl_269 OR and_dcpl_275
      OR and_dcpl_281 OR and_dcpl_287 OR and_dcpl_293 OR and_dcpl_299 OR and_dcpl_305
      OR and_dcpl_311 OR mux_tmp_37);
  result_and_3_cse <= ccs_ccore_en AND (and_dcpl_319 OR and_dcpl_322 OR and_dcpl_325
      OR and_dcpl_329 OR and_dcpl_333 OR and_dcpl_337 OR and_dcpl_341 OR and_dcpl_344
      OR and_dcpl_347 OR mux_tmp_75);
  result_and_5_cse <= ccs_ccore_en AND (and_dcpl_353 OR and_dcpl_357 OR and_dcpl_361
      OR and_dcpl_364 OR and_dcpl_367 OR and_dcpl_370 OR and_dcpl_373 OR and_dcpl_377
      OR and_dcpl_381 OR mux_tmp_113);
  result_and_7_cse <= ccs_ccore_en AND (and_dcpl_387 OR and_dcpl_390 OR and_dcpl_393
      OR and_dcpl_396 OR and_dcpl_399 OR and_dcpl_402 OR and_dcpl_405 OR and_dcpl_408
      OR and_dcpl_411 OR mux_tmp_151);
  result_and_9_cse <= ccs_ccore_en AND (and_dcpl_418 OR and_dcpl_422 OR and_dcpl_426
      OR and_dcpl_430 OR and_dcpl_433 OR and_dcpl_437 OR and_dcpl_441 OR and_dcpl_444
      OR and_dcpl_447 OR mux_tmp_189);
  result_and_11_cse <= ccs_ccore_en AND (and_dcpl_452 OR and_dcpl_455 OR and_dcpl_458
      OR and_dcpl_462 OR and_dcpl_464 OR and_dcpl_468 OR and_dcpl_472 OR and_dcpl_474
      OR and_dcpl_476 OR mux_tmp_227);
  result_and_13_cse <= ccs_ccore_en AND (and_dcpl_480 OR and_dcpl_484 OR and_dcpl_488
      OR and_dcpl_491 OR and_dcpl_493 OR and_dcpl_496 OR and_dcpl_499 OR and_dcpl_501
      OR and_dcpl_503 OR mux_tmp_265);
  result_and_15_cse <= ccs_ccore_en AND (and_dcpl_507 OR and_dcpl_510 OR and_dcpl_513
      OR and_dcpl_516 OR and_dcpl_518 OR and_dcpl_521 OR and_dcpl_524 OR and_dcpl_526
      OR and_dcpl_528 OR mux_tmp_303);
  result_and_17_cse <= ccs_ccore_en AND (and_dcpl_533 OR and_dcpl_536 OR and_dcpl_539
      OR and_dcpl_542 OR and_dcpl_546 OR and_dcpl_549 OR and_dcpl_552 OR and_dcpl_556
      OR and_dcpl_560 OR mux_tmp_348);
  result_and_19_cse <= ccs_ccore_en AND (and_dcpl_566 OR and_dcpl_568 OR and_dcpl_570
      OR and_dcpl_572 OR and_dcpl_576 OR and_dcpl_578 OR and_dcpl_580 OR and_dcpl_583
      OR and_dcpl_586 OR mux_tmp_393);
  result_and_21_cse <= ccs_ccore_en AND (and_dcpl_590 OR and_dcpl_592 OR and_dcpl_594
      OR and_dcpl_596 OR and_dcpl_599 OR and_dcpl_601 OR and_dcpl_603 OR and_dcpl_607
      OR and_dcpl_611 OR mux_tmp_438);
  m_and_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_2;
  m_and_1_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_6;
  m_and_2_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_9;
  m_and_3_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_11;
  m_and_4_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_2;
  m_and_5_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_6;
  m_and_6_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_9;
  m_and_7_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_11;
  m_and_8_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (NOT (result_rem_11cyc_st_9(0)));
  m_and_9_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (result_rem_11cyc_st_9(0));
  m_and_10_cse <= ccs_ccore_en AND and_dcpl_4 AND (result_rem_11cyc_st_9(3)) AND
      (result_rem_11cyc_st_9(1)) AND (NOT (result_rem_11cyc_st_9(0)));
  m_and_11_cse <= ccs_ccore_en AND and_dcpl_30;
  m_and_12_cse <= ccs_ccore_en AND and_dcpl_32;
  m_and_13_cse <= ccs_ccore_en AND and_dcpl_35;
  m_and_14_cse <= ccs_ccore_en AND and_dcpl_37;
  m_and_15_cse <= ccs_ccore_en AND and_dcpl_39;
  m_and_16_cse <= ccs_ccore_en AND and_dcpl_40;
  m_and_17_cse <= ccs_ccore_en AND and_dcpl_41;
  m_and_18_cse <= ccs_ccore_en AND and_dcpl_42;
  m_and_19_cse <= ccs_ccore_en AND and_dcpl_45;
  m_and_20_cse <= ccs_ccore_en AND and_dcpl_47;
  m_and_21_cse <= ccs_ccore_en AND and_dcpl_50;
  m_and_22_cse <= ccs_ccore_en AND and_dcpl_55;
  m_and_23_cse <= ccs_ccore_en AND and_dcpl_58;
  m_and_24_cse <= ccs_ccore_en AND and_dcpl_60;
  m_and_25_cse <= ccs_ccore_en AND and_dcpl_62;
  m_and_26_cse <= ccs_ccore_en AND and_dcpl_65;
  m_and_27_cse <= ccs_ccore_en AND and_dcpl_68;
  m_and_28_cse <= ccs_ccore_en AND and_dcpl_70;
  m_and_29_cse <= ccs_ccore_en AND and_dcpl_72;
  m_and_30_cse <= ccs_ccore_en AND and_dcpl_74;
  m_and_31_cse <= ccs_ccore_en AND and_dcpl_75;
  m_and_32_cse <= ccs_ccore_en AND and_dcpl_76;
  m_and_33_cse <= ccs_ccore_en AND and_dcpl_81;
  m_and_34_cse <= ccs_ccore_en AND and_dcpl_84;
  m_and_35_cse <= ccs_ccore_en AND and_dcpl_86;
  m_and_36_cse <= ccs_ccore_en AND and_dcpl_88;
  m_and_37_cse <= ccs_ccore_en AND and_dcpl_91;
  m_and_38_cse <= ccs_ccore_en AND and_dcpl_94;
  m_and_39_cse <= ccs_ccore_en AND and_dcpl_96;
  m_and_40_cse <= ccs_ccore_en AND and_dcpl_98;
  m_and_41_cse <= ccs_ccore_en AND and_dcpl_100;
  m_and_42_cse <= ccs_ccore_en AND and_dcpl_101;
  m_and_43_cse <= ccs_ccore_en AND and_dcpl_102;
  m_and_44_cse <= ccs_ccore_en AND and_dcpl_107;
  m_and_45_cse <= ccs_ccore_en AND and_dcpl_110;
  m_and_46_cse <= ccs_ccore_en AND and_dcpl_112;
  m_and_47_cse <= ccs_ccore_en AND and_dcpl_114;
  m_and_48_cse <= ccs_ccore_en AND and_dcpl_116;
  m_and_49_cse <= ccs_ccore_en AND and_dcpl_117;
  m_and_50_cse <= ccs_ccore_en AND and_dcpl_118;
  m_and_51_cse <= ccs_ccore_en AND and_dcpl_119;
  m_and_52_cse <= ccs_ccore_en AND and_dcpl_122;
  m_and_53_cse <= ccs_ccore_en AND and_dcpl_125;
  m_and_54_cse <= ccs_ccore_en AND and_dcpl_127;
  m_and_55_cse <= ccs_ccore_en AND and_dcpl_132;
  m_and_56_cse <= ccs_ccore_en AND and_dcpl_135;
  m_and_57_cse <= ccs_ccore_en AND and_dcpl_137;
  m_and_58_cse <= ccs_ccore_en AND and_dcpl_139;
  m_and_59_cse <= ccs_ccore_en AND and_dcpl_142;
  m_and_60_cse <= ccs_ccore_en AND and_dcpl_145;
  m_and_61_cse <= ccs_ccore_en AND and_dcpl_147;
  m_and_62_cse <= ccs_ccore_en AND and_dcpl_149;
  m_and_63_cse <= ccs_ccore_en AND and_dcpl_151;
  m_and_64_cse <= ccs_ccore_en AND and_dcpl_152;
  m_and_65_cse <= ccs_ccore_en AND and_dcpl_153;
  m_and_66_cse <= ccs_ccore_en AND and_dcpl_158;
  m_and_67_cse <= ccs_ccore_en AND and_dcpl_160;
  m_and_68_cse <= ccs_ccore_en AND and_dcpl_163;
  m_and_69_cse <= ccs_ccore_en AND and_dcpl_165;
  m_and_70_cse <= ccs_ccore_en AND and_dcpl_168;
  m_and_71_cse <= ccs_ccore_en AND and_dcpl_170;
  m_and_72_cse <= ccs_ccore_en AND and_dcpl_173;
  m_and_73_cse <= ccs_ccore_en AND and_dcpl_175;
  m_and_74_cse <= ccs_ccore_en AND and_dcpl_177;
  m_and_75_cse <= ccs_ccore_en AND and_dcpl_178;
  m_and_76_cse <= ccs_ccore_en AND and_dcpl_179;
  m_and_77_cse <= ccs_ccore_en AND and_dcpl_184;
  m_and_78_cse <= ccs_ccore_en AND and_dcpl_186;
  m_and_79_cse <= ccs_ccore_en AND and_dcpl_189;
  m_and_80_cse <= ccs_ccore_en AND and_dcpl_191;
  m_and_81_cse <= ccs_ccore_en AND and_dcpl_194;
  m_and_82_cse <= ccs_ccore_en AND and_dcpl_196;
  m_and_83_cse <= ccs_ccore_en AND and_dcpl_199;
  m_and_84_cse <= ccs_ccore_en AND and_dcpl_201;
  m_and_85_cse <= ccs_ccore_en AND and_dcpl_203;
  m_and_86_cse <= ccs_ccore_en AND and_dcpl_204;
  m_and_87_cse <= ccs_ccore_en AND and_dcpl_205;
  m_and_88_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_207;
  m_and_89_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_212;
  m_and_90_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_214;
  m_and_91_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_211 AND (result_rem_11cyc(1));
  m_and_92_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_218 AND (NOT (result_rem_11cyc(1)));
  m_and_93_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_221 AND (NOT (result_rem_11cyc(1)));
  m_and_94_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_218 AND (result_rem_11cyc(1));
  m_and_95_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_221 AND (result_rem_11cyc(1));
  m_and_96_cse <= ccs_ccore_en AND and_dcpl_228 AND and_dcpl_207;
  m_and_97_cse <= ccs_ccore_en AND and_dcpl_228 AND and_dcpl_212;
  m_and_98_cse <= ccs_ccore_en AND and_dcpl_228 AND and_dcpl_214;
  result_result_acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(CONV_SIGNED(CONV_SIGNED(result_acc_imod_1(3),
      1),2)), 2), 4) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(result_acc_imod_1(2 DOWNTO
      0)), 3), 4), 4));
  result_acc_imod_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(result_acc_idiv_1(2
      DOWNTO 0)), 3), 4) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED((NOT (result_acc_idiv_1(3)))
      & STD_LOGIC_VECTOR'( "00")), 3), 4) + CONV_SIGNED(CONV_SIGNED(SIGNED(STD_LOGIC_VECTOR'(
      "10") & (result_acc_idiv_1(3))), 3), 4), 4));
  result_acc_idiv_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(result_rem_11cyc)
      + UNSIGNED'( "0001"), 4));
  and_dcpl_1 <= NOT((result_rem_11cyc_st_9(3)) OR (result_rem_11cyc_st_9(1)));
  and_dcpl_2 <= and_dcpl_1 AND (NOT (result_rem_11cyc_st_9(0)));
  and_dcpl_3 <= main_stage_0_10 AND asn_itm_9;
  and_dcpl_4 <= and_dcpl_3 AND (NOT (result_rem_11cyc_st_9(2)));
  and_dcpl_6 <= and_dcpl_1 AND (result_rem_11cyc_st_9(0));
  and_dcpl_8 <= (NOT (result_rem_11cyc_st_9(3))) AND (result_rem_11cyc_st_9(1));
  and_dcpl_9 <= and_dcpl_8 AND (NOT (result_rem_11cyc_st_9(0)));
  and_dcpl_11 <= and_dcpl_8 AND (result_rem_11cyc_st_9(0));
  and_dcpl_13 <= and_dcpl_3 AND (result_rem_11cyc_st_9(2));
  and_dcpl_18 <= (result_rem_11cyc_st_9(3)) AND (NOT (result_rem_11cyc_st_9(1)));
  and_dcpl_26 <= NOT((result_rem_11cyc_st_8(3)) OR (result_rem_11cyc_st_8(1)));
  and_dcpl_27 <= and_dcpl_26 AND (NOT (result_rem_11cyc_st_8(0)));
  and_dcpl_28 <= main_stage_0_9 AND asn_itm_8;
  and_dcpl_29 <= and_dcpl_28 AND (NOT (result_rem_11cyc_st_8(2)));
  and_dcpl_30 <= and_dcpl_29 AND and_dcpl_27;
  and_dcpl_31 <= and_dcpl_26 AND (result_rem_11cyc_st_8(0));
  and_dcpl_32 <= and_dcpl_29 AND and_dcpl_31;
  and_dcpl_33 <= (NOT (result_rem_11cyc_st_8(3))) AND (result_rem_11cyc_st_8(1));
  and_dcpl_34 <= and_dcpl_33 AND (NOT (result_rem_11cyc_st_8(0)));
  and_dcpl_35 <= and_dcpl_29 AND and_dcpl_34;
  and_dcpl_36 <= and_dcpl_33 AND (result_rem_11cyc_st_8(0));
  and_dcpl_37 <= and_dcpl_29 AND and_dcpl_36;
  and_dcpl_38 <= and_dcpl_28 AND (result_rem_11cyc_st_8(2));
  and_dcpl_39 <= and_dcpl_38 AND and_dcpl_27;
  and_dcpl_40 <= and_dcpl_38 AND and_dcpl_31;
  and_dcpl_41 <= and_dcpl_38 AND and_dcpl_34;
  and_dcpl_42 <= and_dcpl_38 AND and_dcpl_36;
  and_dcpl_43 <= (result_rem_11cyc_st_8(3)) AND (NOT (result_rem_11cyc_st_8(1)));
  and_dcpl_45 <= and_dcpl_29 AND and_dcpl_43 AND (NOT (result_rem_11cyc_st_8(0)));
  and_dcpl_47 <= and_dcpl_29 AND and_dcpl_43 AND (result_rem_11cyc_st_8(0));
  and_dcpl_50 <= and_dcpl_29 AND (result_rem_11cyc_st_8(3)) AND (result_rem_11cyc_st_8(1))
      AND (NOT (result_rem_11cyc_st_8(0)));
  and_dcpl_51 <= NOT((result_rem_11cyc_st_7(2)) OR (result_rem_11cyc_st_7(0)));
  and_dcpl_52 <= and_dcpl_51 AND (NOT (result_rem_11cyc_st_7(1)));
  and_dcpl_53 <= main_stage_0_8 AND asn_itm_7;
  and_dcpl_54 <= and_dcpl_53 AND (NOT (result_rem_11cyc_st_7(3)));
  and_dcpl_55 <= and_dcpl_54 AND and_dcpl_52;
  and_dcpl_56 <= (NOT (result_rem_11cyc_st_7(2))) AND (result_rem_11cyc_st_7(0));
  and_dcpl_57 <= and_dcpl_56 AND (NOT (result_rem_11cyc_st_7(1)));
  and_dcpl_58 <= and_dcpl_54 AND and_dcpl_57;
  and_dcpl_59 <= and_dcpl_51 AND (result_rem_11cyc_st_7(1));
  and_dcpl_60 <= and_dcpl_54 AND and_dcpl_59;
  and_dcpl_62 <= and_dcpl_54 AND and_dcpl_56 AND (result_rem_11cyc_st_7(1));
  and_dcpl_63 <= (result_rem_11cyc_st_7(2)) AND (NOT (result_rem_11cyc_st_7(0)));
  and_dcpl_65 <= and_dcpl_54 AND and_dcpl_63 AND (NOT (result_rem_11cyc_st_7(1)));
  and_dcpl_66 <= (result_rem_11cyc_st_7(2)) AND (result_rem_11cyc_st_7(0));
  and_dcpl_68 <= and_dcpl_54 AND and_dcpl_66 AND (NOT (result_rem_11cyc_st_7(1)));
  and_dcpl_70 <= and_dcpl_54 AND and_dcpl_63 AND (result_rem_11cyc_st_7(1));
  and_dcpl_72 <= and_dcpl_54 AND and_dcpl_66 AND (result_rem_11cyc_st_7(1));
  and_dcpl_73 <= and_dcpl_53 AND (result_rem_11cyc_st_7(3));
  and_dcpl_74 <= and_dcpl_73 AND and_dcpl_52;
  and_dcpl_75 <= and_dcpl_73 AND and_dcpl_57;
  and_dcpl_76 <= and_dcpl_73 AND and_dcpl_59;
  and_dcpl_77 <= NOT((result_rem_11cyc_st_6(2)) OR (result_rem_11cyc_st_6(0)));
  and_dcpl_78 <= and_dcpl_77 AND (NOT (result_rem_11cyc_st_6(1)));
  and_dcpl_79 <= main_stage_0_7 AND asn_itm_6;
  and_dcpl_80 <= and_dcpl_79 AND (NOT (result_rem_11cyc_st_6(3)));
  and_dcpl_81 <= and_dcpl_80 AND and_dcpl_78;
  and_dcpl_82 <= (NOT (result_rem_11cyc_st_6(2))) AND (result_rem_11cyc_st_6(0));
  and_dcpl_83 <= and_dcpl_82 AND (NOT (result_rem_11cyc_st_6(1)));
  and_dcpl_84 <= and_dcpl_80 AND and_dcpl_83;
  and_dcpl_85 <= and_dcpl_77 AND (result_rem_11cyc_st_6(1));
  and_dcpl_86 <= and_dcpl_80 AND and_dcpl_85;
  and_dcpl_88 <= and_dcpl_80 AND and_dcpl_82 AND (result_rem_11cyc_st_6(1));
  and_dcpl_89 <= (result_rem_11cyc_st_6(2)) AND (NOT (result_rem_11cyc_st_6(0)));
  and_dcpl_91 <= and_dcpl_80 AND and_dcpl_89 AND (NOT (result_rem_11cyc_st_6(1)));
  and_dcpl_92 <= (result_rem_11cyc_st_6(2)) AND (result_rem_11cyc_st_6(0));
  and_dcpl_94 <= and_dcpl_80 AND and_dcpl_92 AND (NOT (result_rem_11cyc_st_6(1)));
  and_dcpl_96 <= and_dcpl_80 AND and_dcpl_89 AND (result_rem_11cyc_st_6(1));
  and_dcpl_98 <= and_dcpl_80 AND and_dcpl_92 AND (result_rem_11cyc_st_6(1));
  and_dcpl_99 <= and_dcpl_79 AND (result_rem_11cyc_st_6(3));
  and_dcpl_100 <= and_dcpl_99 AND and_dcpl_78;
  and_dcpl_101 <= and_dcpl_99 AND and_dcpl_83;
  and_dcpl_102 <= and_dcpl_99 AND and_dcpl_85;
  and_dcpl_103 <= NOT((result_rem_11cyc_st_5(3)) OR (result_rem_11cyc_st_5(0)));
  and_dcpl_104 <= and_dcpl_103 AND (NOT (result_rem_11cyc_st_5(1)));
  and_dcpl_105 <= main_stage_0_6 AND asn_itm_5;
  and_dcpl_106 <= and_dcpl_105 AND (NOT (result_rem_11cyc_st_5(2)));
  and_dcpl_107 <= and_dcpl_106 AND and_dcpl_104;
  and_dcpl_108 <= (NOT (result_rem_11cyc_st_5(3))) AND (result_rem_11cyc_st_5(0));
  and_dcpl_109 <= and_dcpl_108 AND (NOT (result_rem_11cyc_st_5(1)));
  and_dcpl_110 <= and_dcpl_106 AND and_dcpl_109;
  and_dcpl_111 <= and_dcpl_103 AND (result_rem_11cyc_st_5(1));
  and_dcpl_112 <= and_dcpl_106 AND and_dcpl_111;
  and_dcpl_113 <= and_dcpl_108 AND (result_rem_11cyc_st_5(1));
  and_dcpl_114 <= and_dcpl_106 AND and_dcpl_113;
  and_dcpl_115 <= and_dcpl_105 AND (result_rem_11cyc_st_5(2));
  and_dcpl_116 <= and_dcpl_115 AND and_dcpl_104;
  and_dcpl_117 <= and_dcpl_115 AND and_dcpl_109;
  and_dcpl_118 <= and_dcpl_115 AND and_dcpl_111;
  and_dcpl_119 <= and_dcpl_115 AND and_dcpl_113;
  and_dcpl_120 <= (result_rem_11cyc_st_5(3)) AND (NOT (result_rem_11cyc_st_5(0)));
  and_dcpl_122 <= and_dcpl_106 AND and_dcpl_120 AND (NOT (result_rem_11cyc_st_5(1)));
  and_dcpl_125 <= and_dcpl_106 AND (result_rem_11cyc_st_5(3)) AND (result_rem_11cyc_st_5(0))
      AND (NOT (result_rem_11cyc_st_5(1)));
  and_dcpl_127 <= and_dcpl_106 AND and_dcpl_120 AND (result_rem_11cyc_st_5(1));
  and_dcpl_128 <= NOT((result_rem_11cyc_st_4(2)) OR (result_rem_11cyc_st_4(0)));
  and_dcpl_129 <= and_dcpl_128 AND (NOT (result_rem_11cyc_st_4(1)));
  and_dcpl_130 <= main_stage_0_5 AND asn_itm_4;
  and_dcpl_131 <= and_dcpl_130 AND (NOT (result_rem_11cyc_st_4(3)));
  and_dcpl_132 <= and_dcpl_131 AND and_dcpl_129;
  and_dcpl_133 <= (NOT (result_rem_11cyc_st_4(2))) AND (result_rem_11cyc_st_4(0));
  and_dcpl_134 <= and_dcpl_133 AND (NOT (result_rem_11cyc_st_4(1)));
  and_dcpl_135 <= and_dcpl_131 AND and_dcpl_134;
  and_dcpl_136 <= and_dcpl_128 AND (result_rem_11cyc_st_4(1));
  and_dcpl_137 <= and_dcpl_131 AND and_dcpl_136;
  and_dcpl_139 <= and_dcpl_131 AND and_dcpl_133 AND (result_rem_11cyc_st_4(1));
  and_dcpl_140 <= (result_rem_11cyc_st_4(2)) AND (NOT (result_rem_11cyc_st_4(0)));
  and_dcpl_142 <= and_dcpl_131 AND and_dcpl_140 AND (NOT (result_rem_11cyc_st_4(1)));
  and_dcpl_143 <= (result_rem_11cyc_st_4(2)) AND (result_rem_11cyc_st_4(0));
  and_dcpl_145 <= and_dcpl_131 AND and_dcpl_143 AND (NOT (result_rem_11cyc_st_4(1)));
  and_dcpl_147 <= and_dcpl_131 AND and_dcpl_140 AND (result_rem_11cyc_st_4(1));
  and_dcpl_149 <= and_dcpl_131 AND and_dcpl_143 AND (result_rem_11cyc_st_4(1));
  and_dcpl_150 <= and_dcpl_130 AND (result_rem_11cyc_st_4(3));
  and_dcpl_151 <= and_dcpl_150 AND and_dcpl_129;
  and_dcpl_152 <= and_dcpl_150 AND and_dcpl_134;
  and_dcpl_153 <= and_dcpl_150 AND and_dcpl_136;
  and_dcpl_154 <= NOT(CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_155 <= and_dcpl_154 AND (NOT (result_rem_11cyc_st_3(0)));
  and_dcpl_156 <= main_stage_0_4 AND asn_itm_3;
  and_dcpl_157 <= and_dcpl_156 AND (NOT (result_rem_11cyc_st_3(3)));
  and_dcpl_158 <= and_dcpl_157 AND and_dcpl_155;
  and_dcpl_159 <= and_dcpl_154 AND (result_rem_11cyc_st_3(0));
  and_dcpl_160 <= and_dcpl_157 AND and_dcpl_159;
  and_dcpl_161 <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_162 <= and_dcpl_161 AND (NOT (result_rem_11cyc_st_3(0)));
  and_dcpl_163 <= and_dcpl_157 AND and_dcpl_162;
  and_dcpl_165 <= and_dcpl_157 AND and_dcpl_161 AND (result_rem_11cyc_st_3(0));
  and_dcpl_166 <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_168 <= and_dcpl_157 AND and_dcpl_166 AND (NOT (result_rem_11cyc_st_3(0)));
  and_dcpl_170 <= and_dcpl_157 AND and_dcpl_166 AND (result_rem_11cyc_st_3(0));
  and_dcpl_171 <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_173 <= and_dcpl_157 AND and_dcpl_171 AND (NOT (result_rem_11cyc_st_3(0)));
  and_dcpl_175 <= and_dcpl_157 AND and_dcpl_171 AND (result_rem_11cyc_st_3(0));
  and_dcpl_176 <= and_dcpl_156 AND (result_rem_11cyc_st_3(3));
  and_dcpl_177 <= and_dcpl_176 AND and_dcpl_155;
  and_dcpl_178 <= and_dcpl_176 AND and_dcpl_159;
  and_dcpl_179 <= and_dcpl_176 AND and_dcpl_162;
  and_dcpl_180 <= NOT(CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_181 <= and_dcpl_180 AND (NOT (result_rem_11cyc_st_2(0)));
  and_dcpl_182 <= main_stage_0_3 AND asn_itm_2;
  and_dcpl_183 <= and_dcpl_182 AND (NOT (result_rem_11cyc_st_2(3)));
  and_dcpl_184 <= and_dcpl_183 AND and_dcpl_181;
  and_dcpl_185 <= and_dcpl_180 AND (result_rem_11cyc_st_2(0));
  and_dcpl_186 <= and_dcpl_183 AND and_dcpl_185;
  and_dcpl_187 <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_188 <= and_dcpl_187 AND (NOT (result_rem_11cyc_st_2(0)));
  and_dcpl_189 <= and_dcpl_183 AND and_dcpl_188;
  and_dcpl_191 <= and_dcpl_183 AND and_dcpl_187 AND (result_rem_11cyc_st_2(0));
  and_dcpl_192 <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_194 <= and_dcpl_183 AND and_dcpl_192 AND (NOT (result_rem_11cyc_st_2(0)));
  and_dcpl_196 <= and_dcpl_183 AND and_dcpl_192 AND (result_rem_11cyc_st_2(0));
  and_dcpl_197 <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_199 <= and_dcpl_183 AND and_dcpl_197 AND (NOT (result_rem_11cyc_st_2(0)));
  and_dcpl_201 <= and_dcpl_183 AND and_dcpl_197 AND (result_rem_11cyc_st_2(0));
  and_dcpl_202 <= and_dcpl_182 AND (result_rem_11cyc_st_2(3));
  and_dcpl_203 <= and_dcpl_202 AND and_dcpl_181;
  and_dcpl_204 <= and_dcpl_202 AND and_dcpl_185;
  and_dcpl_205 <= and_dcpl_202 AND and_dcpl_188;
  and_dcpl_206 <= NOT((result_rem_11cyc(2)) OR (result_rem_11cyc(0)));
  and_dcpl_207 <= and_dcpl_206 AND (NOT (result_rem_11cyc(1)));
  and_dcpl_208 <= main_stage_0_2 AND asn_itm_1;
  and_dcpl_209 <= and_dcpl_208 AND (NOT (result_rem_11cyc(3)));
  and_dcpl_211 <= (NOT (result_rem_11cyc(2))) AND (result_rem_11cyc(0));
  and_dcpl_212 <= and_dcpl_211 AND (NOT (result_rem_11cyc(1)));
  and_dcpl_214 <= and_dcpl_206 AND (result_rem_11cyc(1));
  and_dcpl_218 <= (result_rem_11cyc(2)) AND (NOT (result_rem_11cyc(0)));
  and_dcpl_221 <= (result_rem_11cyc(2)) AND (result_rem_11cyc(0));
  and_dcpl_228 <= and_dcpl_208 AND (result_rem_11cyc(3));
  and_dcpl_232 <= NOT(CONV_SL_1_1(result_rem_11cyc_st_11(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_233 <= and_dcpl_232 AND (NOT (result_rem_11cyc_st_11(0)));
  and_dcpl_234 <= main_stage_0_12 AND asn_itm_11;
  and_dcpl_235 <= and_dcpl_234 AND (NOT (result_rem_11cyc_st_11(3)));
  and_dcpl_237 <= and_dcpl_232 AND (result_rem_11cyc_st_11(0));
  and_dcpl_239 <= CONV_SL_1_1(result_rem_11cyc_st_11(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_240 <= and_dcpl_239 AND (NOT (result_rem_11cyc_st_11(0)));
  and_dcpl_244 <= CONV_SL_1_1(result_rem_11cyc_st_11(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_249 <= CONV_SL_1_1(result_rem_11cyc_st_11(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_254 <= and_dcpl_234 AND (result_rem_11cyc_st_11(3));
  and_dcpl_260 <= NOT(CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_261 <= ccs_ccore_start_rsci_idat AND (NOT (result_result_acc_tmp(2)));
  and_dcpl_262 <= and_dcpl_261 AND (NOT (result_result_acc_tmp(3)));
  and_dcpl_263 <= and_dcpl_262 AND and_dcpl_260;
  or_tmp_2 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0000")) OR (NOT and_dcpl_208);
  or_3_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0000"));
  nor_691_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_2));
  mux_nl <= MUX_s_1_2_2(nor_691_nl, or_tmp_2, or_3_cse);
  and_dcpl_269 <= mux_nl AND and_dcpl_184;
  or_8_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0000"));
  nor_690_nl <= NOT(and_dcpl_208 OR and_dcpl_184);
  or_10_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_182);
  mux_tmp_1 <= MUX_s_1_2_2(nor_690_nl, or_10_nl, or_8_cse);
  nor_689_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_1));
  mux_2_nl <= MUX_s_1_2_2(nor_689_nl, mux_tmp_1, or_3_cse);
  and_dcpl_275 <= mux_2_nl AND and_dcpl_158;
  or_15_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0000"));
  nor_687_nl <= NOT(and_dcpl_182 OR and_dcpl_158);
  or_17_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_156);
  mux_tmp_3 <= MUX_s_1_2_2(nor_687_nl, or_17_nl, or_15_cse);
  nor_688_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_3));
  mux_tmp_4 <= MUX_s_1_2_2(nor_688_nl, mux_tmp_3, or_8_cse);
  nor_686_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_4));
  mux_5_nl <= MUX_s_1_2_2(nor_686_nl, mux_tmp_4, or_3_cse);
  and_dcpl_281 <= mux_5_nl AND and_dcpl_132;
  or_24_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0000"));
  nor_683_nl <= NOT(and_dcpl_156 OR and_dcpl_132);
  or_26_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_130);
  mux_tmp_6 <= MUX_s_1_2_2(nor_683_nl, or_26_nl, or_24_cse);
  nor_684_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_6));
  mux_tmp_7 <= MUX_s_1_2_2(nor_684_nl, mux_tmp_6, or_15_cse);
  nor_685_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_7));
  mux_tmp_8 <= MUX_s_1_2_2(nor_685_nl, mux_tmp_7, or_8_cse);
  nor_682_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_8));
  mux_9_nl <= MUX_s_1_2_2(nor_682_nl, mux_tmp_8, or_3_cse);
  and_dcpl_287 <= mux_9_nl AND and_dcpl_107;
  or_35_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0000"));
  nor_678_nl <= NOT(and_dcpl_130 OR and_dcpl_107);
  or_37_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_105);
  mux_tmp_10 <= MUX_s_1_2_2(nor_678_nl, or_37_nl, or_35_cse);
  nor_679_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_10));
  mux_tmp_11 <= MUX_s_1_2_2(nor_679_nl, mux_tmp_10, or_24_cse);
  nor_680_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_11));
  mux_tmp_12 <= MUX_s_1_2_2(nor_680_nl, mux_tmp_11, or_15_cse);
  nor_681_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_12));
  mux_tmp_13 <= MUX_s_1_2_2(nor_681_nl, mux_tmp_12, or_8_cse);
  nor_677_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_13));
  mux_14_nl <= MUX_s_1_2_2(nor_677_nl, mux_tmp_13, or_3_cse);
  and_dcpl_293 <= mux_14_nl AND and_dcpl_81;
  or_48_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0000"));
  nor_672_nl <= NOT(and_dcpl_105 OR and_dcpl_81);
  or_50_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_79);
  mux_tmp_15 <= MUX_s_1_2_2(nor_672_nl, or_50_nl, or_48_cse);
  nor_673_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_15));
  mux_tmp_16 <= MUX_s_1_2_2(nor_673_nl, mux_tmp_15, or_35_cse);
  nor_674_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_16));
  mux_tmp_17 <= MUX_s_1_2_2(nor_674_nl, mux_tmp_16, or_24_cse);
  nor_675_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_17));
  mux_tmp_18 <= MUX_s_1_2_2(nor_675_nl, mux_tmp_17, or_15_cse);
  nor_676_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_18));
  mux_tmp_19 <= MUX_s_1_2_2(nor_676_nl, mux_tmp_18, or_8_cse);
  nor_671_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_19));
  mux_20_nl <= MUX_s_1_2_2(nor_671_nl, mux_tmp_19, or_3_cse);
  and_dcpl_299 <= mux_20_nl AND and_dcpl_55;
  or_63_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0000"));
  nor_665_nl <= NOT(and_dcpl_79 OR and_dcpl_55);
  or_65_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_53);
  mux_tmp_21 <= MUX_s_1_2_2(nor_665_nl, or_65_nl, or_63_cse);
  nor_666_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_21));
  mux_tmp_22 <= MUX_s_1_2_2(nor_666_nl, mux_tmp_21, or_48_cse);
  nor_667_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_22));
  mux_tmp_23 <= MUX_s_1_2_2(nor_667_nl, mux_tmp_22, or_35_cse);
  nor_668_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_23));
  mux_tmp_24 <= MUX_s_1_2_2(nor_668_nl, mux_tmp_23, or_24_cse);
  nor_669_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_24));
  mux_tmp_25 <= MUX_s_1_2_2(nor_669_nl, mux_tmp_24, or_15_cse);
  nor_670_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_25));
  mux_tmp_26 <= MUX_s_1_2_2(nor_670_nl, mux_tmp_25, or_8_cse);
  nor_664_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_26));
  mux_27_nl <= MUX_s_1_2_2(nor_664_nl, mux_tmp_26, or_3_cse);
  and_dcpl_305 <= mux_27_nl AND and_dcpl_30;
  nor_656_nl <= NOT(and_dcpl_53 OR and_dcpl_30);
  or_82_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_28);
  or_80_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0000"));
  mux_tmp_28 <= MUX_s_1_2_2(nor_656_nl, or_82_nl, or_80_nl);
  nor_657_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_28));
  mux_tmp_29 <= MUX_s_1_2_2(nor_657_nl, mux_tmp_28, or_63_cse);
  nor_658_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_29));
  mux_tmp_30 <= MUX_s_1_2_2(nor_658_nl, mux_tmp_29, or_48_cse);
  nor_659_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_30));
  mux_tmp_31 <= MUX_s_1_2_2(nor_659_nl, mux_tmp_30, or_35_cse);
  nor_660_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_31));
  mux_tmp_32 <= MUX_s_1_2_2(nor_660_nl, mux_tmp_31, or_24_cse);
  nor_661_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_32));
  mux_tmp_33 <= MUX_s_1_2_2(nor_661_nl, mux_tmp_32, or_15_cse);
  nor_662_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_33));
  mux_tmp_34 <= MUX_s_1_2_2(nor_662_nl, mux_tmp_33, or_8_cse);
  nor_663_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_34));
  mux_35_nl <= MUX_s_1_2_2(nor_663_nl, mux_tmp_34, or_3_cse);
  and_dcpl_311 <= mux_35_nl AND and_dcpl_4 AND and_dcpl_2;
  and_tmp_6 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0000")));
  nor_654_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_6));
  mux_tmp_36 <= MUX_s_1_2_2(nor_654_nl, and_tmp_6, or_8_cse);
  nor_655_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_36));
  mux_tmp_37 <= MUX_s_1_2_2(nor_655_nl, mux_tmp_36, or_3_cse);
  and_dcpl_318 <= CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_319 <= and_dcpl_262 AND and_dcpl_318;
  or_tmp_102 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_208);
  or_107_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0001"));
  nor_653_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_102));
  mux_38_nl <= MUX_s_1_2_2(nor_653_nl, or_tmp_102, or_107_cse);
  and_dcpl_322 <= mux_38_nl AND and_dcpl_186;
  or_112_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0001"));
  nor_652_nl <= NOT(and_dcpl_208 OR and_dcpl_186);
  or_114_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_182);
  mux_tmp_39 <= MUX_s_1_2_2(nor_652_nl, or_114_nl, or_112_cse);
  nor_651_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_39));
  mux_40_nl <= MUX_s_1_2_2(nor_651_nl, mux_tmp_39, or_107_cse);
  and_dcpl_325 <= mux_40_nl AND and_dcpl_160;
  or_119_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0001"));
  nor_649_nl <= NOT(and_dcpl_182 OR and_dcpl_160);
  or_121_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_156);
  mux_tmp_41 <= MUX_s_1_2_2(nor_649_nl, or_121_nl, or_119_cse);
  nor_650_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_41));
  mux_tmp_42 <= MUX_s_1_2_2(nor_650_nl, mux_tmp_41, or_112_cse);
  nor_648_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_42));
  mux_43_nl <= MUX_s_1_2_2(nor_648_nl, mux_tmp_42, or_107_cse);
  and_dcpl_329 <= mux_43_nl AND and_dcpl_135;
  or_128_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0001"));
  nor_645_nl <= NOT(and_dcpl_156 OR and_dcpl_135);
  or_130_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_130);
  mux_tmp_44 <= MUX_s_1_2_2(nor_645_nl, or_130_nl, or_128_cse);
  nor_646_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_44));
  mux_tmp_45 <= MUX_s_1_2_2(nor_646_nl, mux_tmp_44, or_119_cse);
  nor_647_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_45));
  mux_tmp_46 <= MUX_s_1_2_2(nor_647_nl, mux_tmp_45, or_112_cse);
  nor_644_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_46));
  mux_47_nl <= MUX_s_1_2_2(nor_644_nl, mux_tmp_46, or_107_cse);
  and_dcpl_333 <= mux_47_nl AND and_dcpl_110;
  or_139_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0001"));
  nor_640_nl <= NOT(and_dcpl_130 OR and_dcpl_110);
  or_141_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_105);
  mux_tmp_48 <= MUX_s_1_2_2(nor_640_nl, or_141_nl, or_139_cse);
  nor_641_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_48));
  mux_tmp_49 <= MUX_s_1_2_2(nor_641_nl, mux_tmp_48, or_128_cse);
  nor_642_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_49));
  mux_tmp_50 <= MUX_s_1_2_2(nor_642_nl, mux_tmp_49, or_119_cse);
  nor_643_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_50));
  mux_tmp_51 <= MUX_s_1_2_2(nor_643_nl, mux_tmp_50, or_112_cse);
  nor_639_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_51));
  mux_52_nl <= MUX_s_1_2_2(nor_639_nl, mux_tmp_51, or_107_cse);
  and_dcpl_337 <= mux_52_nl AND and_dcpl_84;
  or_152_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0001"));
  nor_634_nl <= NOT(and_dcpl_105 OR and_dcpl_84);
  or_154_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_79);
  mux_tmp_53 <= MUX_s_1_2_2(nor_634_nl, or_154_nl, or_152_cse);
  nor_635_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_53));
  mux_tmp_54 <= MUX_s_1_2_2(nor_635_nl, mux_tmp_53, or_139_cse);
  nor_636_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_54));
  mux_tmp_55 <= MUX_s_1_2_2(nor_636_nl, mux_tmp_54, or_128_cse);
  nor_637_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_55));
  mux_tmp_56 <= MUX_s_1_2_2(nor_637_nl, mux_tmp_55, or_119_cse);
  nor_638_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_56));
  mux_tmp_57 <= MUX_s_1_2_2(nor_638_nl, mux_tmp_56, or_112_cse);
  nor_633_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_57));
  mux_58_nl <= MUX_s_1_2_2(nor_633_nl, mux_tmp_57, or_107_cse);
  and_dcpl_341 <= mux_58_nl AND and_dcpl_58;
  or_167_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0001"));
  nor_627_nl <= NOT(and_dcpl_79 OR and_dcpl_58);
  or_169_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_53);
  mux_tmp_59 <= MUX_s_1_2_2(nor_627_nl, or_169_nl, or_167_cse);
  nor_628_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_59));
  mux_tmp_60 <= MUX_s_1_2_2(nor_628_nl, mux_tmp_59, or_152_cse);
  nor_629_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_60));
  mux_tmp_61 <= MUX_s_1_2_2(nor_629_nl, mux_tmp_60, or_139_cse);
  nor_630_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_61));
  mux_tmp_62 <= MUX_s_1_2_2(nor_630_nl, mux_tmp_61, or_128_cse);
  nor_631_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_62));
  mux_tmp_63 <= MUX_s_1_2_2(nor_631_nl, mux_tmp_62, or_119_cse);
  nor_632_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_63));
  mux_tmp_64 <= MUX_s_1_2_2(nor_632_nl, mux_tmp_63, or_112_cse);
  nor_626_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_64));
  mux_65_nl <= MUX_s_1_2_2(nor_626_nl, mux_tmp_64, or_107_cse);
  and_dcpl_344 <= mux_65_nl AND and_dcpl_32;
  nor_618_nl <= NOT(and_dcpl_53 OR and_dcpl_32);
  or_186_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_28);
  or_184_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0001"));
  mux_tmp_66 <= MUX_s_1_2_2(nor_618_nl, or_186_nl, or_184_nl);
  nor_619_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_66));
  mux_tmp_67 <= MUX_s_1_2_2(nor_619_nl, mux_tmp_66, or_167_cse);
  nor_620_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_67));
  mux_tmp_68 <= MUX_s_1_2_2(nor_620_nl, mux_tmp_67, or_152_cse);
  nor_621_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_68));
  mux_tmp_69 <= MUX_s_1_2_2(nor_621_nl, mux_tmp_68, or_139_cse);
  nor_622_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_69));
  mux_tmp_70 <= MUX_s_1_2_2(nor_622_nl, mux_tmp_69, or_128_cse);
  nor_623_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_70));
  mux_tmp_71 <= MUX_s_1_2_2(nor_623_nl, mux_tmp_70, or_119_cse);
  nor_624_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_71));
  mux_tmp_72 <= MUX_s_1_2_2(nor_624_nl, mux_tmp_71, or_112_cse);
  nor_625_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_72));
  mux_73_nl <= MUX_s_1_2_2(nor_625_nl, mux_tmp_72, or_107_cse);
  and_dcpl_347 <= mux_73_nl AND and_dcpl_4 AND and_dcpl_6;
  and_tmp_13 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0001")));
  nor_617_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_13));
  mux_tmp_74 <= MUX_s_1_2_2(nor_617_nl, and_tmp_13, or_112_cse);
  nand_146_cse <= NOT((result_result_acc_tmp(0)) AND ccs_ccore_start_rsci_idat);
  and_797_nl <= nand_146_cse AND mux_tmp_74;
  or_195_nl <= CONV_SL_1_1(result_result_acc_tmp(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_75 <= MUX_s_1_2_2(and_797_nl, mux_tmp_74, or_195_nl);
  and_dcpl_352 <= CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_353 <= and_dcpl_262 AND and_dcpl_352;
  or_tmp_202 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_208);
  or_209_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0010"));
  nor_616_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_202));
  mux_76_nl <= MUX_s_1_2_2(nor_616_nl, or_tmp_202, or_209_cse);
  and_dcpl_357 <= mux_76_nl AND and_dcpl_189;
  or_214_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0010"));
  nor_615_nl <= NOT(and_dcpl_208 OR and_dcpl_189);
  or_216_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_182);
  mux_tmp_77 <= MUX_s_1_2_2(nor_615_nl, or_216_nl, or_214_cse);
  nor_614_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_77));
  mux_78_nl <= MUX_s_1_2_2(nor_614_nl, mux_tmp_77, or_209_cse);
  and_dcpl_361 <= mux_78_nl AND and_dcpl_163;
  or_221_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0010"));
  nor_612_nl <= NOT(and_dcpl_182 OR and_dcpl_163);
  or_223_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_156);
  mux_tmp_79 <= MUX_s_1_2_2(nor_612_nl, or_223_nl, or_221_cse);
  nor_613_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_79));
  mux_tmp_80 <= MUX_s_1_2_2(nor_613_nl, mux_tmp_79, or_214_cse);
  nor_611_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_80));
  mux_81_nl <= MUX_s_1_2_2(nor_611_nl, mux_tmp_80, or_209_cse);
  and_dcpl_364 <= mux_81_nl AND and_dcpl_137;
  or_230_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0010"));
  nor_608_nl <= NOT(and_dcpl_156 OR and_dcpl_137);
  or_232_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_130);
  mux_tmp_82 <= MUX_s_1_2_2(nor_608_nl, or_232_nl, or_230_cse);
  nor_609_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_82));
  mux_tmp_83 <= MUX_s_1_2_2(nor_609_nl, mux_tmp_82, or_221_cse);
  nor_610_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_83));
  mux_tmp_84 <= MUX_s_1_2_2(nor_610_nl, mux_tmp_83, or_214_cse);
  nor_607_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_84));
  mux_85_nl <= MUX_s_1_2_2(nor_607_nl, mux_tmp_84, or_209_cse);
  and_dcpl_367 <= mux_85_nl AND and_dcpl_112;
  or_241_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0010"));
  nor_603_nl <= NOT(and_dcpl_130 OR and_dcpl_112);
  or_243_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_105);
  mux_tmp_86 <= MUX_s_1_2_2(nor_603_nl, or_243_nl, or_241_cse);
  nor_604_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_86));
  mux_tmp_87 <= MUX_s_1_2_2(nor_604_nl, mux_tmp_86, or_230_cse);
  nor_605_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_87));
  mux_tmp_88 <= MUX_s_1_2_2(nor_605_nl, mux_tmp_87, or_221_cse);
  nor_606_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_88));
  mux_tmp_89 <= MUX_s_1_2_2(nor_606_nl, mux_tmp_88, or_214_cse);
  nor_602_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_89));
  mux_90_nl <= MUX_s_1_2_2(nor_602_nl, mux_tmp_89, or_209_cse);
  and_dcpl_370 <= mux_90_nl AND and_dcpl_86;
  or_254_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0010"));
  nor_597_nl <= NOT(and_dcpl_105 OR and_dcpl_86);
  or_256_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_79);
  mux_tmp_91 <= MUX_s_1_2_2(nor_597_nl, or_256_nl, or_254_cse);
  nor_598_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_91));
  mux_tmp_92 <= MUX_s_1_2_2(nor_598_nl, mux_tmp_91, or_241_cse);
  nor_599_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_92));
  mux_tmp_93 <= MUX_s_1_2_2(nor_599_nl, mux_tmp_92, or_230_cse);
  nor_600_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_93));
  mux_tmp_94 <= MUX_s_1_2_2(nor_600_nl, mux_tmp_93, or_221_cse);
  nor_601_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_94));
  mux_tmp_95 <= MUX_s_1_2_2(nor_601_nl, mux_tmp_94, or_214_cse);
  nor_596_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_95));
  mux_96_nl <= MUX_s_1_2_2(nor_596_nl, mux_tmp_95, or_209_cse);
  and_dcpl_373 <= mux_96_nl AND and_dcpl_60;
  or_269_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0010"));
  nor_590_nl <= NOT(and_dcpl_79 OR and_dcpl_60);
  or_271_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_53);
  mux_tmp_97 <= MUX_s_1_2_2(nor_590_nl, or_271_nl, or_269_cse);
  nor_591_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_97));
  mux_tmp_98 <= MUX_s_1_2_2(nor_591_nl, mux_tmp_97, or_254_cse);
  nor_592_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_98));
  mux_tmp_99 <= MUX_s_1_2_2(nor_592_nl, mux_tmp_98, or_241_cse);
  nor_593_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_99));
  mux_tmp_100 <= MUX_s_1_2_2(nor_593_nl, mux_tmp_99, or_230_cse);
  nor_594_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_100));
  mux_tmp_101 <= MUX_s_1_2_2(nor_594_nl, mux_tmp_100, or_221_cse);
  nor_595_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_101));
  mux_tmp_102 <= MUX_s_1_2_2(nor_595_nl, mux_tmp_101, or_214_cse);
  nor_589_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_102));
  mux_103_nl <= MUX_s_1_2_2(nor_589_nl, mux_tmp_102, or_209_cse);
  and_dcpl_377 <= mux_103_nl AND and_dcpl_35;
  nor_581_nl <= NOT(and_dcpl_53 OR and_dcpl_35);
  or_288_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_28);
  or_286_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0010"));
  mux_tmp_104 <= MUX_s_1_2_2(nor_581_nl, or_288_nl, or_286_nl);
  nor_582_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_104));
  mux_tmp_105 <= MUX_s_1_2_2(nor_582_nl, mux_tmp_104, or_269_cse);
  nor_583_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_105));
  mux_tmp_106 <= MUX_s_1_2_2(nor_583_nl, mux_tmp_105, or_254_cse);
  nor_584_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_106));
  mux_tmp_107 <= MUX_s_1_2_2(nor_584_nl, mux_tmp_106, or_241_cse);
  nor_585_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_107));
  mux_tmp_108 <= MUX_s_1_2_2(nor_585_nl, mux_tmp_107, or_230_cse);
  nor_586_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_108));
  mux_tmp_109 <= MUX_s_1_2_2(nor_586_nl, mux_tmp_108, or_221_cse);
  nor_587_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_109));
  mux_tmp_110 <= MUX_s_1_2_2(nor_587_nl, mux_tmp_109, or_214_cse);
  nor_588_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_110));
  mux_111_nl <= MUX_s_1_2_2(nor_588_nl, mux_tmp_110, or_209_cse);
  and_dcpl_381 <= mux_111_nl AND and_dcpl_4 AND and_dcpl_9;
  and_tmp_20 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0010")));
  nor_579_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_20));
  mux_tmp_112 <= MUX_s_1_2_2(nor_579_nl, and_tmp_20, or_214_cse);
  nor_580_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_112));
  mux_tmp_113 <= MUX_s_1_2_2(nor_580_nl, mux_tmp_112, or_209_cse);
  and_dcpl_386 <= CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_387 <= and_dcpl_262 AND and_dcpl_386;
  or_tmp_302 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_208);
  or_311_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0011"));
  nor_578_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_302));
  mux_114_nl <= MUX_s_1_2_2(nor_578_nl, or_tmp_302, or_311_cse);
  and_dcpl_390 <= mux_114_nl AND and_dcpl_191;
  or_316_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0011"));
  nor_577_nl <= NOT(and_dcpl_208 OR and_dcpl_191);
  or_318_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_182);
  mux_tmp_115 <= MUX_s_1_2_2(nor_577_nl, or_318_nl, or_316_cse);
  nor_576_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_115));
  mux_116_nl <= MUX_s_1_2_2(nor_576_nl, mux_tmp_115, or_311_cse);
  and_dcpl_393 <= mux_116_nl AND and_dcpl_165;
  or_323_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0011"));
  nor_574_nl <= NOT(and_dcpl_182 OR and_dcpl_165);
  or_325_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_156);
  mux_tmp_117 <= MUX_s_1_2_2(nor_574_nl, or_325_nl, or_323_cse);
  nor_575_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_117));
  mux_tmp_118 <= MUX_s_1_2_2(nor_575_nl, mux_tmp_117, or_316_cse);
  nor_573_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_118));
  mux_119_nl <= MUX_s_1_2_2(nor_573_nl, mux_tmp_118, or_311_cse);
  and_dcpl_396 <= mux_119_nl AND and_dcpl_139;
  or_332_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0011"));
  nor_570_nl <= NOT(and_dcpl_156 OR and_dcpl_139);
  or_334_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_130);
  mux_tmp_120 <= MUX_s_1_2_2(nor_570_nl, or_334_nl, or_332_cse);
  nor_571_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_120));
  mux_tmp_121 <= MUX_s_1_2_2(nor_571_nl, mux_tmp_120, or_323_cse);
  nor_572_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_121));
  mux_tmp_122 <= MUX_s_1_2_2(nor_572_nl, mux_tmp_121, or_316_cse);
  nor_569_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_122));
  mux_123_nl <= MUX_s_1_2_2(nor_569_nl, mux_tmp_122, or_311_cse);
  and_dcpl_399 <= mux_123_nl AND and_dcpl_114;
  or_343_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0011"));
  nor_565_nl <= NOT(and_dcpl_130 OR and_dcpl_114);
  or_345_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_105);
  mux_tmp_124 <= MUX_s_1_2_2(nor_565_nl, or_345_nl, or_343_cse);
  nor_566_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_124));
  mux_tmp_125 <= MUX_s_1_2_2(nor_566_nl, mux_tmp_124, or_332_cse);
  nor_567_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_125));
  mux_tmp_126 <= MUX_s_1_2_2(nor_567_nl, mux_tmp_125, or_323_cse);
  nor_568_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_126));
  mux_tmp_127 <= MUX_s_1_2_2(nor_568_nl, mux_tmp_126, or_316_cse);
  nor_564_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_127));
  mux_128_nl <= MUX_s_1_2_2(nor_564_nl, mux_tmp_127, or_311_cse);
  and_dcpl_402 <= mux_128_nl AND and_dcpl_88;
  or_356_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0011"));
  nor_559_nl <= NOT(and_dcpl_105 OR and_dcpl_88);
  or_358_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_79);
  mux_tmp_129 <= MUX_s_1_2_2(nor_559_nl, or_358_nl, or_356_cse);
  nor_560_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_129));
  mux_tmp_130 <= MUX_s_1_2_2(nor_560_nl, mux_tmp_129, or_343_cse);
  nor_561_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_130));
  mux_tmp_131 <= MUX_s_1_2_2(nor_561_nl, mux_tmp_130, or_332_cse);
  nor_562_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_131));
  mux_tmp_132 <= MUX_s_1_2_2(nor_562_nl, mux_tmp_131, or_323_cse);
  nor_563_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_132));
  mux_tmp_133 <= MUX_s_1_2_2(nor_563_nl, mux_tmp_132, or_316_cse);
  nor_558_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_133));
  mux_134_nl <= MUX_s_1_2_2(nor_558_nl, mux_tmp_133, or_311_cse);
  and_dcpl_405 <= mux_134_nl AND and_dcpl_62;
  or_371_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0011"));
  nor_552_nl <= NOT(and_dcpl_79 OR and_dcpl_62);
  or_373_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_53);
  mux_tmp_135 <= MUX_s_1_2_2(nor_552_nl, or_373_nl, or_371_cse);
  nor_553_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_135));
  mux_tmp_136 <= MUX_s_1_2_2(nor_553_nl, mux_tmp_135, or_356_cse);
  nor_554_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_136));
  mux_tmp_137 <= MUX_s_1_2_2(nor_554_nl, mux_tmp_136, or_343_cse);
  nor_555_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_137));
  mux_tmp_138 <= MUX_s_1_2_2(nor_555_nl, mux_tmp_137, or_332_cse);
  nor_556_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_138));
  mux_tmp_139 <= MUX_s_1_2_2(nor_556_nl, mux_tmp_138, or_323_cse);
  nor_557_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_139));
  mux_tmp_140 <= MUX_s_1_2_2(nor_557_nl, mux_tmp_139, or_316_cse);
  nor_551_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_140));
  mux_141_nl <= MUX_s_1_2_2(nor_551_nl, mux_tmp_140, or_311_cse);
  and_dcpl_408 <= mux_141_nl AND and_dcpl_37;
  nor_543_nl <= NOT(and_dcpl_53 OR and_dcpl_37);
  or_390_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_28);
  or_388_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0011"));
  mux_tmp_142 <= MUX_s_1_2_2(nor_543_nl, or_390_nl, or_388_nl);
  nor_544_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_142));
  mux_tmp_143 <= MUX_s_1_2_2(nor_544_nl, mux_tmp_142, or_371_cse);
  nor_545_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_143));
  mux_tmp_144 <= MUX_s_1_2_2(nor_545_nl, mux_tmp_143, or_356_cse);
  nor_546_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_144));
  mux_tmp_145 <= MUX_s_1_2_2(nor_546_nl, mux_tmp_144, or_343_cse);
  nor_547_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_145));
  mux_tmp_146 <= MUX_s_1_2_2(nor_547_nl, mux_tmp_145, or_332_cse);
  nor_548_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_146));
  mux_tmp_147 <= MUX_s_1_2_2(nor_548_nl, mux_tmp_146, or_323_cse);
  nor_549_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_147));
  mux_tmp_148 <= MUX_s_1_2_2(nor_549_nl, mux_tmp_147, or_316_cse);
  nor_550_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_148));
  mux_149_nl <= MUX_s_1_2_2(nor_550_nl, mux_tmp_148, or_311_cse);
  and_dcpl_411 <= mux_149_nl AND and_dcpl_4 AND and_dcpl_11;
  and_tmp_27 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0011")));
  nor_542_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_27));
  mux_tmp_150 <= MUX_s_1_2_2(nor_542_nl, and_tmp_27, or_316_cse);
  and_796_nl <= (NOT(CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND ccs_ccore_start_rsci_idat)) AND mux_tmp_150;
  or_399_nl <= CONV_SL_1_1(result_result_acc_tmp(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_151 <= MUX_s_1_2_2(and_796_nl, mux_tmp_150, or_399_nl);
  and_dcpl_417 <= ccs_ccore_start_rsci_idat AND CONV_SL_1_1(result_result_acc_tmp(3
      DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_418 <= and_dcpl_417 AND and_dcpl_260;
  or_tmp_402 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_208);
  nand_144_cse <= NOT((result_result_acc_tmp(2)) AND ccs_ccore_start_rsci_idat);
  or_413_cse <= (result_result_acc_tmp(1)) OR (result_result_acc_tmp(0)) OR (result_result_acc_tmp(3));
  and_795_nl <= nand_144_cse AND or_tmp_402;
  mux_152_nl <= MUX_s_1_2_2(and_795_nl, or_tmp_402, or_413_cse);
  and_dcpl_422 <= mux_152_nl AND and_dcpl_194;
  or_418_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0100"));
  nor_541_nl <= NOT(and_dcpl_208 OR and_dcpl_194);
  or_420_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_182);
  mux_tmp_153 <= MUX_s_1_2_2(nor_541_nl, or_420_nl, or_418_cse);
  and_794_nl <= nand_144_cse AND mux_tmp_153;
  mux_154_nl <= MUX_s_1_2_2(and_794_nl, mux_tmp_153, or_413_cse);
  and_dcpl_426 <= mux_154_nl AND and_dcpl_168;
  or_425_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0100"));
  nor_539_nl <= NOT(and_dcpl_182 OR and_dcpl_168);
  or_427_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_156);
  mux_tmp_155 <= MUX_s_1_2_2(nor_539_nl, or_427_nl, or_425_cse);
  nor_540_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_155));
  mux_tmp_156 <= MUX_s_1_2_2(nor_540_nl, mux_tmp_155, or_418_cse);
  and_793_nl <= nand_144_cse AND mux_tmp_156;
  mux_157_nl <= MUX_s_1_2_2(and_793_nl, mux_tmp_156, or_413_cse);
  and_dcpl_430 <= mux_157_nl AND and_dcpl_142;
  or_434_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0100"));
  nor_536_nl <= NOT(and_dcpl_156 OR and_dcpl_142);
  or_436_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_130);
  mux_tmp_158 <= MUX_s_1_2_2(nor_536_nl, or_436_nl, or_434_cse);
  nor_537_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_158));
  mux_tmp_159 <= MUX_s_1_2_2(nor_537_nl, mux_tmp_158, or_425_cse);
  nor_538_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_159));
  mux_tmp_160 <= MUX_s_1_2_2(nor_538_nl, mux_tmp_159, or_418_cse);
  and_792_nl <= nand_144_cse AND mux_tmp_160;
  mux_161_nl <= MUX_s_1_2_2(and_792_nl, mux_tmp_160, or_413_cse);
  and_dcpl_433 <= mux_161_nl AND and_dcpl_116;
  or_445_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0100"));
  nor_532_nl <= NOT(and_dcpl_130 OR and_dcpl_116);
  or_447_nl <= (result_rem_11cyc_st_5(1)) OR (result_rem_11cyc_st_5(0)) OR (result_rem_11cyc_st_5(3))
      OR (NOT and_dcpl_115);
  mux_tmp_162 <= MUX_s_1_2_2(nor_532_nl, or_447_nl, or_445_cse);
  nor_533_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_162));
  mux_tmp_163 <= MUX_s_1_2_2(nor_533_nl, mux_tmp_162, or_434_cse);
  nor_534_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_163));
  mux_tmp_164 <= MUX_s_1_2_2(nor_534_nl, mux_tmp_163, or_425_cse);
  nor_535_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_164));
  mux_tmp_165 <= MUX_s_1_2_2(nor_535_nl, mux_tmp_164, or_418_cse);
  and_791_nl <= nand_144_cse AND mux_tmp_165;
  mux_166_nl <= MUX_s_1_2_2(and_791_nl, mux_tmp_165, or_413_cse);
  and_dcpl_437 <= mux_166_nl AND and_dcpl_91;
  or_458_cse <= (result_rem_11cyc_st_5(1)) OR (result_rem_11cyc_st_5(0)) OR (result_rem_11cyc_st_5(3));
  and_790_cse <= (result_rem_11cyc_st_5(2)) AND asn_itm_5 AND main_stage_0_6;
  nor_527_nl <= NOT(and_790_cse OR and_dcpl_91);
  or_460_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_79);
  mux_tmp_167 <= MUX_s_1_2_2(nor_527_nl, or_460_nl, or_458_cse);
  nor_528_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_167));
  mux_tmp_168 <= MUX_s_1_2_2(nor_528_nl, mux_tmp_167, or_445_cse);
  nor_529_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_168));
  mux_tmp_169 <= MUX_s_1_2_2(nor_529_nl, mux_tmp_168, or_434_cse);
  nor_530_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_169));
  mux_tmp_170 <= MUX_s_1_2_2(nor_530_nl, mux_tmp_169, or_425_cse);
  nor_531_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_170));
  mux_tmp_171 <= MUX_s_1_2_2(nor_531_nl, mux_tmp_170, or_418_cse);
  and_789_nl <= nand_144_cse AND mux_tmp_171;
  mux_172_nl <= MUX_s_1_2_2(and_789_nl, mux_tmp_171, or_413_cse);
  and_dcpl_441 <= mux_172_nl AND and_dcpl_65;
  or_473_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0100"));
  nor_522_nl <= NOT(and_dcpl_79 OR and_dcpl_65);
  or_475_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_53);
  mux_tmp_173 <= MUX_s_1_2_2(nor_522_nl, or_475_nl, or_473_cse);
  nand_138_cse <= NOT((result_rem_11cyc_st_5(2)) AND asn_itm_5 AND main_stage_0_6);
  and_788_nl <= nand_138_cse AND mux_tmp_173;
  mux_tmp_174 <= MUX_s_1_2_2(and_788_nl, mux_tmp_173, or_458_cse);
  nor_523_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_174));
  mux_tmp_175 <= MUX_s_1_2_2(nor_523_nl, mux_tmp_174, or_445_cse);
  nor_524_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_175));
  mux_tmp_176 <= MUX_s_1_2_2(nor_524_nl, mux_tmp_175, or_434_cse);
  nor_525_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_176));
  mux_tmp_177 <= MUX_s_1_2_2(nor_525_nl, mux_tmp_176, or_425_cse);
  nor_526_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_177));
  mux_tmp_178 <= MUX_s_1_2_2(nor_526_nl, mux_tmp_177, or_418_cse);
  and_787_nl <= nand_144_cse AND mux_tmp_178;
  mux_179_nl <= MUX_s_1_2_2(and_787_nl, mux_tmp_178, or_413_cse);
  and_dcpl_444 <= mux_179_nl AND and_dcpl_39;
  nor_516_nl <= NOT(and_dcpl_53 OR and_dcpl_39);
  or_492_nl <= (result_rem_11cyc_st_8(0)) OR (result_rem_11cyc_st_8(1)) OR (result_rem_11cyc_st_8(3))
      OR (NOT and_dcpl_38);
  or_490_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0100"));
  mux_tmp_180 <= MUX_s_1_2_2(nor_516_nl, or_492_nl, or_490_nl);
  nor_517_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_180));
  mux_tmp_181 <= MUX_s_1_2_2(nor_517_nl, mux_tmp_180, or_473_cse);
  and_785_nl <= nand_138_cse AND mux_tmp_181;
  mux_tmp_182 <= MUX_s_1_2_2(and_785_nl, mux_tmp_181, or_458_cse);
  nor_518_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_182));
  mux_tmp_183 <= MUX_s_1_2_2(nor_518_nl, mux_tmp_182, or_445_cse);
  nor_519_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_183));
  mux_tmp_184 <= MUX_s_1_2_2(nor_519_nl, mux_tmp_183, or_434_cse);
  nor_520_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_184));
  mux_tmp_185 <= MUX_s_1_2_2(nor_520_nl, mux_tmp_184, or_425_cse);
  nor_521_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_185));
  mux_tmp_186 <= MUX_s_1_2_2(nor_521_nl, mux_tmp_185, or_418_cse);
  and_786_nl <= nand_144_cse AND mux_tmp_186;
  mux_187_nl <= MUX_s_1_2_2(and_786_nl, mux_tmp_186, or_413_cse);
  and_dcpl_447 <= mux_187_nl AND and_dcpl_13 AND and_dcpl_2;
  and_tmp_34 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0100")));
  nor_514_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_34));
  mux_tmp_188 <= MUX_s_1_2_2(nor_514_nl, and_tmp_34, or_418_cse);
  nor_515_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_188));
  or_501_nl <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0100"));
  mux_tmp_189 <= MUX_s_1_2_2(nor_515_nl, mux_tmp_188, or_501_nl);
  and_dcpl_452 <= and_dcpl_417 AND and_dcpl_318;
  or_tmp_502 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_208);
  or_516_cse <= (result_result_acc_tmp(1)) OR (NOT (result_result_acc_tmp(0))) OR
      (result_result_acc_tmp(3));
  and_784_nl <= nand_144_cse AND or_tmp_502;
  mux_190_nl <= MUX_s_1_2_2(and_784_nl, or_tmp_502, or_516_cse);
  and_dcpl_455 <= mux_190_nl AND and_dcpl_196;
  or_521_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0101"));
  nor_513_nl <= NOT(and_dcpl_208 OR and_dcpl_196);
  or_523_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_182);
  mux_tmp_191 <= MUX_s_1_2_2(nor_513_nl, or_523_nl, or_521_cse);
  and_783_nl <= nand_144_cse AND mux_tmp_191;
  mux_192_nl <= MUX_s_1_2_2(and_783_nl, mux_tmp_191, or_516_cse);
  and_dcpl_458 <= mux_192_nl AND and_dcpl_170;
  or_528_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0101"));
  nor_511_nl <= NOT(and_dcpl_182 OR and_dcpl_170);
  or_530_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_156);
  mux_tmp_193 <= MUX_s_1_2_2(nor_511_nl, or_530_nl, or_528_cse);
  nor_512_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_193));
  mux_tmp_194 <= MUX_s_1_2_2(nor_512_nl, mux_tmp_193, or_521_cse);
  and_782_nl <= nand_144_cse AND mux_tmp_194;
  mux_195_nl <= MUX_s_1_2_2(and_782_nl, mux_tmp_194, or_516_cse);
  and_dcpl_462 <= mux_195_nl AND and_dcpl_145;
  or_537_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0101"));
  nor_508_nl <= NOT(and_dcpl_156 OR and_dcpl_145);
  or_539_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_130);
  mux_tmp_196 <= MUX_s_1_2_2(nor_508_nl, or_539_nl, or_537_cse);
  nor_509_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_196));
  mux_tmp_197 <= MUX_s_1_2_2(nor_509_nl, mux_tmp_196, or_528_cse);
  nor_510_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_197));
  mux_tmp_198 <= MUX_s_1_2_2(nor_510_nl, mux_tmp_197, or_521_cse);
  and_781_nl <= nand_144_cse AND mux_tmp_198;
  mux_199_nl <= MUX_s_1_2_2(and_781_nl, mux_tmp_198, or_516_cse);
  and_dcpl_464 <= mux_199_nl AND and_dcpl_117;
  or_548_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0101"));
  nor_504_nl <= NOT(and_dcpl_130 OR and_dcpl_117);
  or_550_nl <= (result_rem_11cyc_st_5(1)) OR (NOT (result_rem_11cyc_st_5(0))) OR
      (result_rem_11cyc_st_5(3)) OR (NOT and_dcpl_115);
  mux_tmp_200 <= MUX_s_1_2_2(nor_504_nl, or_550_nl, or_548_cse);
  nor_505_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_200));
  mux_tmp_201 <= MUX_s_1_2_2(nor_505_nl, mux_tmp_200, or_537_cse);
  nor_506_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_201));
  mux_tmp_202 <= MUX_s_1_2_2(nor_506_nl, mux_tmp_201, or_528_cse);
  nor_507_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_202));
  mux_tmp_203 <= MUX_s_1_2_2(nor_507_nl, mux_tmp_202, or_521_cse);
  and_780_nl <= nand_144_cse AND mux_tmp_203;
  mux_204_nl <= MUX_s_1_2_2(and_780_nl, mux_tmp_203, or_516_cse);
  and_dcpl_468 <= mux_204_nl AND and_dcpl_94;
  or_561_cse <= (result_rem_11cyc_st_5(1)) OR (NOT (result_rem_11cyc_st_5(0))) OR
      (result_rem_11cyc_st_5(3));
  nor_499_nl <= NOT(and_790_cse OR and_dcpl_94);
  or_563_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_79);
  mux_tmp_205 <= MUX_s_1_2_2(nor_499_nl, or_563_nl, or_561_cse);
  nor_500_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_205));
  mux_tmp_206 <= MUX_s_1_2_2(nor_500_nl, mux_tmp_205, or_548_cse);
  nor_501_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_206));
  mux_tmp_207 <= MUX_s_1_2_2(nor_501_nl, mux_tmp_206, or_537_cse);
  nor_502_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_207));
  mux_tmp_208 <= MUX_s_1_2_2(nor_502_nl, mux_tmp_207, or_528_cse);
  nor_503_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_208));
  mux_tmp_209 <= MUX_s_1_2_2(nor_503_nl, mux_tmp_208, or_521_cse);
  and_778_nl <= nand_144_cse AND mux_tmp_209;
  mux_210_nl <= MUX_s_1_2_2(and_778_nl, mux_tmp_209, or_516_cse);
  and_dcpl_472 <= mux_210_nl AND and_dcpl_68;
  or_576_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0101"));
  nor_494_nl <= NOT(and_dcpl_79 OR and_dcpl_68);
  or_578_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_53);
  mux_tmp_211 <= MUX_s_1_2_2(nor_494_nl, or_578_nl, or_576_cse);
  and_777_nl <= nand_138_cse AND mux_tmp_211;
  mux_tmp_212 <= MUX_s_1_2_2(and_777_nl, mux_tmp_211, or_561_cse);
  nor_495_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_212));
  mux_tmp_213 <= MUX_s_1_2_2(nor_495_nl, mux_tmp_212, or_548_cse);
  nor_496_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_213));
  mux_tmp_214 <= MUX_s_1_2_2(nor_496_nl, mux_tmp_213, or_537_cse);
  nor_497_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_214));
  mux_tmp_215 <= MUX_s_1_2_2(nor_497_nl, mux_tmp_214, or_528_cse);
  nor_498_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_215));
  mux_tmp_216 <= MUX_s_1_2_2(nor_498_nl, mux_tmp_215, or_521_cse);
  and_776_nl <= nand_144_cse AND mux_tmp_216;
  mux_217_nl <= MUX_s_1_2_2(and_776_nl, mux_tmp_216, or_516_cse);
  and_dcpl_474 <= mux_217_nl AND and_dcpl_40;
  nor_488_nl <= NOT(and_dcpl_53 OR and_dcpl_40);
  or_595_nl <= (NOT (result_rem_11cyc_st_8(0))) OR (result_rem_11cyc_st_8(1)) OR
      (result_rem_11cyc_st_8(3)) OR (NOT and_dcpl_38);
  or_593_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0101"));
  mux_tmp_218 <= MUX_s_1_2_2(nor_488_nl, or_595_nl, or_593_nl);
  nor_489_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_218));
  mux_tmp_219 <= MUX_s_1_2_2(nor_489_nl, mux_tmp_218, or_576_cse);
  and_774_nl <= nand_138_cse AND mux_tmp_219;
  mux_tmp_220 <= MUX_s_1_2_2(and_774_nl, mux_tmp_219, or_561_cse);
  nor_490_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_220));
  mux_tmp_221 <= MUX_s_1_2_2(nor_490_nl, mux_tmp_220, or_548_cse);
  nor_491_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_221));
  mux_tmp_222 <= MUX_s_1_2_2(nor_491_nl, mux_tmp_221, or_537_cse);
  nor_492_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_222));
  mux_tmp_223 <= MUX_s_1_2_2(nor_492_nl, mux_tmp_222, or_528_cse);
  nor_493_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_223));
  mux_tmp_224 <= MUX_s_1_2_2(nor_493_nl, mux_tmp_223, or_521_cse);
  and_775_nl <= nand_144_cse AND mux_tmp_224;
  mux_225_nl <= MUX_s_1_2_2(and_775_nl, mux_tmp_224, or_516_cse);
  and_dcpl_476 <= mux_225_nl AND and_dcpl_13 AND and_dcpl_6;
  and_tmp_41 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0101")));
  nor_487_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_41));
  mux_tmp_226 <= MUX_s_1_2_2(nor_487_nl, and_tmp_41, or_521_cse);
  and_773_nl <= nand_146_cse AND mux_tmp_226;
  or_604_nl <= CONV_SL_1_1(result_result_acc_tmp(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_227 <= MUX_s_1_2_2(and_773_nl, mux_tmp_226, or_604_nl);
  and_dcpl_480 <= and_dcpl_417 AND and_dcpl_352;
  or_tmp_602 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_208);
  or_617_cse <= (NOT (result_result_acc_tmp(1))) OR (result_result_acc_tmp(0)) OR
      (result_result_acc_tmp(3));
  and_772_nl <= nand_144_cse AND or_tmp_602;
  mux_228_nl <= MUX_s_1_2_2(and_772_nl, or_tmp_602, or_617_cse);
  and_dcpl_484 <= mux_228_nl AND and_dcpl_199;
  or_622_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0110"));
  nor_486_nl <= NOT(and_dcpl_208 OR and_dcpl_199);
  or_624_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_182);
  mux_tmp_229 <= MUX_s_1_2_2(nor_486_nl, or_624_nl, or_622_cse);
  and_771_nl <= nand_144_cse AND mux_tmp_229;
  mux_230_nl <= MUX_s_1_2_2(and_771_nl, mux_tmp_229, or_617_cse);
  and_dcpl_488 <= mux_230_nl AND and_dcpl_173;
  or_629_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0110"));
  nor_484_nl <= NOT(and_dcpl_182 OR and_dcpl_173);
  or_631_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_156);
  mux_tmp_231 <= MUX_s_1_2_2(nor_484_nl, or_631_nl, or_629_cse);
  nor_485_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_231));
  mux_tmp_232 <= MUX_s_1_2_2(nor_485_nl, mux_tmp_231, or_622_cse);
  and_770_nl <= nand_144_cse AND mux_tmp_232;
  mux_233_nl <= MUX_s_1_2_2(and_770_nl, mux_tmp_232, or_617_cse);
  and_dcpl_491 <= mux_233_nl AND and_dcpl_147;
  or_638_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0110"));
  nor_481_nl <= NOT(and_dcpl_156 OR and_dcpl_147);
  or_640_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_130);
  mux_tmp_234 <= MUX_s_1_2_2(nor_481_nl, or_640_nl, or_638_cse);
  nor_482_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_234));
  mux_tmp_235 <= MUX_s_1_2_2(nor_482_nl, mux_tmp_234, or_629_cse);
  nor_483_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_235));
  mux_tmp_236 <= MUX_s_1_2_2(nor_483_nl, mux_tmp_235, or_622_cse);
  and_769_nl <= nand_144_cse AND mux_tmp_236;
  mux_237_nl <= MUX_s_1_2_2(and_769_nl, mux_tmp_236, or_617_cse);
  and_dcpl_493 <= mux_237_nl AND and_dcpl_118;
  or_649_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0110"));
  nor_477_nl <= NOT(and_dcpl_130 OR and_dcpl_118);
  or_651_nl <= (NOT (result_rem_11cyc_st_5(1))) OR (result_rem_11cyc_st_5(0)) OR
      (result_rem_11cyc_st_5(3)) OR (NOT and_dcpl_115);
  mux_tmp_238 <= MUX_s_1_2_2(nor_477_nl, or_651_nl, or_649_cse);
  nor_478_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_238));
  mux_tmp_239 <= MUX_s_1_2_2(nor_478_nl, mux_tmp_238, or_638_cse);
  nor_479_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_239));
  mux_tmp_240 <= MUX_s_1_2_2(nor_479_nl, mux_tmp_239, or_629_cse);
  nor_480_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_240));
  mux_tmp_241 <= MUX_s_1_2_2(nor_480_nl, mux_tmp_240, or_622_cse);
  and_768_nl <= nand_144_cse AND mux_tmp_241;
  mux_242_nl <= MUX_s_1_2_2(and_768_nl, mux_tmp_241, or_617_cse);
  and_dcpl_496 <= mux_242_nl AND and_dcpl_96;
  or_662_cse <= (NOT (result_rem_11cyc_st_5(1))) OR (result_rem_11cyc_st_5(0)) OR
      (result_rem_11cyc_st_5(3));
  nor_472_nl <= NOT(and_790_cse OR and_dcpl_96);
  or_664_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_79);
  mux_tmp_243 <= MUX_s_1_2_2(nor_472_nl, or_664_nl, or_662_cse);
  nor_473_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_243));
  mux_tmp_244 <= MUX_s_1_2_2(nor_473_nl, mux_tmp_243, or_649_cse);
  nor_474_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_244));
  mux_tmp_245 <= MUX_s_1_2_2(nor_474_nl, mux_tmp_244, or_638_cse);
  nor_475_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_245));
  mux_tmp_246 <= MUX_s_1_2_2(nor_475_nl, mux_tmp_245, or_629_cse);
  nor_476_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_246));
  mux_tmp_247 <= MUX_s_1_2_2(nor_476_nl, mux_tmp_246, or_622_cse);
  and_766_nl <= nand_144_cse AND mux_tmp_247;
  mux_248_nl <= MUX_s_1_2_2(and_766_nl, mux_tmp_247, or_617_cse);
  and_dcpl_499 <= mux_248_nl AND and_dcpl_70;
  or_677_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0110"));
  nor_467_nl <= NOT(and_dcpl_79 OR and_dcpl_70);
  or_679_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_53);
  mux_tmp_249 <= MUX_s_1_2_2(nor_467_nl, or_679_nl, or_677_cse);
  and_765_nl <= nand_138_cse AND mux_tmp_249;
  mux_tmp_250 <= MUX_s_1_2_2(and_765_nl, mux_tmp_249, or_662_cse);
  nor_468_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_250));
  mux_tmp_251 <= MUX_s_1_2_2(nor_468_nl, mux_tmp_250, or_649_cse);
  nor_469_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_251));
  mux_tmp_252 <= MUX_s_1_2_2(nor_469_nl, mux_tmp_251, or_638_cse);
  nor_470_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_252));
  mux_tmp_253 <= MUX_s_1_2_2(nor_470_nl, mux_tmp_252, or_629_cse);
  nor_471_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_253));
  mux_tmp_254 <= MUX_s_1_2_2(nor_471_nl, mux_tmp_253, or_622_cse);
  and_764_nl <= nand_144_cse AND mux_tmp_254;
  mux_255_nl <= MUX_s_1_2_2(and_764_nl, mux_tmp_254, or_617_cse);
  and_dcpl_501 <= mux_255_nl AND and_dcpl_41;
  nor_461_nl <= NOT(and_dcpl_53 OR and_dcpl_41);
  or_696_nl <= (result_rem_11cyc_st_8(0)) OR (NOT (result_rem_11cyc_st_8(1))) OR
      (result_rem_11cyc_st_8(3)) OR (NOT and_dcpl_38);
  or_694_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0110"));
  mux_tmp_256 <= MUX_s_1_2_2(nor_461_nl, or_696_nl, or_694_nl);
  nor_462_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_256));
  mux_tmp_257 <= MUX_s_1_2_2(nor_462_nl, mux_tmp_256, or_677_cse);
  and_762_nl <= nand_138_cse AND mux_tmp_257;
  mux_tmp_258 <= MUX_s_1_2_2(and_762_nl, mux_tmp_257, or_662_cse);
  nor_463_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_258));
  mux_tmp_259 <= MUX_s_1_2_2(nor_463_nl, mux_tmp_258, or_649_cse);
  nor_464_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_259));
  mux_tmp_260 <= MUX_s_1_2_2(nor_464_nl, mux_tmp_259, or_638_cse);
  nor_465_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_260));
  mux_tmp_261 <= MUX_s_1_2_2(nor_465_nl, mux_tmp_260, or_629_cse);
  nor_466_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_261));
  mux_tmp_262 <= MUX_s_1_2_2(nor_466_nl, mux_tmp_261, or_622_cse);
  and_763_nl <= nand_144_cse AND mux_tmp_262;
  mux_263_nl <= MUX_s_1_2_2(and_763_nl, mux_tmp_262, or_617_cse);
  and_dcpl_503 <= mux_263_nl AND and_dcpl_13 AND and_dcpl_9;
  and_tmp_48 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0110")));
  nor_459_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_48));
  mux_tmp_264 <= MUX_s_1_2_2(nor_459_nl, and_tmp_48, or_622_cse);
  nor_460_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_264));
  or_705_nl <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0110"));
  mux_tmp_265 <= MUX_s_1_2_2(nor_460_nl, mux_tmp_264, or_705_nl);
  and_dcpl_507 <= and_dcpl_417 AND and_dcpl_386;
  or_tmp_702 <= NOT(CONV_SL_1_1(result_rem_11cyc=STD_LOGIC_VECTOR'("0111")) AND and_dcpl_208);
  or_718_cse <= (NOT (result_result_acc_tmp(1))) OR (NOT (result_result_acc_tmp(0)))
      OR (result_result_acc_tmp(3));
  and_761_nl <= nand_144_cse AND or_tmp_702;
  mux_266_nl <= MUX_s_1_2_2(and_761_nl, or_tmp_702, or_718_cse);
  and_dcpl_510 <= mux_266_nl AND and_dcpl_201;
  nand_112_cse <= NOT(CONV_SL_1_1(result_rem_11cyc=STD_LOGIC_VECTOR'("0111")));
  nor_458_nl <= NOT(and_dcpl_208 OR and_dcpl_201);
  nand_153_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_2=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_182);
  mux_tmp_267 <= MUX_s_1_2_2(nor_458_nl, nand_153_nl, nand_112_cse);
  and_760_nl <= nand_144_cse AND mux_tmp_267;
  mux_268_nl <= MUX_s_1_2_2(and_760_nl, mux_tmp_267, or_718_cse);
  and_dcpl_513 <= mux_268_nl AND and_dcpl_175;
  nand_108_cse <= NOT(CONV_SL_1_1(result_rem_11cyc_st_2=STD_LOGIC_VECTOR'("0111")));
  nor_456_nl <= NOT(and_dcpl_182 OR and_dcpl_175);
  nand_152_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_3=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_156);
  mux_tmp_269 <= MUX_s_1_2_2(nor_456_nl, nand_152_nl, nand_108_cse);
  nor_457_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_269));
  mux_tmp_270 <= MUX_s_1_2_2(nor_457_nl, mux_tmp_269, nand_112_cse);
  and_759_nl <= nand_144_cse AND mux_tmp_270;
  mux_271_nl <= MUX_s_1_2_2(and_759_nl, mux_tmp_270, or_718_cse);
  and_dcpl_516 <= mux_271_nl AND and_dcpl_149;
  nand_103_cse <= NOT(CONV_SL_1_1(result_rem_11cyc_st_3=STD_LOGIC_VECTOR'("0111")));
  nor_453_nl <= NOT(and_dcpl_156 OR and_dcpl_149);
  nand_151_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_4=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_130);
  mux_tmp_272 <= MUX_s_1_2_2(nor_453_nl, nand_151_nl, nand_103_cse);
  nor_454_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_272));
  mux_tmp_273 <= MUX_s_1_2_2(nor_454_nl, mux_tmp_272, nand_108_cse);
  nor_455_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_273));
  mux_tmp_274 <= MUX_s_1_2_2(nor_455_nl, mux_tmp_273, nand_112_cse);
  and_758_nl <= nand_144_cse AND mux_tmp_274;
  mux_275_nl <= MUX_s_1_2_2(and_758_nl, mux_tmp_274, or_718_cse);
  and_dcpl_518 <= mux_275_nl AND and_dcpl_119;
  nand_97_cse <= NOT(CONV_SL_1_1(result_rem_11cyc_st_4=STD_LOGIC_VECTOR'("0111")));
  nor_449_nl <= NOT(and_dcpl_130 OR and_dcpl_119);
  nand_96_nl <= NOT((result_rem_11cyc_st_5(1)) AND (result_rem_11cyc_st_5(0)) AND
      (NOT (result_rem_11cyc_st_5(3))) AND and_dcpl_115);
  mux_tmp_276 <= MUX_s_1_2_2(nor_449_nl, nand_96_nl, nand_97_cse);
  nor_450_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_276));
  mux_tmp_277 <= MUX_s_1_2_2(nor_450_nl, mux_tmp_276, nand_103_cse);
  nor_451_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_277));
  mux_tmp_278 <= MUX_s_1_2_2(nor_451_nl, mux_tmp_277, nand_108_cse);
  nor_452_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_278));
  mux_tmp_279 <= MUX_s_1_2_2(nor_452_nl, mux_tmp_278, nand_112_cse);
  and_757_nl <= nand_144_cse AND mux_tmp_279;
  mux_280_nl <= MUX_s_1_2_2(and_757_nl, mux_tmp_279, or_718_cse);
  and_dcpl_521 <= mux_280_nl AND and_dcpl_98;
  or_763_cse <= (NOT (result_rem_11cyc_st_5(1))) OR (NOT (result_rem_11cyc_st_5(0)))
      OR (result_rem_11cyc_st_5(3));
  nor_444_nl <= NOT(and_790_cse OR and_dcpl_98);
  nand_150_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_6=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_79);
  mux_tmp_281 <= MUX_s_1_2_2(nor_444_nl, nand_150_nl, or_763_cse);
  nor_445_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_281));
  mux_tmp_282 <= MUX_s_1_2_2(nor_445_nl, mux_tmp_281, nand_97_cse);
  nor_446_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_282));
  mux_tmp_283 <= MUX_s_1_2_2(nor_446_nl, mux_tmp_282, nand_103_cse);
  nor_447_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_283));
  mux_tmp_284 <= MUX_s_1_2_2(nor_447_nl, mux_tmp_283, nand_108_cse);
  nor_448_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_284));
  mux_tmp_285 <= MUX_s_1_2_2(nor_448_nl, mux_tmp_284, nand_112_cse);
  and_755_nl <= nand_144_cse AND mux_tmp_285;
  mux_286_nl <= MUX_s_1_2_2(and_755_nl, mux_tmp_285, or_718_cse);
  and_dcpl_524 <= mux_286_nl AND and_dcpl_72;
  nand_83_cse <= NOT(CONV_SL_1_1(result_rem_11cyc_st_6=STD_LOGIC_VECTOR'("0111")));
  nor_439_nl <= NOT(and_dcpl_79 OR and_dcpl_72);
  nand_149_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_7=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_53);
  mux_tmp_287 <= MUX_s_1_2_2(nor_439_nl, nand_149_nl, nand_83_cse);
  and_754_nl <= nand_138_cse AND mux_tmp_287;
  mux_tmp_288 <= MUX_s_1_2_2(and_754_nl, mux_tmp_287, or_763_cse);
  nor_440_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_288));
  mux_tmp_289 <= MUX_s_1_2_2(nor_440_nl, mux_tmp_288, nand_97_cse);
  nor_441_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_289));
  mux_tmp_290 <= MUX_s_1_2_2(nor_441_nl, mux_tmp_289, nand_103_cse);
  nor_442_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_290));
  mux_tmp_291 <= MUX_s_1_2_2(nor_442_nl, mux_tmp_290, nand_108_cse);
  nor_443_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_291));
  mux_tmp_292 <= MUX_s_1_2_2(nor_443_nl, mux_tmp_291, nand_112_cse);
  and_753_nl <= nand_144_cse AND mux_tmp_292;
  mux_293_nl <= MUX_s_1_2_2(and_753_nl, mux_tmp_292, or_718_cse);
  and_dcpl_526 <= mux_293_nl AND and_dcpl_42;
  nor_433_nl <= NOT(and_dcpl_53 OR and_dcpl_42);
  nand_72_nl <= NOT((result_rem_11cyc_st_8(0)) AND (result_rem_11cyc_st_8(1)) AND
      (NOT (result_rem_11cyc_st_8(3))) AND and_dcpl_38);
  nand_73_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_7=STD_LOGIC_VECTOR'("0111")));
  mux_tmp_294 <= MUX_s_1_2_2(nor_433_nl, nand_72_nl, nand_73_nl);
  nor_434_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_294));
  mux_tmp_295 <= MUX_s_1_2_2(nor_434_nl, mux_tmp_294, nand_83_cse);
  and_751_nl <= nand_138_cse AND mux_tmp_295;
  mux_tmp_296 <= MUX_s_1_2_2(and_751_nl, mux_tmp_295, or_763_cse);
  nor_435_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_296));
  mux_tmp_297 <= MUX_s_1_2_2(nor_435_nl, mux_tmp_296, nand_97_cse);
  nor_436_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_297));
  mux_tmp_298 <= MUX_s_1_2_2(nor_436_nl, mux_tmp_297, nand_103_cse);
  nor_437_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_298));
  mux_tmp_299 <= MUX_s_1_2_2(nor_437_nl, mux_tmp_298, nand_108_cse);
  nor_438_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_299));
  mux_tmp_300 <= MUX_s_1_2_2(nor_438_nl, mux_tmp_299, nand_112_cse);
  and_752_nl <= nand_144_cse AND mux_tmp_300;
  mux_301_nl <= MUX_s_1_2_2(and_752_nl, mux_tmp_300, or_718_cse);
  and_dcpl_528 <= mux_301_nl AND and_dcpl_13 AND and_dcpl_11;
  and_tmp_55 <= (NOT(main_stage_0_3 AND asn_itm_2 AND CONV_SL_1_1(result_rem_11cyc_st_2=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_4 AND asn_itm_3 AND CONV_SL_1_1(result_rem_11cyc_st_3=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_5 AND asn_itm_4 AND CONV_SL_1_1(result_rem_11cyc_st_4=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_6 AND asn_itm_5 AND CONV_SL_1_1(result_rem_11cyc_st_5=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_7 AND asn_itm_6 AND CONV_SL_1_1(result_rem_11cyc_st_6=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_8 AND asn_itm_7 AND CONV_SL_1_1(result_rem_11cyc_st_7=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_9 AND asn_itm_8 AND CONV_SL_1_1(result_rem_11cyc_st_8=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_10 AND asn_itm_9 AND CONV_SL_1_1(result_rem_11cyc_st_9=STD_LOGIC_VECTOR'("0111"))));
  nor_432_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_55));
  mux_tmp_302 <= MUX_s_1_2_2(nor_432_nl, and_tmp_55, nand_112_cse);
  and_750_nl <= (NOT(CONV_SL_1_1(result_result_acc_tmp(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND ccs_ccore_start_rsci_idat)) AND mux_tmp_302;
  mux_tmp_303 <= MUX_s_1_2_2(and_750_nl, mux_tmp_302, result_result_acc_tmp(3));
  and_dcpl_532 <= and_dcpl_261 AND (result_result_acc_tmp(3));
  and_dcpl_533 <= and_dcpl_532 AND and_dcpl_260;
  not_tmp_645 <= NOT((result_rem_11cyc(3)) AND asn_itm_1 AND main_stage_0_2);
  or_tmp_801 <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR not_tmp_645;
  or_818_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("1000"));
  nor_431_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_801));
  mux_304_nl <= MUX_s_1_2_2(nor_431_nl, or_tmp_801, or_818_cse);
  and_dcpl_536 <= mux_304_nl AND and_dcpl_203;
  or_823_cse <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_749_cse <= (result_rem_11cyc(3)) AND asn_itm_1 AND main_stage_0_2;
  nor_430_nl <= NOT(and_749_cse OR and_dcpl_203);
  or_825_nl <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_202);
  mux_tmp_305 <= MUX_s_1_2_2(nor_430_nl, or_825_nl, or_823_cse);
  nor_429_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_305));
  mux_306_nl <= MUX_s_1_2_2(nor_429_nl, mux_tmp_305, or_818_cse);
  and_dcpl_539 <= mux_306_nl AND and_dcpl_177;
  or_830_cse <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_747_cse <= (result_rem_11cyc_st_2(3)) AND asn_itm_2 AND main_stage_0_3;
  nor_428_nl <= NOT(and_747_cse OR and_dcpl_177);
  or_832_nl <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_176);
  mux_tmp_307 <= MUX_s_1_2_2(nor_428_nl, or_832_nl, or_830_cse);
  and_748_nl <= not_tmp_645 AND mux_tmp_307;
  mux_tmp_308 <= MUX_s_1_2_2(and_748_nl, mux_tmp_307, or_823_cse);
  nor_427_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_308));
  mux_309_nl <= MUX_s_1_2_2(nor_427_nl, mux_tmp_308, or_818_cse);
  and_dcpl_542 <= mux_309_nl AND and_dcpl_151;
  or_839_cse <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_744_cse <= (result_rem_11cyc_st_3(3)) AND asn_itm_3 AND main_stage_0_4;
  nor_426_nl <= NOT(and_744_cse OR and_dcpl_151);
  or_841_nl <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_150);
  mux_tmp_310 <= MUX_s_1_2_2(nor_426_nl, or_841_nl, or_839_cse);
  nand_58_cse <= NOT((result_rem_11cyc_st_2(3)) AND asn_itm_2 AND main_stage_0_3);
  and_745_nl <= nand_58_cse AND mux_tmp_310;
  mux_tmp_311 <= MUX_s_1_2_2(and_745_nl, mux_tmp_310, or_830_cse);
  and_746_nl <= not_tmp_645 AND mux_tmp_311;
  mux_tmp_312 <= MUX_s_1_2_2(and_746_nl, mux_tmp_311, or_823_cse);
  nor_425_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_312));
  mux_313_nl <= MUX_s_1_2_2(nor_425_nl, mux_tmp_312, or_818_cse);
  and_dcpl_546 <= mux_313_nl AND and_dcpl_122;
  or_850_cse <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_740_cse <= (result_rem_11cyc_st_4(3)) AND asn_itm_4 AND main_stage_0_5;
  nor_424_nl <= NOT(and_740_cse OR and_dcpl_122);
  or_852_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      and_dcpl_105);
  mux_tmp_314 <= MUX_s_1_2_2(nor_424_nl, or_852_nl, or_850_cse);
  nand_55_cse <= NOT((result_rem_11cyc_st_3(3)) AND asn_itm_3 AND main_stage_0_4);
  and_741_nl <= nand_55_cse AND mux_tmp_314;
  mux_tmp_315 <= MUX_s_1_2_2(and_741_nl, mux_tmp_314, or_839_cse);
  and_742_nl <= nand_58_cse AND mux_tmp_315;
  mux_tmp_316 <= MUX_s_1_2_2(and_742_nl, mux_tmp_315, or_830_cse);
  and_743_nl <= not_tmp_645 AND mux_tmp_316;
  mux_tmp_317 <= MUX_s_1_2_2(and_743_nl, mux_tmp_316, or_823_cse);
  nor_423_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_317));
  mux_318_nl <= MUX_s_1_2_2(nor_423_nl, mux_tmp_317, or_818_cse);
  and_dcpl_549 <= mux_318_nl AND and_dcpl_100;
  or_863_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1000"));
  nor_422_nl <= NOT(and_dcpl_105 OR and_dcpl_100);
  or_865_nl <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_99);
  mux_tmp_319 <= MUX_s_1_2_2(nor_422_nl, or_865_nl, or_863_cse);
  nand_51_cse <= NOT((result_rem_11cyc_st_4(3)) AND asn_itm_4 AND main_stage_0_5);
  and_736_nl <= nand_51_cse AND mux_tmp_319;
  mux_tmp_320 <= MUX_s_1_2_2(and_736_nl, mux_tmp_319, or_850_cse);
  and_737_nl <= nand_55_cse AND mux_tmp_320;
  mux_tmp_321 <= MUX_s_1_2_2(and_737_nl, mux_tmp_320, or_839_cse);
  and_738_nl <= nand_58_cse AND mux_tmp_321;
  mux_tmp_322 <= MUX_s_1_2_2(and_738_nl, mux_tmp_321, or_830_cse);
  and_739_nl <= not_tmp_645 AND mux_tmp_322;
  mux_tmp_323 <= MUX_s_1_2_2(and_739_nl, mux_tmp_322, or_823_cse);
  nor_421_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_323));
  mux_324_nl <= MUX_s_1_2_2(nor_421_nl, mux_tmp_323, or_818_cse);
  and_dcpl_552 <= mux_324_nl AND and_dcpl_74;
  or_878_cse <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_731_cse <= (result_rem_11cyc_st_6(3)) AND asn_itm_6 AND main_stage_0_7;
  nor_419_nl <= NOT(and_731_cse OR and_dcpl_74);
  or_880_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_73);
  mux_tmp_325 <= MUX_s_1_2_2(nor_419_nl, or_880_nl, or_878_cse);
  nor_420_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_325));
  mux_tmp_326 <= MUX_s_1_2_2(nor_420_nl, mux_tmp_325, or_863_cse);
  and_732_nl <= nand_51_cse AND mux_tmp_326;
  mux_tmp_327 <= MUX_s_1_2_2(and_732_nl, mux_tmp_326, or_850_cse);
  and_733_nl <= nand_55_cse AND mux_tmp_327;
  mux_tmp_328 <= MUX_s_1_2_2(and_733_nl, mux_tmp_327, or_839_cse);
  and_734_nl <= nand_58_cse AND mux_tmp_328;
  mux_tmp_329 <= MUX_s_1_2_2(and_734_nl, mux_tmp_328, or_830_cse);
  and_735_nl <= not_tmp_645 AND mux_tmp_329;
  mux_tmp_330 <= MUX_s_1_2_2(and_735_nl, mux_tmp_329, or_823_cse);
  nor_418_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_330));
  mux_331_nl <= MUX_s_1_2_2(nor_418_nl, mux_tmp_330, or_818_cse);
  and_dcpl_556 <= mux_331_nl AND and_dcpl_45;
  and_725_cse <= (result_rem_11cyc_st_7(3)) AND asn_itm_7 AND main_stage_0_8;
  nor_415_nl <= NOT(and_725_cse OR and_dcpl_45);
  or_897_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      and_dcpl_28);
  or_895_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_332 <= MUX_s_1_2_2(nor_415_nl, or_897_nl, or_895_nl);
  nand_42_cse <= NOT((result_rem_11cyc_st_6(3)) AND asn_itm_6 AND main_stage_0_7);
  and_726_nl <= nand_42_cse AND mux_tmp_332;
  mux_tmp_333 <= MUX_s_1_2_2(and_726_nl, mux_tmp_332, or_878_cse);
  nor_416_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_333));
  mux_tmp_334 <= MUX_s_1_2_2(nor_416_nl, mux_tmp_333, or_863_cse);
  and_727_nl <= nand_51_cse AND mux_tmp_334;
  mux_tmp_335 <= MUX_s_1_2_2(and_727_nl, mux_tmp_334, or_850_cse);
  and_728_nl <= nand_55_cse AND mux_tmp_335;
  mux_tmp_336 <= MUX_s_1_2_2(and_728_nl, mux_tmp_335, or_839_cse);
  and_729_nl <= nand_58_cse AND mux_tmp_336;
  mux_tmp_337 <= MUX_s_1_2_2(and_729_nl, mux_tmp_336, or_830_cse);
  and_730_nl <= not_tmp_645 AND mux_tmp_337;
  mux_tmp_338 <= MUX_s_1_2_2(and_730_nl, mux_tmp_337, or_823_cse);
  nor_417_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_338));
  mux_339_nl <= MUX_s_1_2_2(nor_417_nl, mux_tmp_338, or_818_cse);
  and_dcpl_560 <= mux_339_nl AND and_dcpl_4 AND and_dcpl_18 AND (NOT (result_rem_11cyc_st_9(0)));
  or_tmp_897 <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("1000"));
  nor_407_nl <= NOT((result_rem_11cyc_st_8(3)) OR (NOT or_tmp_897));
  or_914_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_340 <= MUX_s_1_2_2(nor_407_nl, or_tmp_897, or_914_nl);
  nor_408_nl <= NOT((result_rem_11cyc_st_7(3)) OR (NOT mux_tmp_340));
  or_913_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_341 <= MUX_s_1_2_2(nor_408_nl, mux_tmp_340, or_913_nl);
  nor_409_nl <= NOT((result_rem_11cyc_st_6(3)) OR (NOT mux_tmp_341));
  or_912_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_342 <= MUX_s_1_2_2(nor_409_nl, mux_tmp_341, or_912_nl);
  nor_410_nl <= NOT((result_rem_11cyc_st_5(3)) OR (NOT mux_tmp_342));
  or_911_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_343 <= MUX_s_1_2_2(nor_410_nl, mux_tmp_342, or_911_nl);
  nor_411_nl <= NOT((result_rem_11cyc_st_4(3)) OR (NOT mux_tmp_343));
  or_910_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_344 <= MUX_s_1_2_2(nor_411_nl, mux_tmp_343, or_910_nl);
  nor_412_nl <= NOT((result_rem_11cyc_st_3(3)) OR (NOT mux_tmp_344));
  or_909_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_345 <= MUX_s_1_2_2(nor_412_nl, mux_tmp_344, or_909_nl);
  nor_413_nl <= NOT((result_rem_11cyc_st_2(3)) OR (NOT mux_tmp_345));
  or_908_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_346 <= MUX_s_1_2_2(nor_413_nl, mux_tmp_345, or_908_nl);
  and_724_nl <= not_tmp_645 AND mux_tmp_346;
  mux_tmp_347 <= MUX_s_1_2_2(and_724_nl, mux_tmp_346, or_823_cse);
  nor_414_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_347));
  mux_tmp_348 <= MUX_s_1_2_2(nor_414_nl, mux_tmp_347, or_818_cse);
  and_dcpl_566 <= and_dcpl_532 AND and_dcpl_318;
  or_tmp_909 <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR not_tmp_645;
  or_928_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("1001"));
  nor_406_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_909));
  mux_349_nl <= MUX_s_1_2_2(nor_406_nl, or_tmp_909, or_928_cse);
  and_dcpl_568 <= mux_349_nl AND and_dcpl_204;
  or_933_cse <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_405_nl <= NOT(and_749_cse OR and_dcpl_204);
  or_935_nl <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_202);
  mux_tmp_350 <= MUX_s_1_2_2(nor_405_nl, or_935_nl, or_933_cse);
  nor_404_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_350));
  mux_351_nl <= MUX_s_1_2_2(nor_404_nl, mux_tmp_350, or_928_cse);
  and_dcpl_570 <= mux_351_nl AND and_dcpl_178;
  or_940_cse <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_403_nl <= NOT(and_747_cse OR and_dcpl_178);
  or_942_nl <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_176);
  mux_tmp_352 <= MUX_s_1_2_2(nor_403_nl, or_942_nl, or_940_cse);
  and_722_nl <= not_tmp_645 AND mux_tmp_352;
  mux_tmp_353 <= MUX_s_1_2_2(and_722_nl, mux_tmp_352, or_933_cse);
  nor_402_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_353));
  mux_354_nl <= MUX_s_1_2_2(nor_402_nl, mux_tmp_353, or_928_cse);
  and_dcpl_572 <= mux_354_nl AND and_dcpl_152;
  or_949_cse <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_401_nl <= NOT(and_744_cse OR and_dcpl_152);
  or_951_nl <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_150);
  mux_tmp_355 <= MUX_s_1_2_2(nor_401_nl, or_951_nl, or_949_cse);
  and_719_nl <= nand_58_cse AND mux_tmp_355;
  mux_tmp_356 <= MUX_s_1_2_2(and_719_nl, mux_tmp_355, or_940_cse);
  and_720_nl <= not_tmp_645 AND mux_tmp_356;
  mux_tmp_357 <= MUX_s_1_2_2(and_720_nl, mux_tmp_356, or_933_cse);
  nor_400_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_357));
  mux_358_nl <= MUX_s_1_2_2(nor_400_nl, mux_tmp_357, or_928_cse);
  and_dcpl_576 <= mux_358_nl AND and_dcpl_125;
  or_960_cse <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_399_nl <= NOT(and_740_cse OR and_dcpl_125);
  or_962_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1001")) OR (NOT
      and_dcpl_105);
  mux_tmp_359 <= MUX_s_1_2_2(nor_399_nl, or_962_nl, or_960_cse);
  and_715_nl <= nand_55_cse AND mux_tmp_359;
  mux_tmp_360 <= MUX_s_1_2_2(and_715_nl, mux_tmp_359, or_949_cse);
  and_716_nl <= nand_58_cse AND mux_tmp_360;
  mux_tmp_361 <= MUX_s_1_2_2(and_716_nl, mux_tmp_360, or_940_cse);
  and_717_nl <= not_tmp_645 AND mux_tmp_361;
  mux_tmp_362 <= MUX_s_1_2_2(and_717_nl, mux_tmp_361, or_933_cse);
  nor_398_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_362));
  mux_363_nl <= MUX_s_1_2_2(nor_398_nl, mux_tmp_362, or_928_cse);
  and_dcpl_578 <= mux_363_nl AND and_dcpl_101;
  or_973_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1001"));
  nor_397_nl <= NOT(and_dcpl_105 OR and_dcpl_101);
  or_975_nl <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_99);
  mux_tmp_364 <= MUX_s_1_2_2(nor_397_nl, or_975_nl, or_973_cse);
  and_710_nl <= nand_51_cse AND mux_tmp_364;
  mux_tmp_365 <= MUX_s_1_2_2(and_710_nl, mux_tmp_364, or_960_cse);
  and_711_nl <= nand_55_cse AND mux_tmp_365;
  mux_tmp_366 <= MUX_s_1_2_2(and_711_nl, mux_tmp_365, or_949_cse);
  and_712_nl <= nand_58_cse AND mux_tmp_366;
  mux_tmp_367 <= MUX_s_1_2_2(and_712_nl, mux_tmp_366, or_940_cse);
  and_713_nl <= not_tmp_645 AND mux_tmp_367;
  mux_tmp_368 <= MUX_s_1_2_2(and_713_nl, mux_tmp_367, or_933_cse);
  nor_396_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_368));
  mux_369_nl <= MUX_s_1_2_2(nor_396_nl, mux_tmp_368, or_928_cse);
  and_dcpl_580 <= mux_369_nl AND and_dcpl_75;
  or_988_cse <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_394_nl <= NOT(and_731_cse OR and_dcpl_75);
  or_990_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_73);
  mux_tmp_370 <= MUX_s_1_2_2(nor_394_nl, or_990_nl, or_988_cse);
  nor_395_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_370));
  mux_tmp_371 <= MUX_s_1_2_2(nor_395_nl, mux_tmp_370, or_973_cse);
  and_706_nl <= nand_51_cse AND mux_tmp_371;
  mux_tmp_372 <= MUX_s_1_2_2(and_706_nl, mux_tmp_371, or_960_cse);
  and_707_nl <= nand_55_cse AND mux_tmp_372;
  mux_tmp_373 <= MUX_s_1_2_2(and_707_nl, mux_tmp_372, or_949_cse);
  and_708_nl <= nand_58_cse AND mux_tmp_373;
  mux_tmp_374 <= MUX_s_1_2_2(and_708_nl, mux_tmp_373, or_940_cse);
  and_709_nl <= not_tmp_645 AND mux_tmp_374;
  mux_tmp_375 <= MUX_s_1_2_2(and_709_nl, mux_tmp_374, or_933_cse);
  nor_393_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_375));
  mux_376_nl <= MUX_s_1_2_2(nor_393_nl, mux_tmp_375, or_928_cse);
  and_dcpl_583 <= mux_376_nl AND and_dcpl_47;
  nor_390_nl <= NOT(and_725_cse OR and_dcpl_47);
  or_1007_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("1001")) OR
      (NOT and_dcpl_28);
  or_1005_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_377 <= MUX_s_1_2_2(nor_390_nl, or_1007_nl, or_1005_nl);
  and_700_nl <= nand_42_cse AND mux_tmp_377;
  mux_tmp_378 <= MUX_s_1_2_2(and_700_nl, mux_tmp_377, or_988_cse);
  nor_391_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_378));
  mux_tmp_379 <= MUX_s_1_2_2(nor_391_nl, mux_tmp_378, or_973_cse);
  and_701_nl <= nand_51_cse AND mux_tmp_379;
  mux_tmp_380 <= MUX_s_1_2_2(and_701_nl, mux_tmp_379, or_960_cse);
  and_702_nl <= nand_55_cse AND mux_tmp_380;
  mux_tmp_381 <= MUX_s_1_2_2(and_702_nl, mux_tmp_380, or_949_cse);
  and_703_nl <= nand_58_cse AND mux_tmp_381;
  mux_tmp_382 <= MUX_s_1_2_2(and_703_nl, mux_tmp_381, or_940_cse);
  and_704_nl <= not_tmp_645 AND mux_tmp_382;
  mux_tmp_383 <= MUX_s_1_2_2(and_704_nl, mux_tmp_382, or_933_cse);
  nor_392_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_383));
  mux_384_nl <= MUX_s_1_2_2(nor_392_nl, mux_tmp_383, or_928_cse);
  and_dcpl_586 <= mux_384_nl AND and_dcpl_4 AND and_dcpl_18 AND (result_rem_11cyc_st_9(0));
  or_tmp_1005 <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("1001"));
  nor_383_nl <= NOT((result_rem_11cyc_st_8(3)) OR (NOT or_tmp_1005));
  or_1024_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_385 <= MUX_s_1_2_2(nor_383_nl, or_tmp_1005, or_1024_nl);
  nor_384_nl <= NOT((result_rem_11cyc_st_7(3)) OR (NOT mux_tmp_385));
  or_1023_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_386 <= MUX_s_1_2_2(nor_384_nl, mux_tmp_385, or_1023_nl);
  nor_385_nl <= NOT((result_rem_11cyc_st_6(3)) OR (NOT mux_tmp_386));
  or_1022_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_387 <= MUX_s_1_2_2(nor_385_nl, mux_tmp_386, or_1022_nl);
  nor_386_nl <= NOT((result_rem_11cyc_st_5(3)) OR (NOT mux_tmp_387));
  or_1021_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_388 <= MUX_s_1_2_2(nor_386_nl, mux_tmp_387, or_1021_nl);
  nor_387_nl <= NOT((result_rem_11cyc_st_4(3)) OR (NOT mux_tmp_388));
  or_1020_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_389 <= MUX_s_1_2_2(nor_387_nl, mux_tmp_388, or_1020_nl);
  nor_388_nl <= NOT((result_rem_11cyc_st_3(3)) OR (NOT mux_tmp_389));
  or_1019_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_390 <= MUX_s_1_2_2(nor_388_nl, mux_tmp_389, or_1019_nl);
  nor_389_nl <= NOT((result_rem_11cyc_st_2(3)) OR (NOT mux_tmp_390));
  or_1018_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_391 <= MUX_s_1_2_2(nor_389_nl, mux_tmp_390, or_1018_nl);
  and_697_nl <= not_tmp_645 AND mux_tmp_391;
  mux_tmp_392 <= MUX_s_1_2_2(and_697_nl, mux_tmp_391, or_933_cse);
  and_698_nl <= nand_146_cse AND mux_tmp_392;
  or_1016_nl <= CONV_SL_1_1(result_result_acc_tmp(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_393 <= MUX_s_1_2_2(and_698_nl, mux_tmp_392, or_1016_nl);
  and_dcpl_590 <= and_dcpl_532 AND and_dcpl_352;
  or_tmp_1017 <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR not_tmp_645;
  or_1037_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("1010"));
  nor_382_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_1017));
  mux_394_nl <= MUX_s_1_2_2(nor_382_nl, or_tmp_1017, or_1037_cse);
  and_dcpl_592 <= mux_394_nl AND and_dcpl_205;
  or_1042_cse <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_381_nl <= NOT(and_749_cse OR and_dcpl_205);
  or_1044_nl <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_202);
  mux_tmp_395 <= MUX_s_1_2_2(nor_381_nl, or_1044_nl, or_1042_cse);
  nor_380_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_395));
  mux_396_nl <= MUX_s_1_2_2(nor_380_nl, mux_tmp_395, or_1037_cse);
  and_dcpl_594 <= mux_396_nl AND and_dcpl_179;
  or_1049_cse <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_379_nl <= NOT(and_747_cse OR and_dcpl_179);
  or_1051_nl <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_176);
  mux_tmp_397 <= MUX_s_1_2_2(nor_379_nl, or_1051_nl, or_1049_cse);
  and_695_nl <= not_tmp_645 AND mux_tmp_397;
  mux_tmp_398 <= MUX_s_1_2_2(and_695_nl, mux_tmp_397, or_1042_cse);
  nor_378_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_398));
  mux_399_nl <= MUX_s_1_2_2(nor_378_nl, mux_tmp_398, or_1037_cse);
  and_dcpl_596 <= mux_399_nl AND and_dcpl_153;
  or_1058_cse <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_377_nl <= NOT(and_744_cse OR and_dcpl_153);
  or_1060_nl <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_150);
  mux_tmp_400 <= MUX_s_1_2_2(nor_377_nl, or_1060_nl, or_1058_cse);
  and_692_nl <= nand_58_cse AND mux_tmp_400;
  mux_tmp_401 <= MUX_s_1_2_2(and_692_nl, mux_tmp_400, or_1049_cse);
  and_693_nl <= not_tmp_645 AND mux_tmp_401;
  mux_tmp_402 <= MUX_s_1_2_2(and_693_nl, mux_tmp_401, or_1042_cse);
  nor_376_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_402));
  mux_403_nl <= MUX_s_1_2_2(nor_376_nl, mux_tmp_402, or_1037_cse);
  and_dcpl_599 <= mux_403_nl AND and_dcpl_127;
  or_1069_cse <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_375_nl <= NOT(and_740_cse OR and_dcpl_127);
  or_1071_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1010")) OR
      (NOT and_dcpl_105);
  mux_tmp_404 <= MUX_s_1_2_2(nor_375_nl, or_1071_nl, or_1069_cse);
  and_688_nl <= nand_55_cse AND mux_tmp_404;
  mux_tmp_405 <= MUX_s_1_2_2(and_688_nl, mux_tmp_404, or_1058_cse);
  and_689_nl <= nand_58_cse AND mux_tmp_405;
  mux_tmp_406 <= MUX_s_1_2_2(and_689_nl, mux_tmp_405, or_1049_cse);
  and_690_nl <= not_tmp_645 AND mux_tmp_406;
  mux_tmp_407 <= MUX_s_1_2_2(and_690_nl, mux_tmp_406, or_1042_cse);
  nor_374_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_407));
  mux_408_nl <= MUX_s_1_2_2(nor_374_nl, mux_tmp_407, or_1037_cse);
  and_dcpl_601 <= mux_408_nl AND and_dcpl_102;
  or_1082_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1010"));
  nor_373_nl <= NOT(and_dcpl_105 OR and_dcpl_102);
  or_1084_nl <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_99);
  mux_tmp_409 <= MUX_s_1_2_2(nor_373_nl, or_1084_nl, or_1082_cse);
  and_683_nl <= nand_51_cse AND mux_tmp_409;
  mux_tmp_410 <= MUX_s_1_2_2(and_683_nl, mux_tmp_409, or_1069_cse);
  and_684_nl <= nand_55_cse AND mux_tmp_410;
  mux_tmp_411 <= MUX_s_1_2_2(and_684_nl, mux_tmp_410, or_1058_cse);
  and_685_nl <= nand_58_cse AND mux_tmp_411;
  mux_tmp_412 <= MUX_s_1_2_2(and_685_nl, mux_tmp_411, or_1049_cse);
  and_686_nl <= not_tmp_645 AND mux_tmp_412;
  mux_tmp_413 <= MUX_s_1_2_2(and_686_nl, mux_tmp_412, or_1042_cse);
  nor_372_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_413));
  mux_414_nl <= MUX_s_1_2_2(nor_372_nl, mux_tmp_413, or_1037_cse);
  and_dcpl_603 <= mux_414_nl AND and_dcpl_76;
  or_1097_cse <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_370_nl <= NOT(and_731_cse OR and_dcpl_76);
  or_1099_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_73);
  mux_tmp_415 <= MUX_s_1_2_2(nor_370_nl, or_1099_nl, or_1097_cse);
  nor_371_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_415));
  mux_tmp_416 <= MUX_s_1_2_2(nor_371_nl, mux_tmp_415, or_1082_cse);
  and_679_nl <= nand_51_cse AND mux_tmp_416;
  mux_tmp_417 <= MUX_s_1_2_2(and_679_nl, mux_tmp_416, or_1069_cse);
  and_680_nl <= nand_55_cse AND mux_tmp_417;
  mux_tmp_418 <= MUX_s_1_2_2(and_680_nl, mux_tmp_417, or_1058_cse);
  and_681_nl <= nand_58_cse AND mux_tmp_418;
  mux_tmp_419 <= MUX_s_1_2_2(and_681_nl, mux_tmp_418, or_1049_cse);
  and_682_nl <= not_tmp_645 AND mux_tmp_419;
  mux_tmp_420 <= MUX_s_1_2_2(and_682_nl, mux_tmp_419, or_1042_cse);
  nor_369_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_420));
  mux_421_nl <= MUX_s_1_2_2(nor_369_nl, mux_tmp_420, or_1037_cse);
  and_dcpl_607 <= mux_421_nl AND and_dcpl_50;
  nor_366_nl <= NOT(and_725_cse OR and_dcpl_50);
  or_1116_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("1010")) OR
      (NOT and_dcpl_28);
  or_1114_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_422 <= MUX_s_1_2_2(nor_366_nl, or_1116_nl, or_1114_nl);
  and_673_nl <= nand_42_cse AND mux_tmp_422;
  mux_tmp_423 <= MUX_s_1_2_2(and_673_nl, mux_tmp_422, or_1097_cse);
  nor_367_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_423));
  mux_tmp_424 <= MUX_s_1_2_2(nor_367_nl, mux_tmp_423, or_1082_cse);
  and_674_nl <= nand_51_cse AND mux_tmp_424;
  mux_tmp_425 <= MUX_s_1_2_2(and_674_nl, mux_tmp_424, or_1069_cse);
  and_675_nl <= nand_55_cse AND mux_tmp_425;
  mux_tmp_426 <= MUX_s_1_2_2(and_675_nl, mux_tmp_425, or_1058_cse);
  and_676_nl <= nand_58_cse AND mux_tmp_426;
  mux_tmp_427 <= MUX_s_1_2_2(and_676_nl, mux_tmp_426, or_1049_cse);
  and_677_nl <= not_tmp_645 AND mux_tmp_427;
  mux_tmp_428 <= MUX_s_1_2_2(and_677_nl, mux_tmp_427, or_1042_cse);
  nor_368_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_428));
  mux_429_nl <= MUX_s_1_2_2(nor_368_nl, mux_tmp_428, or_1037_cse);
  and_dcpl_611 <= mux_429_nl AND and_dcpl_4 AND (result_rem_11cyc_st_9(3)) AND (result_rem_11cyc_st_9(1))
      AND (NOT (result_rem_11cyc_st_9(0)));
  or_tmp_1113 <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("1010"));
  nor_358_nl <= NOT((result_rem_11cyc_st_8(3)) OR (NOT or_tmp_1113));
  or_1133_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_430 <= MUX_s_1_2_2(nor_358_nl, or_tmp_1113, or_1133_nl);
  nor_359_nl <= NOT((result_rem_11cyc_st_7(3)) OR (NOT mux_tmp_430));
  or_1132_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_431 <= MUX_s_1_2_2(nor_359_nl, mux_tmp_430, or_1132_nl);
  nor_360_nl <= NOT((result_rem_11cyc_st_6(3)) OR (NOT mux_tmp_431));
  or_1131_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_432 <= MUX_s_1_2_2(nor_360_nl, mux_tmp_431, or_1131_nl);
  nor_361_nl <= NOT((result_rem_11cyc_st_5(3)) OR (NOT mux_tmp_432));
  or_1130_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_433 <= MUX_s_1_2_2(nor_361_nl, mux_tmp_432, or_1130_nl);
  nor_362_nl <= NOT((result_rem_11cyc_st_4(3)) OR (NOT mux_tmp_433));
  or_1129_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_434 <= MUX_s_1_2_2(nor_362_nl, mux_tmp_433, or_1129_nl);
  nor_363_nl <= NOT((result_rem_11cyc_st_3(3)) OR (NOT mux_tmp_434));
  or_1128_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_435 <= MUX_s_1_2_2(nor_363_nl, mux_tmp_434, or_1128_nl);
  nor_364_nl <= NOT((result_rem_11cyc_st_2(3)) OR (NOT mux_tmp_435));
  or_1127_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_436 <= MUX_s_1_2_2(nor_364_nl, mux_tmp_435, or_1127_nl);
  and_671_nl <= not_tmp_645 AND mux_tmp_436;
  mux_tmp_437 <= MUX_s_1_2_2(and_671_nl, mux_tmp_436, or_1042_cse);
  nor_365_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_437));
  mux_tmp_438 <= MUX_s_1_2_2(nor_365_nl, mux_tmp_437, or_1037_cse);
  return_rsci_d_mx0c0 <= and_dcpl_235 AND and_dcpl_233;
  return_rsci_d_mx0c1 <= and_dcpl_235 AND and_dcpl_237;
  return_rsci_d_mx0c2 <= and_dcpl_235 AND and_dcpl_240;
  return_rsci_d_mx0c3 <= and_dcpl_235 AND and_dcpl_239 AND (result_rem_11cyc_st_11(0));
  return_rsci_d_mx0c4 <= and_dcpl_235 AND and_dcpl_244 AND (NOT (result_rem_11cyc_st_11(0)));
  return_rsci_d_mx0c5 <= and_dcpl_235 AND and_dcpl_244 AND (result_rem_11cyc_st_11(0));
  return_rsci_d_mx0c6 <= and_dcpl_235 AND and_dcpl_249 AND (NOT (result_rem_11cyc_st_11(0)));
  return_rsci_d_mx0c7 <= and_dcpl_235 AND and_dcpl_249 AND (result_rem_11cyc_st_11(0));
  return_rsci_d_mx0c8 <= and_dcpl_254 AND and_dcpl_233;
  return_rsci_d_mx0c9 <= and_dcpl_254 AND and_dcpl_237;
  return_rsci_d_mx0c10 <= and_dcpl_254 AND and_dcpl_240;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( (ccs_ccore_en AND (return_rsci_d_mx0c0 OR return_rsci_d_mx0c1 OR return_rsci_d_mx0c2
          OR return_rsci_d_mx0c3 OR return_rsci_d_mx0c4 OR return_rsci_d_mx0c5 OR
          return_rsci_d_mx0c6 OR return_rsci_d_mx0c7 OR return_rsci_d_mx0c8 OR return_rsci_d_mx0c9
          OR return_rsci_d_mx0c10)) = '1' ) THEN
        return_rsci_d <= MUX1HOT_v_64_11_2(result_rem_12_cmp_1_z, result_rem_12_cmp_2_z,
            result_rem_12_cmp_3_z, result_rem_12_cmp_4_z, result_rem_12_cmp_5_z,
            result_rem_12_cmp_6_z, result_rem_12_cmp_7_z, result_rem_12_cmp_8_z,
            result_rem_12_cmp_9_z, result_rem_12_cmp_10_z, result_rem_12_cmp_z, STD_LOGIC_VECTOR'(
            return_rsci_d_mx0c0 & return_rsci_d_mx0c1 & return_rsci_d_mx0c2 & return_rsci_d_mx0c3
            & return_rsci_d_mx0c4 & return_rsci_d_mx0c5 & return_rsci_d_mx0c6 & return_rsci_d_mx0c7
            & return_rsci_d_mx0c8 & return_rsci_d_mx0c9 & return_rsci_d_mx0c10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_11 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND main_stage_0_11 AND asn_itm_10) = '1' ) THEN
        result_rem_11cyc_st_11 <= result_rem_11cyc_st_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        asn_itm_11 <= '0';
        asn_itm_10 <= '0';
        asn_itm_9 <= '0';
        asn_itm_8 <= '0';
        asn_itm_7 <= '0';
        asn_itm_6 <= '0';
        asn_itm_5 <= '0';
        asn_itm_4 <= '0';
        asn_itm_3 <= '0';
        asn_itm_2 <= '0';
        asn_itm_1 <= '0';
        main_stage_0_2 <= '0';
        main_stage_0_3 <= '0';
        main_stage_0_4 <= '0';
        main_stage_0_5 <= '0';
        main_stage_0_6 <= '0';
        main_stage_0_7 <= '0';
        main_stage_0_8 <= '0';
        main_stage_0_9 <= '0';
        main_stage_0_10 <= '0';
        main_stage_0_11 <= '0';
        main_stage_0_12 <= '0';
      ELSIF ( ccs_ccore_en = '1' ) THEN
        asn_itm_11 <= asn_itm_10;
        asn_itm_10 <= asn_itm_9;
        asn_itm_9 <= asn_itm_8;
        asn_itm_8 <= asn_itm_7;
        asn_itm_7 <= asn_itm_6;
        asn_itm_6 <= asn_itm_5;
        asn_itm_5 <= asn_itm_4;
        asn_itm_4 <= asn_itm_3;
        asn_itm_3 <= asn_itm_2;
        asn_itm_2 <= asn_itm_1;
        asn_itm_1 <= ccs_ccore_start_rsci_idat;
        main_stage_0_2 <= '1';
        main_stage_0_3 <= main_stage_0_2;
        main_stage_0_4 <= main_stage_0_3;
        main_stage_0_5 <= main_stage_0_4;
        main_stage_0_6 <= main_stage_0_5;
        main_stage_0_7 <= main_stage_0_6;
        main_stage_0_8 <= main_stage_0_7;
        main_stage_0_9 <= main_stage_0_8;
        main_stage_0_10 <= main_stage_0_9;
        main_stage_0_11 <= main_stage_0_10;
        main_stage_0_12 <= main_stage_0_11;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_1_cse = '1' ) THEN
        result_rem_12_cmp_1_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_1_2,
            m_buf_sva_mut_1_3, m_buf_sva_mut_1_4, m_buf_sva_mut_1_5, m_buf_sva_mut_1_6,
            m_buf_sva_mut_1_7, m_buf_sva_mut_1_8, m_buf_sva_mut_1_9, m_buf_sva_mut_1_10,
            STD_LOGIC_VECTOR'( and_dcpl_263 & and_dcpl_269 & and_dcpl_275 & and_dcpl_281
            & and_dcpl_287 & and_dcpl_293 & and_dcpl_299 & and_dcpl_305 & and_dcpl_311
            & mux_tmp_37));
        result_rem_12_cmp_1_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_1_2,
            base_buf_sva_mut_1_3, base_buf_sva_mut_1_4, base_buf_sva_mut_1_5, base_buf_sva_mut_1_6,
            base_buf_sva_mut_1_7, base_buf_sva_mut_1_8, base_buf_sva_mut_1_9, base_buf_sva_mut_1_10,
            STD_LOGIC_VECTOR'( and_dcpl_263 & and_dcpl_269 & and_dcpl_275 & and_dcpl_281
            & and_dcpl_287 & and_dcpl_293 & and_dcpl_299 & and_dcpl_305 & and_dcpl_311
            & mux_tmp_37));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_3_cse = '1' ) THEN
        result_rem_12_cmp_2_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_2_2,
            m_buf_sva_mut_2_3, m_buf_sva_mut_2_4, m_buf_sva_mut_2_5, m_buf_sva_mut_2_6,
            m_buf_sva_mut_2_7, m_buf_sva_mut_2_8, m_buf_sva_mut_2_9, m_buf_sva_mut_2_10,
            STD_LOGIC_VECTOR'( and_dcpl_319 & and_dcpl_322 & and_dcpl_325 & and_dcpl_329
            & and_dcpl_333 & and_dcpl_337 & and_dcpl_341 & and_dcpl_344 & and_dcpl_347
            & mux_tmp_75));
        result_rem_12_cmp_2_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_2_2,
            base_buf_sva_mut_2_3, base_buf_sva_mut_2_4, base_buf_sva_mut_2_5, base_buf_sva_mut_2_6,
            base_buf_sva_mut_2_7, base_buf_sva_mut_2_8, base_buf_sva_mut_2_9, base_buf_sva_mut_2_10,
            STD_LOGIC_VECTOR'( and_dcpl_319 & and_dcpl_322 & and_dcpl_325 & and_dcpl_329
            & and_dcpl_333 & and_dcpl_337 & and_dcpl_341 & and_dcpl_344 & and_dcpl_347
            & mux_tmp_75));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_5_cse = '1' ) THEN
        result_rem_12_cmp_3_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_3_2,
            m_buf_sva_mut_3_3, m_buf_sva_mut_3_4, m_buf_sva_mut_3_5, m_buf_sva_mut_3_6,
            m_buf_sva_mut_3_7, m_buf_sva_mut_3_8, m_buf_sva_mut_3_9, m_buf_sva_mut_3_10,
            STD_LOGIC_VECTOR'( and_dcpl_353 & and_dcpl_357 & and_dcpl_361 & and_dcpl_364
            & and_dcpl_367 & and_dcpl_370 & and_dcpl_373 & and_dcpl_377 & and_dcpl_381
            & mux_tmp_113));
        result_rem_12_cmp_3_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_3_2,
            base_buf_sva_mut_3_3, base_buf_sva_mut_3_4, base_buf_sva_mut_3_5, base_buf_sva_mut_3_6,
            base_buf_sva_mut_3_7, base_buf_sva_mut_3_8, base_buf_sva_mut_3_9, base_buf_sva_mut_3_10,
            STD_LOGIC_VECTOR'( and_dcpl_353 & and_dcpl_357 & and_dcpl_361 & and_dcpl_364
            & and_dcpl_367 & and_dcpl_370 & and_dcpl_373 & and_dcpl_377 & and_dcpl_381
            & mux_tmp_113));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_7_cse = '1' ) THEN
        result_rem_12_cmp_4_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_4_2,
            m_buf_sva_mut_4_3, m_buf_sva_mut_4_4, m_buf_sva_mut_4_5, m_buf_sva_mut_4_6,
            m_buf_sva_mut_4_7, m_buf_sva_mut_4_8, m_buf_sva_mut_4_9, m_buf_sva_mut_4_10,
            STD_LOGIC_VECTOR'( and_dcpl_387 & and_dcpl_390 & and_dcpl_393 & and_dcpl_396
            & and_dcpl_399 & and_dcpl_402 & and_dcpl_405 & and_dcpl_408 & and_dcpl_411
            & mux_tmp_151));
        result_rem_12_cmp_4_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_4_2,
            base_buf_sva_mut_4_3, base_buf_sva_mut_4_4, base_buf_sva_mut_4_5, base_buf_sva_mut_4_6,
            base_buf_sva_mut_4_7, base_buf_sva_mut_4_8, base_buf_sva_mut_4_9, base_buf_sva_mut_4_10,
            STD_LOGIC_VECTOR'( and_dcpl_387 & and_dcpl_390 & and_dcpl_393 & and_dcpl_396
            & and_dcpl_399 & and_dcpl_402 & and_dcpl_405 & and_dcpl_408 & and_dcpl_411
            & mux_tmp_151));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_9_cse = '1' ) THEN
        result_rem_12_cmp_5_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_5_2,
            m_buf_sva_mut_5_3, m_buf_sva_mut_5_4, m_buf_sva_mut_5_5, m_buf_sva_mut_5_6,
            m_buf_sva_mut_5_7, m_buf_sva_mut_5_8, m_buf_sva_mut_5_9, m_buf_sva_mut_5_10,
            STD_LOGIC_VECTOR'( and_dcpl_418 & and_dcpl_422 & and_dcpl_426 & and_dcpl_430
            & and_dcpl_433 & and_dcpl_437 & and_dcpl_441 & and_dcpl_444 & and_dcpl_447
            & mux_tmp_189));
        result_rem_12_cmp_5_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_5_2,
            base_buf_sva_mut_5_3, base_buf_sva_mut_5_4, base_buf_sva_mut_5_5, base_buf_sva_mut_5_6,
            base_buf_sva_mut_5_7, base_buf_sva_mut_5_8, base_buf_sva_mut_5_9, base_buf_sva_mut_5_10,
            STD_LOGIC_VECTOR'( and_dcpl_418 & and_dcpl_422 & and_dcpl_426 & and_dcpl_430
            & and_dcpl_433 & and_dcpl_437 & and_dcpl_441 & and_dcpl_444 & and_dcpl_447
            & mux_tmp_189));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_11_cse = '1' ) THEN
        result_rem_12_cmp_6_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_6_2,
            m_buf_sva_mut_6_3, m_buf_sva_mut_6_4, m_buf_sva_mut_6_5, m_buf_sva_mut_6_6,
            m_buf_sva_mut_6_7, m_buf_sva_mut_6_8, m_buf_sva_mut_6_9, m_buf_sva_mut_6_10,
            STD_LOGIC_VECTOR'( and_dcpl_452 & and_dcpl_455 & and_dcpl_458 & and_dcpl_462
            & and_dcpl_464 & and_dcpl_468 & and_dcpl_472 & and_dcpl_474 & and_dcpl_476
            & mux_tmp_227));
        result_rem_12_cmp_6_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_6_2,
            base_buf_sva_mut_6_3, base_buf_sva_mut_6_4, base_buf_sva_mut_6_5, base_buf_sva_mut_6_6,
            base_buf_sva_mut_6_7, base_buf_sva_mut_6_8, base_buf_sva_mut_6_9, base_buf_sva_mut_6_10,
            STD_LOGIC_VECTOR'( and_dcpl_452 & and_dcpl_455 & and_dcpl_458 & and_dcpl_462
            & and_dcpl_464 & and_dcpl_468 & and_dcpl_472 & and_dcpl_474 & and_dcpl_476
            & mux_tmp_227));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_13_cse = '1' ) THEN
        result_rem_12_cmp_7_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_7_2,
            m_buf_sva_mut_7_3, m_buf_sva_mut_7_4, m_buf_sva_mut_7_5, m_buf_sva_mut_7_6,
            m_buf_sva_mut_7_7, m_buf_sva_mut_7_8, m_buf_sva_mut_7_9, m_buf_sva_mut_7_10,
            STD_LOGIC_VECTOR'( and_dcpl_480 & and_dcpl_484 & and_dcpl_488 & and_dcpl_491
            & and_dcpl_493 & and_dcpl_496 & and_dcpl_499 & and_dcpl_501 & and_dcpl_503
            & mux_tmp_265));
        result_rem_12_cmp_7_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_7_2,
            base_buf_sva_mut_7_3, base_buf_sva_mut_7_4, base_buf_sva_mut_7_5, base_buf_sva_mut_7_6,
            base_buf_sva_mut_7_7, base_buf_sva_mut_7_8, base_buf_sva_mut_7_9, base_buf_sva_mut_7_10,
            STD_LOGIC_VECTOR'( and_dcpl_480 & and_dcpl_484 & and_dcpl_488 & and_dcpl_491
            & and_dcpl_493 & and_dcpl_496 & and_dcpl_499 & and_dcpl_501 & and_dcpl_503
            & mux_tmp_265));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_15_cse = '1' ) THEN
        result_rem_12_cmp_8_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_8_2,
            m_buf_sva_mut_8_3, m_buf_sva_mut_8_4, m_buf_sva_mut_8_5, m_buf_sva_mut_8_6,
            m_buf_sva_mut_8_7, m_buf_sva_mut_8_8, m_buf_sva_mut_8_9, m_buf_sva_mut_8_10,
            STD_LOGIC_VECTOR'( and_dcpl_507 & and_dcpl_510 & and_dcpl_513 & and_dcpl_516
            & and_dcpl_518 & and_dcpl_521 & and_dcpl_524 & and_dcpl_526 & and_dcpl_528
            & mux_tmp_303));
        result_rem_12_cmp_8_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_8_2,
            base_buf_sva_mut_8_3, base_buf_sva_mut_8_4, base_buf_sva_mut_8_5, base_buf_sva_mut_8_6,
            base_buf_sva_mut_8_7, base_buf_sva_mut_8_8, base_buf_sva_mut_8_9, base_buf_sva_mut_8_10,
            STD_LOGIC_VECTOR'( and_dcpl_507 & and_dcpl_510 & and_dcpl_513 & and_dcpl_516
            & and_dcpl_518 & and_dcpl_521 & and_dcpl_524 & and_dcpl_526 & and_dcpl_528
            & mux_tmp_303));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_17_cse = '1' ) THEN
        result_rem_12_cmp_9_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_9_2,
            m_buf_sva_mut_9_3, m_buf_sva_mut_9_4, m_buf_sva_mut_9_5, m_buf_sva_mut_9_6,
            m_buf_sva_mut_9_7, m_buf_sva_mut_9_8, m_buf_sva_mut_9_9, m_buf_sva_mut_9_10,
            STD_LOGIC_VECTOR'( and_dcpl_533 & and_dcpl_536 & and_dcpl_539 & and_dcpl_542
            & and_dcpl_546 & and_dcpl_549 & and_dcpl_552 & and_dcpl_556 & and_dcpl_560
            & mux_tmp_348));
        result_rem_12_cmp_9_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_9_2,
            base_buf_sva_mut_9_3, base_buf_sva_mut_9_4, base_buf_sva_mut_9_5, base_buf_sva_mut_9_6,
            base_buf_sva_mut_9_7, base_buf_sva_mut_9_8, base_buf_sva_mut_9_9, base_buf_sva_mut_9_10,
            STD_LOGIC_VECTOR'( and_dcpl_533 & and_dcpl_536 & and_dcpl_539 & and_dcpl_542
            & and_dcpl_546 & and_dcpl_549 & and_dcpl_552 & and_dcpl_556 & and_dcpl_560
            & mux_tmp_348));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_19_cse = '1' ) THEN
        result_rem_12_cmp_10_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_10_2,
            m_buf_sva_mut_10_3, m_buf_sva_mut_10_4, m_buf_sva_mut_10_5, m_buf_sva_mut_10_6,
            m_buf_sva_mut_10_7, m_buf_sva_mut_10_8, m_buf_sva_mut_10_9, m_buf_sva_mut_10_10,
            STD_LOGIC_VECTOR'( and_dcpl_566 & and_dcpl_568 & and_dcpl_570 & and_dcpl_572
            & and_dcpl_576 & and_dcpl_578 & and_dcpl_580 & and_dcpl_583 & and_dcpl_586
            & mux_tmp_393));
        result_rem_12_cmp_10_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_10_2,
            base_buf_sva_mut_10_3, base_buf_sva_mut_10_4, base_buf_sva_mut_10_5,
            base_buf_sva_mut_10_6, base_buf_sva_mut_10_7, base_buf_sva_mut_10_8,
            base_buf_sva_mut_10_9, base_buf_sva_mut_10_10, STD_LOGIC_VECTOR'( and_dcpl_566
            & and_dcpl_568 & and_dcpl_570 & and_dcpl_572 & and_dcpl_576 & and_dcpl_578
            & and_dcpl_580 & and_dcpl_583 & and_dcpl_586 & mux_tmp_393));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_21_cse = '1' ) THEN
        result_rem_12_cmp_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_2, m_buf_sva_mut_3,
            m_buf_sva_mut_4, m_buf_sva_mut_5, m_buf_sva_mut_6, m_buf_sva_mut_7, m_buf_sva_mut_8,
            m_buf_sva_mut_9, m_buf_sva_mut_10, STD_LOGIC_VECTOR'( and_dcpl_590 &
            and_dcpl_592 & and_dcpl_594 & and_dcpl_596 & and_dcpl_599 & and_dcpl_601
            & and_dcpl_603 & and_dcpl_607 & and_dcpl_611 & mux_tmp_438));
        result_rem_12_cmp_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_2,
            base_buf_sva_mut_3, base_buf_sva_mut_4, base_buf_sva_mut_5, base_buf_sva_mut_6,
            base_buf_sva_mut_7, base_buf_sva_mut_8, base_buf_sva_mut_9, base_buf_sva_mut_10,
            STD_LOGIC_VECTOR'( and_dcpl_590 & and_dcpl_592 & and_dcpl_594 & and_dcpl_596
            & and_dcpl_599 & and_dcpl_601 & and_dcpl_603 & and_dcpl_607 & and_dcpl_611
            & mux_tmp_438));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_cse = '1' ) THEN
        m_buf_sva_mut_1_10 <= m_buf_sva_mut_1_9;
        base_buf_sva_mut_1_10 <= base_buf_sva_mut_1_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_1_cse = '1' ) THEN
        m_buf_sva_mut_2_10 <= m_buf_sva_mut_2_9;
        base_buf_sva_mut_2_10 <= base_buf_sva_mut_2_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_2_cse = '1' ) THEN
        m_buf_sva_mut_3_10 <= m_buf_sva_mut_3_9;
        base_buf_sva_mut_3_10 <= base_buf_sva_mut_3_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_3_cse = '1' ) THEN
        m_buf_sva_mut_4_10 <= m_buf_sva_mut_4_9;
        base_buf_sva_mut_4_10 <= base_buf_sva_mut_4_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_4_cse = '1' ) THEN
        m_buf_sva_mut_5_10 <= m_buf_sva_mut_5_9;
        base_buf_sva_mut_5_10 <= base_buf_sva_mut_5_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_5_cse = '1' ) THEN
        m_buf_sva_mut_6_10 <= m_buf_sva_mut_6_9;
        base_buf_sva_mut_6_10 <= base_buf_sva_mut_6_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_6_cse = '1' ) THEN
        m_buf_sva_mut_7_10 <= m_buf_sva_mut_7_9;
        base_buf_sva_mut_7_10 <= base_buf_sva_mut_7_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_7_cse = '1' ) THEN
        m_buf_sva_mut_8_10 <= m_buf_sva_mut_8_9;
        base_buf_sva_mut_8_10 <= base_buf_sva_mut_8_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_8_cse = '1' ) THEN
        m_buf_sva_mut_9_10 <= m_buf_sva_mut_9_9;
        base_buf_sva_mut_9_10 <= base_buf_sva_mut_9_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_9_cse = '1' ) THEN
        m_buf_sva_mut_10_10 <= m_buf_sva_mut_10_9;
        base_buf_sva_mut_10_10 <= base_buf_sva_mut_10_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_10_cse = '1' ) THEN
        m_buf_sva_mut_10 <= m_buf_sva_mut_9;
        base_buf_sva_mut_10 <= base_buf_sva_mut_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_10 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_3) = '1' ) THEN
        result_rem_11cyc_st_10 <= result_rem_11cyc_st_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_11_cse = '1' ) THEN
        m_buf_sva_mut_1_9 <= m_buf_sva_mut_1_8;
        base_buf_sva_mut_1_9 <= base_buf_sva_mut_1_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_12_cse = '1' ) THEN
        m_buf_sva_mut_2_9 <= m_buf_sva_mut_2_8;
        base_buf_sva_mut_2_9 <= base_buf_sva_mut_2_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_13_cse = '1' ) THEN
        m_buf_sva_mut_3_9 <= m_buf_sva_mut_3_8;
        base_buf_sva_mut_3_9 <= base_buf_sva_mut_3_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_14_cse = '1' ) THEN
        m_buf_sva_mut_4_9 <= m_buf_sva_mut_4_8;
        base_buf_sva_mut_4_9 <= base_buf_sva_mut_4_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_15_cse = '1' ) THEN
        m_buf_sva_mut_5_9 <= m_buf_sva_mut_5_8;
        base_buf_sva_mut_5_9 <= base_buf_sva_mut_5_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_16_cse = '1' ) THEN
        m_buf_sva_mut_6_9 <= m_buf_sva_mut_6_8;
        base_buf_sva_mut_6_9 <= base_buf_sva_mut_6_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_17_cse = '1' ) THEN
        m_buf_sva_mut_7_9 <= m_buf_sva_mut_7_8;
        base_buf_sva_mut_7_9 <= base_buf_sva_mut_7_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_18_cse = '1' ) THEN
        m_buf_sva_mut_8_9 <= m_buf_sva_mut_8_8;
        base_buf_sva_mut_8_9 <= base_buf_sva_mut_8_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_19_cse = '1' ) THEN
        m_buf_sva_mut_9_9 <= m_buf_sva_mut_9_8;
        base_buf_sva_mut_9_9 <= base_buf_sva_mut_9_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_20_cse = '1' ) THEN
        m_buf_sva_mut_10_9 <= m_buf_sva_mut_10_8;
        base_buf_sva_mut_10_9 <= base_buf_sva_mut_10_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_21_cse = '1' ) THEN
        m_buf_sva_mut_9 <= m_buf_sva_mut_8;
        base_buf_sva_mut_9 <= base_buf_sva_mut_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_9 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_28) = '1' ) THEN
        result_rem_11cyc_st_9 <= result_rem_11cyc_st_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_22_cse = '1' ) THEN
        m_buf_sva_mut_1_8 <= m_buf_sva_mut_1_7;
        base_buf_sva_mut_1_8 <= base_buf_sva_mut_1_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_23_cse = '1' ) THEN
        m_buf_sva_mut_2_8 <= m_buf_sva_mut_2_7;
        base_buf_sva_mut_2_8 <= base_buf_sva_mut_2_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_24_cse = '1' ) THEN
        m_buf_sva_mut_3_8 <= m_buf_sva_mut_3_7;
        base_buf_sva_mut_3_8 <= base_buf_sva_mut_3_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_25_cse = '1' ) THEN
        m_buf_sva_mut_4_8 <= m_buf_sva_mut_4_7;
        base_buf_sva_mut_4_8 <= base_buf_sva_mut_4_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_26_cse = '1' ) THEN
        m_buf_sva_mut_5_8 <= m_buf_sva_mut_5_7;
        base_buf_sva_mut_5_8 <= base_buf_sva_mut_5_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_27_cse = '1' ) THEN
        m_buf_sva_mut_6_8 <= m_buf_sva_mut_6_7;
        base_buf_sva_mut_6_8 <= base_buf_sva_mut_6_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_28_cse = '1' ) THEN
        m_buf_sva_mut_7_8 <= m_buf_sva_mut_7_7;
        base_buf_sva_mut_7_8 <= base_buf_sva_mut_7_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_29_cse = '1' ) THEN
        m_buf_sva_mut_8_8 <= m_buf_sva_mut_8_7;
        base_buf_sva_mut_8_8 <= base_buf_sva_mut_8_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_30_cse = '1' ) THEN
        m_buf_sva_mut_9_8 <= m_buf_sva_mut_9_7;
        base_buf_sva_mut_9_8 <= base_buf_sva_mut_9_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_31_cse = '1' ) THEN
        m_buf_sva_mut_10_8 <= m_buf_sva_mut_10_7;
        base_buf_sva_mut_10_8 <= base_buf_sva_mut_10_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_32_cse = '1' ) THEN
        m_buf_sva_mut_8 <= m_buf_sva_mut_7;
        base_buf_sva_mut_8 <= base_buf_sva_mut_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_8 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_53) = '1' ) THEN
        result_rem_11cyc_st_8 <= result_rem_11cyc_st_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_33_cse = '1' ) THEN
        m_buf_sva_mut_1_7 <= m_buf_sva_mut_1_6;
        base_buf_sva_mut_1_7 <= base_buf_sva_mut_1_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_34_cse = '1' ) THEN
        m_buf_sva_mut_2_7 <= m_buf_sva_mut_2_6;
        base_buf_sva_mut_2_7 <= base_buf_sva_mut_2_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_35_cse = '1' ) THEN
        m_buf_sva_mut_3_7 <= m_buf_sva_mut_3_6;
        base_buf_sva_mut_3_7 <= base_buf_sva_mut_3_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_36_cse = '1' ) THEN
        m_buf_sva_mut_4_7 <= m_buf_sva_mut_4_6;
        base_buf_sva_mut_4_7 <= base_buf_sva_mut_4_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_37_cse = '1' ) THEN
        m_buf_sva_mut_5_7 <= m_buf_sva_mut_5_6;
        base_buf_sva_mut_5_7 <= base_buf_sva_mut_5_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_38_cse = '1' ) THEN
        m_buf_sva_mut_6_7 <= m_buf_sva_mut_6_6;
        base_buf_sva_mut_6_7 <= base_buf_sva_mut_6_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_39_cse = '1' ) THEN
        m_buf_sva_mut_7_7 <= m_buf_sva_mut_7_6;
        base_buf_sva_mut_7_7 <= base_buf_sva_mut_7_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_40_cse = '1' ) THEN
        m_buf_sva_mut_8_7 <= m_buf_sva_mut_8_6;
        base_buf_sva_mut_8_7 <= base_buf_sva_mut_8_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_41_cse = '1' ) THEN
        m_buf_sva_mut_9_7 <= m_buf_sva_mut_9_6;
        base_buf_sva_mut_9_7 <= base_buf_sva_mut_9_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_42_cse = '1' ) THEN
        m_buf_sva_mut_10_7 <= m_buf_sva_mut_10_6;
        base_buf_sva_mut_10_7 <= base_buf_sva_mut_10_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_43_cse = '1' ) THEN
        m_buf_sva_mut_7 <= m_buf_sva_mut_6;
        base_buf_sva_mut_7 <= base_buf_sva_mut_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_7 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_79) = '1' ) THEN
        result_rem_11cyc_st_7 <= result_rem_11cyc_st_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_44_cse = '1' ) THEN
        m_buf_sva_mut_1_6 <= m_buf_sva_mut_1_5;
        base_buf_sva_mut_1_6 <= base_buf_sva_mut_1_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_45_cse = '1' ) THEN
        m_buf_sva_mut_2_6 <= m_buf_sva_mut_2_5;
        base_buf_sva_mut_2_6 <= base_buf_sva_mut_2_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_46_cse = '1' ) THEN
        m_buf_sva_mut_3_6 <= m_buf_sva_mut_3_5;
        base_buf_sva_mut_3_6 <= base_buf_sva_mut_3_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_47_cse = '1' ) THEN
        m_buf_sva_mut_4_6 <= m_buf_sva_mut_4_5;
        base_buf_sva_mut_4_6 <= base_buf_sva_mut_4_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_48_cse = '1' ) THEN
        m_buf_sva_mut_5_6 <= m_buf_sva_mut_5_5;
        base_buf_sva_mut_5_6 <= base_buf_sva_mut_5_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_49_cse = '1' ) THEN
        m_buf_sva_mut_6_6 <= m_buf_sva_mut_6_5;
        base_buf_sva_mut_6_6 <= base_buf_sva_mut_6_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_50_cse = '1' ) THEN
        m_buf_sva_mut_7_6 <= m_buf_sva_mut_7_5;
        base_buf_sva_mut_7_6 <= base_buf_sva_mut_7_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_51_cse = '1' ) THEN
        m_buf_sva_mut_8_6 <= m_buf_sva_mut_8_5;
        base_buf_sva_mut_8_6 <= base_buf_sva_mut_8_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_52_cse = '1' ) THEN
        m_buf_sva_mut_9_6 <= m_buf_sva_mut_9_5;
        base_buf_sva_mut_9_6 <= base_buf_sva_mut_9_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_53_cse = '1' ) THEN
        m_buf_sva_mut_10_6 <= m_buf_sva_mut_10_5;
        base_buf_sva_mut_10_6 <= base_buf_sva_mut_10_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_54_cse = '1' ) THEN
        m_buf_sva_mut_6 <= m_buf_sva_mut_5;
        base_buf_sva_mut_6 <= base_buf_sva_mut_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_6 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_105) = '1' ) THEN
        result_rem_11cyc_st_6 <= result_rem_11cyc_st_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_55_cse = '1' ) THEN
        m_buf_sva_mut_1_5 <= m_buf_sva_mut_1_4;
        base_buf_sva_mut_1_5 <= base_buf_sva_mut_1_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_56_cse = '1' ) THEN
        m_buf_sva_mut_2_5 <= m_buf_sva_mut_2_4;
        base_buf_sva_mut_2_5 <= base_buf_sva_mut_2_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_57_cse = '1' ) THEN
        m_buf_sva_mut_3_5 <= m_buf_sva_mut_3_4;
        base_buf_sva_mut_3_5 <= base_buf_sva_mut_3_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_58_cse = '1' ) THEN
        m_buf_sva_mut_4_5 <= m_buf_sva_mut_4_4;
        base_buf_sva_mut_4_5 <= base_buf_sva_mut_4_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_59_cse = '1' ) THEN
        m_buf_sva_mut_5_5 <= m_buf_sva_mut_5_4;
        base_buf_sva_mut_5_5 <= base_buf_sva_mut_5_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_60_cse = '1' ) THEN
        m_buf_sva_mut_6_5 <= m_buf_sva_mut_6_4;
        base_buf_sva_mut_6_5 <= base_buf_sva_mut_6_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_61_cse = '1' ) THEN
        m_buf_sva_mut_7_5 <= m_buf_sva_mut_7_4;
        base_buf_sva_mut_7_5 <= base_buf_sva_mut_7_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_62_cse = '1' ) THEN
        m_buf_sva_mut_8_5 <= m_buf_sva_mut_8_4;
        base_buf_sva_mut_8_5 <= base_buf_sva_mut_8_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_63_cse = '1' ) THEN
        m_buf_sva_mut_9_5 <= m_buf_sva_mut_9_4;
        base_buf_sva_mut_9_5 <= base_buf_sva_mut_9_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_64_cse = '1' ) THEN
        m_buf_sva_mut_10_5 <= m_buf_sva_mut_10_4;
        base_buf_sva_mut_10_5 <= base_buf_sva_mut_10_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_65_cse = '1' ) THEN
        m_buf_sva_mut_5 <= m_buf_sva_mut_4;
        base_buf_sva_mut_5 <= base_buf_sva_mut_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_5 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_130) = '1' ) THEN
        result_rem_11cyc_st_5 <= result_rem_11cyc_st_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_66_cse = '1' ) THEN
        m_buf_sva_mut_1_4 <= m_buf_sva_mut_1_3;
        base_buf_sva_mut_1_4 <= base_buf_sva_mut_1_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_67_cse = '1' ) THEN
        m_buf_sva_mut_2_4 <= m_buf_sva_mut_2_3;
        base_buf_sva_mut_2_4 <= base_buf_sva_mut_2_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_68_cse = '1' ) THEN
        m_buf_sva_mut_3_4 <= m_buf_sva_mut_3_3;
        base_buf_sva_mut_3_4 <= base_buf_sva_mut_3_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_69_cse = '1' ) THEN
        m_buf_sva_mut_4_4 <= m_buf_sva_mut_4_3;
        base_buf_sva_mut_4_4 <= base_buf_sva_mut_4_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_70_cse = '1' ) THEN
        m_buf_sva_mut_5_4 <= m_buf_sva_mut_5_3;
        base_buf_sva_mut_5_4 <= base_buf_sva_mut_5_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_71_cse = '1' ) THEN
        m_buf_sva_mut_6_4 <= m_buf_sva_mut_6_3;
        base_buf_sva_mut_6_4 <= base_buf_sva_mut_6_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_72_cse = '1' ) THEN
        m_buf_sva_mut_7_4 <= m_buf_sva_mut_7_3;
        base_buf_sva_mut_7_4 <= base_buf_sva_mut_7_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_73_cse = '1' ) THEN
        m_buf_sva_mut_8_4 <= m_buf_sva_mut_8_3;
        base_buf_sva_mut_8_4 <= base_buf_sva_mut_8_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_74_cse = '1' ) THEN
        m_buf_sva_mut_9_4 <= m_buf_sva_mut_9_3;
        base_buf_sva_mut_9_4 <= base_buf_sva_mut_9_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_75_cse = '1' ) THEN
        m_buf_sva_mut_10_4 <= m_buf_sva_mut_10_3;
        base_buf_sva_mut_10_4 <= base_buf_sva_mut_10_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_76_cse = '1' ) THEN
        m_buf_sva_mut_4 <= m_buf_sva_mut_3;
        base_buf_sva_mut_4 <= base_buf_sva_mut_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_4 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_156) = '1' ) THEN
        result_rem_11cyc_st_4 <= result_rem_11cyc_st_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_77_cse = '1' ) THEN
        m_buf_sva_mut_1_3 <= m_buf_sva_mut_1_2;
        base_buf_sva_mut_1_3 <= base_buf_sva_mut_1_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_78_cse = '1' ) THEN
        m_buf_sva_mut_2_3 <= m_buf_sva_mut_2_2;
        base_buf_sva_mut_2_3 <= base_buf_sva_mut_2_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_79_cse = '1' ) THEN
        m_buf_sva_mut_3_3 <= m_buf_sva_mut_3_2;
        base_buf_sva_mut_3_3 <= base_buf_sva_mut_3_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_80_cse = '1' ) THEN
        m_buf_sva_mut_4_3 <= m_buf_sva_mut_4_2;
        base_buf_sva_mut_4_3 <= base_buf_sva_mut_4_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_81_cse = '1' ) THEN
        m_buf_sva_mut_5_3 <= m_buf_sva_mut_5_2;
        base_buf_sva_mut_5_3 <= base_buf_sva_mut_5_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_82_cse = '1' ) THEN
        m_buf_sva_mut_6_3 <= m_buf_sva_mut_6_2;
        base_buf_sva_mut_6_3 <= base_buf_sva_mut_6_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_83_cse = '1' ) THEN
        m_buf_sva_mut_7_3 <= m_buf_sva_mut_7_2;
        base_buf_sva_mut_7_3 <= base_buf_sva_mut_7_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_84_cse = '1' ) THEN
        m_buf_sva_mut_8_3 <= m_buf_sva_mut_8_2;
        base_buf_sva_mut_8_3 <= base_buf_sva_mut_8_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_85_cse = '1' ) THEN
        m_buf_sva_mut_9_3 <= m_buf_sva_mut_9_2;
        base_buf_sva_mut_9_3 <= base_buf_sva_mut_9_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_86_cse = '1' ) THEN
        m_buf_sva_mut_10_3 <= m_buf_sva_mut_10_2;
        base_buf_sva_mut_10_3 <= base_buf_sva_mut_10_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_87_cse = '1' ) THEN
        m_buf_sva_mut_3 <= m_buf_sva_mut_2;
        base_buf_sva_mut_3 <= base_buf_sva_mut_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_3 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_182) = '1' ) THEN
        result_rem_11cyc_st_3 <= result_rem_11cyc_st_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_88_cse = '1' ) THEN
        m_buf_sva_mut_1_2 <= result_rem_12_cmp_1_b;
        base_buf_sva_mut_1_2 <= result_rem_12_cmp_1_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_89_cse = '1' ) THEN
        m_buf_sva_mut_2_2 <= result_rem_12_cmp_2_b;
        base_buf_sva_mut_2_2 <= result_rem_12_cmp_2_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_90_cse = '1' ) THEN
        m_buf_sva_mut_3_2 <= result_rem_12_cmp_3_b;
        base_buf_sva_mut_3_2 <= result_rem_12_cmp_3_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_91_cse = '1' ) THEN
        m_buf_sva_mut_4_2 <= result_rem_12_cmp_4_b;
        base_buf_sva_mut_4_2 <= result_rem_12_cmp_4_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_92_cse = '1' ) THEN
        m_buf_sva_mut_5_2 <= result_rem_12_cmp_5_b;
        base_buf_sva_mut_5_2 <= result_rem_12_cmp_5_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_93_cse = '1' ) THEN
        m_buf_sva_mut_6_2 <= result_rem_12_cmp_6_b;
        base_buf_sva_mut_6_2 <= result_rem_12_cmp_6_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_94_cse = '1' ) THEN
        m_buf_sva_mut_7_2 <= result_rem_12_cmp_7_b;
        base_buf_sva_mut_7_2 <= result_rem_12_cmp_7_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_95_cse = '1' ) THEN
        m_buf_sva_mut_8_2 <= result_rem_12_cmp_8_b;
        base_buf_sva_mut_8_2 <= result_rem_12_cmp_8_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_96_cse = '1' ) THEN
        m_buf_sva_mut_9_2 <= result_rem_12_cmp_9_b;
        base_buf_sva_mut_9_2 <= result_rem_12_cmp_9_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_97_cse = '1' ) THEN
        m_buf_sva_mut_10_2 <= result_rem_12_cmp_10_b;
        base_buf_sva_mut_10_2 <= result_rem_12_cmp_10_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_98_cse = '1' ) THEN
        m_buf_sva_mut_2 <= result_rem_12_cmp_b;
        base_buf_sva_mut_2 <= result_rem_12_cmp_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_2 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_208) = '1' ) THEN
        result_rem_11cyc_st_2 <= result_rem_11cyc;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND ccs_ccore_start_rsci_idat) = '1' ) THEN
        result_rem_11cyc <= result_result_acc_tmp;
      END IF;
    END IF;
  END PROCESS;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    modulo_dev
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_dev IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_dev;

ARCHITECTURE v1 OF modulo_dev IS
  -- Default Constants

  COMPONENT modulo_dev_core
    PORT(
      base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_dev_core_inst_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_core_inst_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_core_inst_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  modulo_dev_core_inst : modulo_dev_core
    PORT MAP(
      base_rsc_dat => modulo_dev_core_inst_base_rsc_dat,
      m_rsc_dat => modulo_dev_core_inst_m_rsc_dat,
      return_rsc_z => modulo_dev_core_inst_return_rsc_z,
      ccs_ccore_start_rsc_dat => ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_srst => ccs_ccore_srst,
      ccs_ccore_en => ccs_ccore_en
    );
  modulo_dev_core_inst_base_rsc_dat <= base_rsc_dat;
  modulo_dev_core_inst_m_rsc_dat <= m_rsc_dat;
  return_rsc_z <= modulo_dev_core_inst_return_rsc_z;

END v1;




--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Thu Aug 26 04:28:40 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen;

ARCHITECTURE v13 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    COMP_LOOP_C_28_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_56_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_84_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_112_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_140_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_168_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_196_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_224_tr0 : IN STD_LOGIC;
    VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_1_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_core_core_fsm;

ARCHITECTURE v13 OF inPlaceNTT_DIF_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIF_core_core_fsm_1
  TYPE inPlaceNTT_DIF_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, COMP_LOOP_C_0,
      COMP_LOOP_C_1, COMP_LOOP_C_2, COMP_LOOP_C_3, COMP_LOOP_C_4, COMP_LOOP_C_5,
      COMP_LOOP_C_6, COMP_LOOP_C_7, COMP_LOOP_C_8, COMP_LOOP_C_9, COMP_LOOP_C_10,
      COMP_LOOP_C_11, COMP_LOOP_C_12, COMP_LOOP_C_13, COMP_LOOP_C_14, COMP_LOOP_C_15,
      COMP_LOOP_C_16, COMP_LOOP_C_17, COMP_LOOP_C_18, COMP_LOOP_C_19, COMP_LOOP_C_20,
      COMP_LOOP_C_21, COMP_LOOP_C_22, COMP_LOOP_C_23, COMP_LOOP_C_24, COMP_LOOP_C_25,
      COMP_LOOP_C_26, COMP_LOOP_C_27, COMP_LOOP_C_28, COMP_LOOP_C_29, COMP_LOOP_C_30,
      COMP_LOOP_C_31, COMP_LOOP_C_32, COMP_LOOP_C_33, COMP_LOOP_C_34, COMP_LOOP_C_35,
      COMP_LOOP_C_36, COMP_LOOP_C_37, COMP_LOOP_C_38, COMP_LOOP_C_39, COMP_LOOP_C_40,
      COMP_LOOP_C_41, COMP_LOOP_C_42, COMP_LOOP_C_43, COMP_LOOP_C_44, COMP_LOOP_C_45,
      COMP_LOOP_C_46, COMP_LOOP_C_47, COMP_LOOP_C_48, COMP_LOOP_C_49, COMP_LOOP_C_50,
      COMP_LOOP_C_51, COMP_LOOP_C_52, COMP_LOOP_C_53, COMP_LOOP_C_54, COMP_LOOP_C_55,
      COMP_LOOP_C_56, COMP_LOOP_C_57, COMP_LOOP_C_58, COMP_LOOP_C_59, COMP_LOOP_C_60,
      COMP_LOOP_C_61, COMP_LOOP_C_62, COMP_LOOP_C_63, COMP_LOOP_C_64, COMP_LOOP_C_65,
      COMP_LOOP_C_66, COMP_LOOP_C_67, COMP_LOOP_C_68, COMP_LOOP_C_69, COMP_LOOP_C_70,
      COMP_LOOP_C_71, COMP_LOOP_C_72, COMP_LOOP_C_73, COMP_LOOP_C_74, COMP_LOOP_C_75,
      COMP_LOOP_C_76, COMP_LOOP_C_77, COMP_LOOP_C_78, COMP_LOOP_C_79, COMP_LOOP_C_80,
      COMP_LOOP_C_81, COMP_LOOP_C_82, COMP_LOOP_C_83, COMP_LOOP_C_84, COMP_LOOP_C_85,
      COMP_LOOP_C_86, COMP_LOOP_C_87, COMP_LOOP_C_88, COMP_LOOP_C_89, COMP_LOOP_C_90,
      COMP_LOOP_C_91, COMP_LOOP_C_92, COMP_LOOP_C_93, COMP_LOOP_C_94, COMP_LOOP_C_95,
      COMP_LOOP_C_96, COMP_LOOP_C_97, COMP_LOOP_C_98, COMP_LOOP_C_99, COMP_LOOP_C_100,
      COMP_LOOP_C_101, COMP_LOOP_C_102, COMP_LOOP_C_103, COMP_LOOP_C_104, COMP_LOOP_C_105,
      COMP_LOOP_C_106, COMP_LOOP_C_107, COMP_LOOP_C_108, COMP_LOOP_C_109, COMP_LOOP_C_110,
      COMP_LOOP_C_111, COMP_LOOP_C_112, COMP_LOOP_C_113, COMP_LOOP_C_114, COMP_LOOP_C_115,
      COMP_LOOP_C_116, COMP_LOOP_C_117, COMP_LOOP_C_118, COMP_LOOP_C_119, COMP_LOOP_C_120,
      COMP_LOOP_C_121, COMP_LOOP_C_122, COMP_LOOP_C_123, COMP_LOOP_C_124, COMP_LOOP_C_125,
      COMP_LOOP_C_126, COMP_LOOP_C_127, COMP_LOOP_C_128, COMP_LOOP_C_129, COMP_LOOP_C_130,
      COMP_LOOP_C_131, COMP_LOOP_C_132, COMP_LOOP_C_133, COMP_LOOP_C_134, COMP_LOOP_C_135,
      COMP_LOOP_C_136, COMP_LOOP_C_137, COMP_LOOP_C_138, COMP_LOOP_C_139, COMP_LOOP_C_140,
      COMP_LOOP_C_141, COMP_LOOP_C_142, COMP_LOOP_C_143, COMP_LOOP_C_144, COMP_LOOP_C_145,
      COMP_LOOP_C_146, COMP_LOOP_C_147, COMP_LOOP_C_148, COMP_LOOP_C_149, COMP_LOOP_C_150,
      COMP_LOOP_C_151, COMP_LOOP_C_152, COMP_LOOP_C_153, COMP_LOOP_C_154, COMP_LOOP_C_155,
      COMP_LOOP_C_156, COMP_LOOP_C_157, COMP_LOOP_C_158, COMP_LOOP_C_159, COMP_LOOP_C_160,
      COMP_LOOP_C_161, COMP_LOOP_C_162, COMP_LOOP_C_163, COMP_LOOP_C_164, COMP_LOOP_C_165,
      COMP_LOOP_C_166, COMP_LOOP_C_167, COMP_LOOP_C_168, COMP_LOOP_C_169, COMP_LOOP_C_170,
      COMP_LOOP_C_171, COMP_LOOP_C_172, COMP_LOOP_C_173, COMP_LOOP_C_174, COMP_LOOP_C_175,
      COMP_LOOP_C_176, COMP_LOOP_C_177, COMP_LOOP_C_178, COMP_LOOP_C_179, COMP_LOOP_C_180,
      COMP_LOOP_C_181, COMP_LOOP_C_182, COMP_LOOP_C_183, COMP_LOOP_C_184, COMP_LOOP_C_185,
      COMP_LOOP_C_186, COMP_LOOP_C_187, COMP_LOOP_C_188, COMP_LOOP_C_189, COMP_LOOP_C_190,
      COMP_LOOP_C_191, COMP_LOOP_C_192, COMP_LOOP_C_193, COMP_LOOP_C_194, COMP_LOOP_C_195,
      COMP_LOOP_C_196, COMP_LOOP_C_197, COMP_LOOP_C_198, COMP_LOOP_C_199, COMP_LOOP_C_200,
      COMP_LOOP_C_201, COMP_LOOP_C_202, COMP_LOOP_C_203, COMP_LOOP_C_204, COMP_LOOP_C_205,
      COMP_LOOP_C_206, COMP_LOOP_C_207, COMP_LOOP_C_208, COMP_LOOP_C_209, COMP_LOOP_C_210,
      COMP_LOOP_C_211, COMP_LOOP_C_212, COMP_LOOP_C_213, COMP_LOOP_C_214, COMP_LOOP_C_215,
      COMP_LOOP_C_216, COMP_LOOP_C_217, COMP_LOOP_C_218, COMP_LOOP_C_219, COMP_LOOP_C_220,
      COMP_LOOP_C_221, COMP_LOOP_C_222, COMP_LOOP_C_223, COMP_LOOP_C_224, VEC_LOOP_C_0,
      STAGE_LOOP_C_1, main_C_1);

  SIGNAL state_var : inPlaceNTT_DIF_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIF_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIF_core_core_fsm_1 : PROCESS (COMP_LOOP_C_28_tr0, COMP_LOOP_C_56_tr0,
      COMP_LOOP_C_84_tr0, COMP_LOOP_C_112_tr0, COMP_LOOP_C_140_tr0, COMP_LOOP_C_168_tr0,
      COMP_LOOP_C_196_tr0, COMP_LOOP_C_224_tr0, VEC_LOOP_C_0_tr0, STAGE_LOOP_C_1_tr0,
      state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001");
        state_var_NS <= COMP_LOOP_C_0;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011");
        state_var_NS <= COMP_LOOP_C_2;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101");
        state_var_NS <= COMP_LOOP_C_4;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110");
        state_var_NS <= COMP_LOOP_C_5;
      WHEN COMP_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111");
        state_var_NS <= COMP_LOOP_C_6;
      WHEN COMP_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000");
        state_var_NS <= COMP_LOOP_C_7;
      WHEN COMP_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001");
        state_var_NS <= COMP_LOOP_C_8;
      WHEN COMP_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010");
        state_var_NS <= COMP_LOOP_C_9;
      WHEN COMP_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011");
        state_var_NS <= COMP_LOOP_C_10;
      WHEN COMP_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100");
        state_var_NS <= COMP_LOOP_C_11;
      WHEN COMP_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101");
        state_var_NS <= COMP_LOOP_C_12;
      WHEN COMP_LOOP_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110");
        state_var_NS <= COMP_LOOP_C_13;
      WHEN COMP_LOOP_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111");
        state_var_NS <= COMP_LOOP_C_14;
      WHEN COMP_LOOP_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000");
        state_var_NS <= COMP_LOOP_C_15;
      WHEN COMP_LOOP_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001");
        state_var_NS <= COMP_LOOP_C_16;
      WHEN COMP_LOOP_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010");
        state_var_NS <= COMP_LOOP_C_17;
      WHEN COMP_LOOP_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011");
        state_var_NS <= COMP_LOOP_C_18;
      WHEN COMP_LOOP_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100");
        state_var_NS <= COMP_LOOP_C_19;
      WHEN COMP_LOOP_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101");
        state_var_NS <= COMP_LOOP_C_20;
      WHEN COMP_LOOP_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110");
        state_var_NS <= COMP_LOOP_C_21;
      WHEN COMP_LOOP_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111");
        state_var_NS <= COMP_LOOP_C_22;
      WHEN COMP_LOOP_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000");
        state_var_NS <= COMP_LOOP_C_23;
      WHEN COMP_LOOP_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001");
        state_var_NS <= COMP_LOOP_C_24;
      WHEN COMP_LOOP_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010");
        state_var_NS <= COMP_LOOP_C_25;
      WHEN COMP_LOOP_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011");
        state_var_NS <= COMP_LOOP_C_26;
      WHEN COMP_LOOP_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100");
        state_var_NS <= COMP_LOOP_C_27;
      WHEN COMP_LOOP_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101");
        state_var_NS <= COMP_LOOP_C_28;
      WHEN COMP_LOOP_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110");
        IF ( COMP_LOOP_C_28_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_29;
        END IF;
      WHEN COMP_LOOP_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111");
        state_var_NS <= COMP_LOOP_C_30;
      WHEN COMP_LOOP_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000");
        state_var_NS <= COMP_LOOP_C_31;
      WHEN COMP_LOOP_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001");
        state_var_NS <= COMP_LOOP_C_32;
      WHEN COMP_LOOP_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010");
        state_var_NS <= COMP_LOOP_C_33;
      WHEN COMP_LOOP_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011");
        state_var_NS <= COMP_LOOP_C_34;
      WHEN COMP_LOOP_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100");
        state_var_NS <= COMP_LOOP_C_35;
      WHEN COMP_LOOP_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101");
        state_var_NS <= COMP_LOOP_C_36;
      WHEN COMP_LOOP_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110");
        state_var_NS <= COMP_LOOP_C_37;
      WHEN COMP_LOOP_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111");
        state_var_NS <= COMP_LOOP_C_38;
      WHEN COMP_LOOP_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000");
        state_var_NS <= COMP_LOOP_C_39;
      WHEN COMP_LOOP_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001");
        state_var_NS <= COMP_LOOP_C_40;
      WHEN COMP_LOOP_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010");
        state_var_NS <= COMP_LOOP_C_41;
      WHEN COMP_LOOP_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011");
        state_var_NS <= COMP_LOOP_C_42;
      WHEN COMP_LOOP_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100");
        state_var_NS <= COMP_LOOP_C_43;
      WHEN COMP_LOOP_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101");
        state_var_NS <= COMP_LOOP_C_44;
      WHEN COMP_LOOP_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110");
        state_var_NS <= COMP_LOOP_C_45;
      WHEN COMP_LOOP_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111");
        state_var_NS <= COMP_LOOP_C_46;
      WHEN COMP_LOOP_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000");
        state_var_NS <= COMP_LOOP_C_47;
      WHEN COMP_LOOP_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001");
        state_var_NS <= COMP_LOOP_C_48;
      WHEN COMP_LOOP_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010");
        state_var_NS <= COMP_LOOP_C_49;
      WHEN COMP_LOOP_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011");
        state_var_NS <= COMP_LOOP_C_50;
      WHEN COMP_LOOP_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100");
        state_var_NS <= COMP_LOOP_C_51;
      WHEN COMP_LOOP_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101");
        state_var_NS <= COMP_LOOP_C_52;
      WHEN COMP_LOOP_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110");
        state_var_NS <= COMP_LOOP_C_53;
      WHEN COMP_LOOP_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111");
        state_var_NS <= COMP_LOOP_C_54;
      WHEN COMP_LOOP_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000");
        state_var_NS <= COMP_LOOP_C_55;
      WHEN COMP_LOOP_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001");
        state_var_NS <= COMP_LOOP_C_56;
      WHEN COMP_LOOP_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010");
        IF ( COMP_LOOP_C_56_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_57;
        END IF;
      WHEN COMP_LOOP_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011");
        state_var_NS <= COMP_LOOP_C_58;
      WHEN COMP_LOOP_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100");
        state_var_NS <= COMP_LOOP_C_59;
      WHEN COMP_LOOP_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101");
        state_var_NS <= COMP_LOOP_C_60;
      WHEN COMP_LOOP_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110");
        state_var_NS <= COMP_LOOP_C_61;
      WHEN COMP_LOOP_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111");
        state_var_NS <= COMP_LOOP_C_62;
      WHEN COMP_LOOP_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000");
        state_var_NS <= COMP_LOOP_C_63;
      WHEN COMP_LOOP_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001");
        state_var_NS <= COMP_LOOP_C_64;
      WHEN COMP_LOOP_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010");
        state_var_NS <= COMP_LOOP_C_65;
      WHEN COMP_LOOP_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011");
        state_var_NS <= COMP_LOOP_C_66;
      WHEN COMP_LOOP_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100");
        state_var_NS <= COMP_LOOP_C_67;
      WHEN COMP_LOOP_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101");
        state_var_NS <= COMP_LOOP_C_68;
      WHEN COMP_LOOP_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110");
        state_var_NS <= COMP_LOOP_C_69;
      WHEN COMP_LOOP_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111");
        state_var_NS <= COMP_LOOP_C_70;
      WHEN COMP_LOOP_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000");
        state_var_NS <= COMP_LOOP_C_71;
      WHEN COMP_LOOP_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001");
        state_var_NS <= COMP_LOOP_C_72;
      WHEN COMP_LOOP_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010");
        state_var_NS <= COMP_LOOP_C_73;
      WHEN COMP_LOOP_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011");
        state_var_NS <= COMP_LOOP_C_74;
      WHEN COMP_LOOP_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100");
        state_var_NS <= COMP_LOOP_C_75;
      WHEN COMP_LOOP_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101");
        state_var_NS <= COMP_LOOP_C_76;
      WHEN COMP_LOOP_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110");
        state_var_NS <= COMP_LOOP_C_77;
      WHEN COMP_LOOP_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111");
        state_var_NS <= COMP_LOOP_C_78;
      WHEN COMP_LOOP_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000");
        state_var_NS <= COMP_LOOP_C_79;
      WHEN COMP_LOOP_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001");
        state_var_NS <= COMP_LOOP_C_80;
      WHEN COMP_LOOP_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010");
        state_var_NS <= COMP_LOOP_C_81;
      WHEN COMP_LOOP_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011");
        state_var_NS <= COMP_LOOP_C_82;
      WHEN COMP_LOOP_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100");
        state_var_NS <= COMP_LOOP_C_83;
      WHEN COMP_LOOP_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101");
        state_var_NS <= COMP_LOOP_C_84;
      WHEN COMP_LOOP_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110");
        IF ( COMP_LOOP_C_84_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_85;
        END IF;
      WHEN COMP_LOOP_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111");
        state_var_NS <= COMP_LOOP_C_86;
      WHEN COMP_LOOP_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000");
        state_var_NS <= COMP_LOOP_C_87;
      WHEN COMP_LOOP_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001");
        state_var_NS <= COMP_LOOP_C_88;
      WHEN COMP_LOOP_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010");
        state_var_NS <= COMP_LOOP_C_89;
      WHEN COMP_LOOP_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011");
        state_var_NS <= COMP_LOOP_C_90;
      WHEN COMP_LOOP_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100");
        state_var_NS <= COMP_LOOP_C_91;
      WHEN COMP_LOOP_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101");
        state_var_NS <= COMP_LOOP_C_92;
      WHEN COMP_LOOP_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110");
        state_var_NS <= COMP_LOOP_C_93;
      WHEN COMP_LOOP_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111");
        state_var_NS <= COMP_LOOP_C_94;
      WHEN COMP_LOOP_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000");
        state_var_NS <= COMP_LOOP_C_95;
      WHEN COMP_LOOP_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001");
        state_var_NS <= COMP_LOOP_C_96;
      WHEN COMP_LOOP_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010");
        state_var_NS <= COMP_LOOP_C_97;
      WHEN COMP_LOOP_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011");
        state_var_NS <= COMP_LOOP_C_98;
      WHEN COMP_LOOP_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100");
        state_var_NS <= COMP_LOOP_C_99;
      WHEN COMP_LOOP_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101");
        state_var_NS <= COMP_LOOP_C_100;
      WHEN COMP_LOOP_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110");
        state_var_NS <= COMP_LOOP_C_101;
      WHEN COMP_LOOP_C_101 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111");
        state_var_NS <= COMP_LOOP_C_102;
      WHEN COMP_LOOP_C_102 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000");
        state_var_NS <= COMP_LOOP_C_103;
      WHEN COMP_LOOP_C_103 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001");
        state_var_NS <= COMP_LOOP_C_104;
      WHEN COMP_LOOP_C_104 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010");
        state_var_NS <= COMP_LOOP_C_105;
      WHEN COMP_LOOP_C_105 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011");
        state_var_NS <= COMP_LOOP_C_106;
      WHEN COMP_LOOP_C_106 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100");
        state_var_NS <= COMP_LOOP_C_107;
      WHEN COMP_LOOP_C_107 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101");
        state_var_NS <= COMP_LOOP_C_108;
      WHEN COMP_LOOP_C_108 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110");
        state_var_NS <= COMP_LOOP_C_109;
      WHEN COMP_LOOP_C_109 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111");
        state_var_NS <= COMP_LOOP_C_110;
      WHEN COMP_LOOP_C_110 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000");
        state_var_NS <= COMP_LOOP_C_111;
      WHEN COMP_LOOP_C_111 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001");
        state_var_NS <= COMP_LOOP_C_112;
      WHEN COMP_LOOP_C_112 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010");
        IF ( COMP_LOOP_C_112_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_113;
        END IF;
      WHEN COMP_LOOP_C_113 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011");
        state_var_NS <= COMP_LOOP_C_114;
      WHEN COMP_LOOP_C_114 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100");
        state_var_NS <= COMP_LOOP_C_115;
      WHEN COMP_LOOP_C_115 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101");
        state_var_NS <= COMP_LOOP_C_116;
      WHEN COMP_LOOP_C_116 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110");
        state_var_NS <= COMP_LOOP_C_117;
      WHEN COMP_LOOP_C_117 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111");
        state_var_NS <= COMP_LOOP_C_118;
      WHEN COMP_LOOP_C_118 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000");
        state_var_NS <= COMP_LOOP_C_119;
      WHEN COMP_LOOP_C_119 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001");
        state_var_NS <= COMP_LOOP_C_120;
      WHEN COMP_LOOP_C_120 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010");
        state_var_NS <= COMP_LOOP_C_121;
      WHEN COMP_LOOP_C_121 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011");
        state_var_NS <= COMP_LOOP_C_122;
      WHEN COMP_LOOP_C_122 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100");
        state_var_NS <= COMP_LOOP_C_123;
      WHEN COMP_LOOP_C_123 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101");
        state_var_NS <= COMP_LOOP_C_124;
      WHEN COMP_LOOP_C_124 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110");
        state_var_NS <= COMP_LOOP_C_125;
      WHEN COMP_LOOP_C_125 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111");
        state_var_NS <= COMP_LOOP_C_126;
      WHEN COMP_LOOP_C_126 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000");
        state_var_NS <= COMP_LOOP_C_127;
      WHEN COMP_LOOP_C_127 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001");
        state_var_NS <= COMP_LOOP_C_128;
      WHEN COMP_LOOP_C_128 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010");
        state_var_NS <= COMP_LOOP_C_129;
      WHEN COMP_LOOP_C_129 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011");
        state_var_NS <= COMP_LOOP_C_130;
      WHEN COMP_LOOP_C_130 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100");
        state_var_NS <= COMP_LOOP_C_131;
      WHEN COMP_LOOP_C_131 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101");
        state_var_NS <= COMP_LOOP_C_132;
      WHEN COMP_LOOP_C_132 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110");
        state_var_NS <= COMP_LOOP_C_133;
      WHEN COMP_LOOP_C_133 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111");
        state_var_NS <= COMP_LOOP_C_134;
      WHEN COMP_LOOP_C_134 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000");
        state_var_NS <= COMP_LOOP_C_135;
      WHEN COMP_LOOP_C_135 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001");
        state_var_NS <= COMP_LOOP_C_136;
      WHEN COMP_LOOP_C_136 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010");
        state_var_NS <= COMP_LOOP_C_137;
      WHEN COMP_LOOP_C_137 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011");
        state_var_NS <= COMP_LOOP_C_138;
      WHEN COMP_LOOP_C_138 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100");
        state_var_NS <= COMP_LOOP_C_139;
      WHEN COMP_LOOP_C_139 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101");
        state_var_NS <= COMP_LOOP_C_140;
      WHEN COMP_LOOP_C_140 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110");
        IF ( COMP_LOOP_C_140_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_141;
        END IF;
      WHEN COMP_LOOP_C_141 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111");
        state_var_NS <= COMP_LOOP_C_142;
      WHEN COMP_LOOP_C_142 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000");
        state_var_NS <= COMP_LOOP_C_143;
      WHEN COMP_LOOP_C_143 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001");
        state_var_NS <= COMP_LOOP_C_144;
      WHEN COMP_LOOP_C_144 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010");
        state_var_NS <= COMP_LOOP_C_145;
      WHEN COMP_LOOP_C_145 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011");
        state_var_NS <= COMP_LOOP_C_146;
      WHEN COMP_LOOP_C_146 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100");
        state_var_NS <= COMP_LOOP_C_147;
      WHEN COMP_LOOP_C_147 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101");
        state_var_NS <= COMP_LOOP_C_148;
      WHEN COMP_LOOP_C_148 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110");
        state_var_NS <= COMP_LOOP_C_149;
      WHEN COMP_LOOP_C_149 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111");
        state_var_NS <= COMP_LOOP_C_150;
      WHEN COMP_LOOP_C_150 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000");
        state_var_NS <= COMP_LOOP_C_151;
      WHEN COMP_LOOP_C_151 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001");
        state_var_NS <= COMP_LOOP_C_152;
      WHEN COMP_LOOP_C_152 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010");
        state_var_NS <= COMP_LOOP_C_153;
      WHEN COMP_LOOP_C_153 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011");
        state_var_NS <= COMP_LOOP_C_154;
      WHEN COMP_LOOP_C_154 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100");
        state_var_NS <= COMP_LOOP_C_155;
      WHEN COMP_LOOP_C_155 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101");
        state_var_NS <= COMP_LOOP_C_156;
      WHEN COMP_LOOP_C_156 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110");
        state_var_NS <= COMP_LOOP_C_157;
      WHEN COMP_LOOP_C_157 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111");
        state_var_NS <= COMP_LOOP_C_158;
      WHEN COMP_LOOP_C_158 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000");
        state_var_NS <= COMP_LOOP_C_159;
      WHEN COMP_LOOP_C_159 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001");
        state_var_NS <= COMP_LOOP_C_160;
      WHEN COMP_LOOP_C_160 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010");
        state_var_NS <= COMP_LOOP_C_161;
      WHEN COMP_LOOP_C_161 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011");
        state_var_NS <= COMP_LOOP_C_162;
      WHEN COMP_LOOP_C_162 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100");
        state_var_NS <= COMP_LOOP_C_163;
      WHEN COMP_LOOP_C_163 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101");
        state_var_NS <= COMP_LOOP_C_164;
      WHEN COMP_LOOP_C_164 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110");
        state_var_NS <= COMP_LOOP_C_165;
      WHEN COMP_LOOP_C_165 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111");
        state_var_NS <= COMP_LOOP_C_166;
      WHEN COMP_LOOP_C_166 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000");
        state_var_NS <= COMP_LOOP_C_167;
      WHEN COMP_LOOP_C_167 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001");
        state_var_NS <= COMP_LOOP_C_168;
      WHEN COMP_LOOP_C_168 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010");
        IF ( COMP_LOOP_C_168_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_169;
        END IF;
      WHEN COMP_LOOP_C_169 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011");
        state_var_NS <= COMP_LOOP_C_170;
      WHEN COMP_LOOP_C_170 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100");
        state_var_NS <= COMP_LOOP_C_171;
      WHEN COMP_LOOP_C_171 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101");
        state_var_NS <= COMP_LOOP_C_172;
      WHEN COMP_LOOP_C_172 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110");
        state_var_NS <= COMP_LOOP_C_173;
      WHEN COMP_LOOP_C_173 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111");
        state_var_NS <= COMP_LOOP_C_174;
      WHEN COMP_LOOP_C_174 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000");
        state_var_NS <= COMP_LOOP_C_175;
      WHEN COMP_LOOP_C_175 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001");
        state_var_NS <= COMP_LOOP_C_176;
      WHEN COMP_LOOP_C_176 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010");
        state_var_NS <= COMP_LOOP_C_177;
      WHEN COMP_LOOP_C_177 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011");
        state_var_NS <= COMP_LOOP_C_178;
      WHEN COMP_LOOP_C_178 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100");
        state_var_NS <= COMP_LOOP_C_179;
      WHEN COMP_LOOP_C_179 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101");
        state_var_NS <= COMP_LOOP_C_180;
      WHEN COMP_LOOP_C_180 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110");
        state_var_NS <= COMP_LOOP_C_181;
      WHEN COMP_LOOP_C_181 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111");
        state_var_NS <= COMP_LOOP_C_182;
      WHEN COMP_LOOP_C_182 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000");
        state_var_NS <= COMP_LOOP_C_183;
      WHEN COMP_LOOP_C_183 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001");
        state_var_NS <= COMP_LOOP_C_184;
      WHEN COMP_LOOP_C_184 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010");
        state_var_NS <= COMP_LOOP_C_185;
      WHEN COMP_LOOP_C_185 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011");
        state_var_NS <= COMP_LOOP_C_186;
      WHEN COMP_LOOP_C_186 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100");
        state_var_NS <= COMP_LOOP_C_187;
      WHEN COMP_LOOP_C_187 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101");
        state_var_NS <= COMP_LOOP_C_188;
      WHEN COMP_LOOP_C_188 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110");
        state_var_NS <= COMP_LOOP_C_189;
      WHEN COMP_LOOP_C_189 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111");
        state_var_NS <= COMP_LOOP_C_190;
      WHEN COMP_LOOP_C_190 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000");
        state_var_NS <= COMP_LOOP_C_191;
      WHEN COMP_LOOP_C_191 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001");
        state_var_NS <= COMP_LOOP_C_192;
      WHEN COMP_LOOP_C_192 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010");
        state_var_NS <= COMP_LOOP_C_193;
      WHEN COMP_LOOP_C_193 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011");
        state_var_NS <= COMP_LOOP_C_194;
      WHEN COMP_LOOP_C_194 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100");
        state_var_NS <= COMP_LOOP_C_195;
      WHEN COMP_LOOP_C_195 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101");
        state_var_NS <= COMP_LOOP_C_196;
      WHEN COMP_LOOP_C_196 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110");
        IF ( COMP_LOOP_C_196_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_197;
        END IF;
      WHEN COMP_LOOP_C_197 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111");
        state_var_NS <= COMP_LOOP_C_198;
      WHEN COMP_LOOP_C_198 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000");
        state_var_NS <= COMP_LOOP_C_199;
      WHEN COMP_LOOP_C_199 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001");
        state_var_NS <= COMP_LOOP_C_200;
      WHEN COMP_LOOP_C_200 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010");
        state_var_NS <= COMP_LOOP_C_201;
      WHEN COMP_LOOP_C_201 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011");
        state_var_NS <= COMP_LOOP_C_202;
      WHEN COMP_LOOP_C_202 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100");
        state_var_NS <= COMP_LOOP_C_203;
      WHEN COMP_LOOP_C_203 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101");
        state_var_NS <= COMP_LOOP_C_204;
      WHEN COMP_LOOP_C_204 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110");
        state_var_NS <= COMP_LOOP_C_205;
      WHEN COMP_LOOP_C_205 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111");
        state_var_NS <= COMP_LOOP_C_206;
      WHEN COMP_LOOP_C_206 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000");
        state_var_NS <= COMP_LOOP_C_207;
      WHEN COMP_LOOP_C_207 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001");
        state_var_NS <= COMP_LOOP_C_208;
      WHEN COMP_LOOP_C_208 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010");
        state_var_NS <= COMP_LOOP_C_209;
      WHEN COMP_LOOP_C_209 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011");
        state_var_NS <= COMP_LOOP_C_210;
      WHEN COMP_LOOP_C_210 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010100");
        state_var_NS <= COMP_LOOP_C_211;
      WHEN COMP_LOOP_C_211 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010101");
        state_var_NS <= COMP_LOOP_C_212;
      WHEN COMP_LOOP_C_212 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010110");
        state_var_NS <= COMP_LOOP_C_213;
      WHEN COMP_LOOP_C_213 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010111");
        state_var_NS <= COMP_LOOP_C_214;
      WHEN COMP_LOOP_C_214 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011000");
        state_var_NS <= COMP_LOOP_C_215;
      WHEN COMP_LOOP_C_215 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011001");
        state_var_NS <= COMP_LOOP_C_216;
      WHEN COMP_LOOP_C_216 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011010");
        state_var_NS <= COMP_LOOP_C_217;
      WHEN COMP_LOOP_C_217 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011011");
        state_var_NS <= COMP_LOOP_C_218;
      WHEN COMP_LOOP_C_218 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011100");
        state_var_NS <= COMP_LOOP_C_219;
      WHEN COMP_LOOP_C_219 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011101");
        state_var_NS <= COMP_LOOP_C_220;
      WHEN COMP_LOOP_C_220 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011110");
        state_var_NS <= COMP_LOOP_C_221;
      WHEN COMP_LOOP_C_221 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011111");
        state_var_NS <= COMP_LOOP_C_222;
      WHEN COMP_LOOP_C_222 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100000");
        state_var_NS <= COMP_LOOP_C_223;
      WHEN COMP_LOOP_C_223 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100001");
        state_var_NS <= COMP_LOOP_C_224;
      WHEN COMP_LOOP_C_224 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100010");
        IF ( COMP_LOOP_C_224_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100011");
        IF ( VEC_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100100");
        IF ( STAGE_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100101");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS inPlaceNTT_DIF_core_core_fsm_1;

  inPlaceNTT_DIF_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIF_core_core_fsm_1_REG;

END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core_wait_dp IS
  PORT(
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_core_wait_dp;

ARCHITECTURE v13 OF inPlaceNTT_DIF_core_wait_dp IS
  -- Default Constants

BEGIN
  COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en <= ensig_cgo OR ensig_cgo_iro;
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    vec_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_1_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_2_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_3_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_4_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_5_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_6_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_7_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_8_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_9_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_10_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_11_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_12_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_13_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_14_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_15_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_16_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_17_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_18_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_19_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_20_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_21_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_22_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_23_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_24_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_25_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_26_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_27_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_28_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_29_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_30_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_31_i_we_d_pff : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_1_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_2_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_4_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0)
  );
END inPlaceNTT_DIF_core;

ARCHITECTURE v13 OF inPlaceNTT_DIF_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : STD_LOGIC;
  SIGNAL fsm_output : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL nor_tmp_53 : STD_LOGIC;
  SIGNAL or_tmp_142 : STD_LOGIC;
  SIGNAL and_dcpl_28 : STD_LOGIC;
  SIGNAL and_dcpl_29 : STD_LOGIC;
  SIGNAL and_dcpl_30 : STD_LOGIC;
  SIGNAL and_dcpl_31 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_35 : STD_LOGIC;
  SIGNAL and_dcpl_36 : STD_LOGIC;
  SIGNAL and_dcpl_38 : STD_LOGIC;
  SIGNAL nor_tmp_95 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_44 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_46 : STD_LOGIC;
  SIGNAL and_dcpl_48 : STD_LOGIC;
  SIGNAL and_dcpl_49 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL and_dcpl_52 : STD_LOGIC;
  SIGNAL and_dcpl_54 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_56 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_59 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_61 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL and_dcpl_64 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_dcpl_68 : STD_LOGIC;
  SIGNAL and_dcpl_69 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL and_dcpl_71 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_74 : STD_LOGIC;
  SIGNAL and_dcpl_75 : STD_LOGIC;
  SIGNAL and_dcpl_76 : STD_LOGIC;
  SIGNAL and_dcpl_78 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_95 : STD_LOGIC;
  SIGNAL and_dcpl_97 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL mux_tmp_311 : STD_LOGIC;
  SIGNAL mux_tmp_373 : STD_LOGIC;
  SIGNAL mux_tmp_435 : STD_LOGIC;
  SIGNAL mux_tmp_497 : STD_LOGIC;
  SIGNAL mux_tmp_559 : STD_LOGIC;
  SIGNAL mux_tmp_621 : STD_LOGIC;
  SIGNAL mux_tmp_683 : STD_LOGIC;
  SIGNAL mux_tmp_745 : STD_LOGIC;
  SIGNAL mux_tmp_807 : STD_LOGIC;
  SIGNAL mux_tmp_869 : STD_LOGIC;
  SIGNAL mux_tmp_931 : STD_LOGIC;
  SIGNAL mux_tmp_993 : STD_LOGIC;
  SIGNAL mux_tmp_1055 : STD_LOGIC;
  SIGNAL mux_tmp_1117 : STD_LOGIC;
  SIGNAL mux_tmp_1179 : STD_LOGIC;
  SIGNAL mux_tmp_1241 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_172 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_174 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_176 : STD_LOGIC;
  SIGNAL and_dcpl_177 : STD_LOGIC;
  SIGNAL and_dcpl_178 : STD_LOGIC;
  SIGNAL and_dcpl_179 : STD_LOGIC;
  SIGNAL not_tmp_617 : STD_LOGIC;
  SIGNAL not_tmp_618 : STD_LOGIC;
  SIGNAL not_tmp_625 : STD_LOGIC;
  SIGNAL not_tmp_632 : STD_LOGIC;
  SIGNAL mux_tmp_1423 : STD_LOGIC;
  SIGNAL or_tmp_2024 : STD_LOGIC;
  SIGNAL mux_tmp_1424 : STD_LOGIC;
  SIGNAL or_tmp_2025 : STD_LOGIC;
  SIGNAL mux_tmp_1430 : STD_LOGIC;
  SIGNAL and_dcpl_220 : STD_LOGIC;
  SIGNAL and_dcpl_222 : STD_LOGIC;
  SIGNAL and_dcpl_223 : STD_LOGIC;
  SIGNAL and_dcpl_226 : STD_LOGIC;
  SIGNAL and_dcpl_229 : STD_LOGIC;
  SIGNAL and_dcpl_232 : STD_LOGIC;
  SIGNAL and_dcpl_234 : STD_LOGIC;
  SIGNAL and_dcpl_236 : STD_LOGIC;
  SIGNAL and_dcpl_238 : STD_LOGIC;
  SIGNAL nand_tmp_184 : STD_LOGIC;
  SIGNAL mux_tmp_1437 : STD_LOGIC;
  SIGNAL and_dcpl_244 : STD_LOGIC;
  SIGNAL or_dcpl_84 : STD_LOGIC;
  SIGNAL or_tmp_2048 : STD_LOGIC;
  SIGNAL mux_tmp_1452 : STD_LOGIC;
  SIGNAL mux_tmp_1456 : STD_LOGIC;
  SIGNAL mux_tmp_1459 : STD_LOGIC;
  SIGNAL and_tmp_11 : STD_LOGIC;
  SIGNAL or_tmp_2054 : STD_LOGIC;
  SIGNAL not_tmp_692 : STD_LOGIC;
  SIGNAL or_tmp_2057 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL mux_tmp_1468 : STD_LOGIC;
  SIGNAL and_tmp_13 : STD_LOGIC;
  SIGNAL and_dcpl_256 : STD_LOGIC;
  SIGNAL nor_tmp_324 : STD_LOGIC;
  SIGNAL and_dcpl_259 : STD_LOGIC;
  SIGNAL mux_tmp_1482 : STD_LOGIC;
  SIGNAL mux_tmp_1487 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL not_tmp_717 : STD_LOGIC;
  SIGNAL and_dcpl_262 : STD_LOGIC;
  SIGNAL and_dcpl_264 : STD_LOGIC;
  SIGNAL and_dcpl_278 : STD_LOGIC;
  SIGNAL or_tmp_2075 : STD_LOGIC;
  SIGNAL or_dcpl_109 : STD_LOGIC;
  SIGNAL COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_1_cse_6_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL VEC_LOOP_j_10_0_sva_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_k_10_3_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_2_tmp_lshift_ncse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_42_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_2_tmp_mul_idiv_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_3_tmp_lshift_ncse_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_25_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_49_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_psp_sva : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_13_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_1_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_5_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_14_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_3_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_7_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_5_tmp_mul_idiv_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_mul_idiv_sva_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_psp_sva_mx0w0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_119_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_121_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_125_rgt : STD_LOGIC;
  SIGNAL mux_1592_tmp : STD_LOGIC;
  SIGNAL and_298_m1c : STD_LOGIC;
  SIGNAL nor_1117_tmp : STD_LOGIC;
  SIGNAL nor_tmp : STD_LOGIC;
  SIGNAL nor_1119_tmp : STD_LOGIC;
  SIGNAL and_294_tmp : STD_LOGIC;
  SIGNAL reg_COMP_LOOP_k_10_3_ftd : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL or_285_cse : STD_LOGIC;
  SIGNAL nand_443_cse : STD_LOGIC;
  SIGNAL nand_444_cse : STD_LOGIC;
  SIGNAL or_493_cse : STD_LOGIC;
  SIGNAL or_701_cse : STD_LOGIC;
  SIGNAL nand_394_cse : STD_LOGIC;
  SIGNAL or_1113_cse : STD_LOGIC;
  SIGNAL nand_356_cse : STD_LOGIC;
  SIGNAL nand_336_cse : STD_LOGIC;
  SIGNAL nand_300_cse : STD_LOGIC;
  SIGNAL nand_293_cse : STD_LOGIC;
  SIGNAL nand_264_cse : STD_LOGIC;
  SIGNAL nand_204_cse : STD_LOGIC;
  SIGNAL nand_205_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_0_31_obj_ld_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL or_220_cse : STD_LOGIC;
  SIGNAL or_212_cse : STD_LOGIC;
  SIGNAL and_496_cse : STD_LOGIC;
  SIGNAL and_316_cse : STD_LOGIC;
  SIGNAL or_32_cse : STD_LOGIC;
  SIGNAL mux_189_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_12_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_17_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_35_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_40_cse : STD_LOGIC;
  SIGNAL and_4_cse : STD_LOGIC;
  SIGNAL and_1_cse : STD_LOGIC;
  SIGNAL nor_1025_cse : STD_LOGIC;
  SIGNAL and_464_cse : STD_LOGIC;
  SIGNAL and_490_cse : STD_LOGIC;
  SIGNAL and_449_cse : STD_LOGIC;
  SIGNAL and_479_cse : STD_LOGIC;
  SIGNAL mux_322_cse : STD_LOGIC;
  SIGNAL nand_445_cse : STD_LOGIC;
  SIGNAL nand_447_cse : STD_LOGIC;
  SIGNAL nand_441_cse : STD_LOGIC;
  SIGNAL nand_442_cse : STD_LOGIC;
  SIGNAL mux_353_cse : STD_LOGIC;
  SIGNAL nand_446_cse : STD_LOGIC;
  SIGNAL nand_448_cse : STD_LOGIC;
  SIGNAL nor_98_cse : STD_LOGIC;
  SIGNAL mux_446_cse : STD_LOGIC;
  SIGNAL nand_423_cse : STD_LOGIC;
  SIGNAL mux_477_cse : STD_LOGIC;
  SIGNAL mux_570_cse : STD_LOGIC;
  SIGNAL nand_435_cse : STD_LOGIC;
  SIGNAL nand_411_cse : STD_LOGIC;
  SIGNAL nand_437_cse : STD_LOGIC;
  SIGNAL mux_601_cse : STD_LOGIC;
  SIGNAL mux_694_cse : STD_LOGIC;
  SIGNAL nand_371_cse : STD_LOGIC;
  SIGNAL nand_385_cse : STD_LOGIC;
  SIGNAL mux_725_cse : STD_LOGIC;
  SIGNAL nand_364_cse : STD_LOGIC;
  SIGNAL nand_365_cse : STD_LOGIC;
  SIGNAL nand_357_cse : STD_LOGIC;
  SIGNAL nand_353_cse : STD_LOGIC;
  SIGNAL nand_417_cse : STD_LOGIC;
  SIGNAL nand_419_cse : STD_LOGIC;
  SIGNAL nand_302_cse : STD_LOGIC;
  SIGNAL nand_303_cse : STD_LOGIC;
  SIGNAL nand_294_cse : STD_LOGIC;
  SIGNAL nand_289_cse : STD_LOGIC;
  SIGNAL nand_266_cse : STD_LOGIC;
  SIGNAL nand_297_cse : STD_LOGIC;
  SIGNAL mux_1190_cse : STD_LOGIC;
  SIGNAL mux_1221_cse : STD_LOGIC;
  SIGNAL or_167_cse : STD_LOGIC;
  SIGNAL or_145_cse : STD_LOGIC;
  SIGNAL nor_1023_cse : STD_LOGIC;
  SIGNAL and_491_cse : STD_LOGIC;
  SIGNAL and_485_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm : STD_LOGIC;
  SIGNAL mux_348_cse : STD_LOGIC;
  SIGNAL mux_410_cse : STD_LOGIC;
  SIGNAL mux_472_cse : STD_LOGIC;
  SIGNAL mux_534_cse : STD_LOGIC;
  SIGNAL mux_596_cse : STD_LOGIC;
  SIGNAL mux_658_cse : STD_LOGIC;
  SIGNAL mux_720_cse : STD_LOGIC;
  SIGNAL mux_782_cse : STD_LOGIC;
  SIGNAL mux_844_cse : STD_LOGIC;
  SIGNAL mux_818_cse : STD_LOGIC;
  SIGNAL mux_849_cse : STD_LOGIC;
  SIGNAL mux_906_cse : STD_LOGIC;
  SIGNAL mux_968_cse : STD_LOGIC;
  SIGNAL mux_942_cse : STD_LOGIC;
  SIGNAL mux_973_cse : STD_LOGIC;
  SIGNAL mux_1030_cse : STD_LOGIC;
  SIGNAL mux_1092_cse : STD_LOGIC;
  SIGNAL mux_1066_cse : STD_LOGIC;
  SIGNAL mux_1097_cse : STD_LOGIC;
  SIGNAL mux_1154_cse : STD_LOGIC;
  SIGNAL mux_1216_cse : STD_LOGIC;
  SIGNAL mux_1278_cse : STD_LOGIC;
  SIGNAL and_33_cse : STD_LOGIC;
  SIGNAL and_456_cse : STD_LOGIC;
  SIGNAL mux_1462_rmff : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_8_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_1_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_2_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_3_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_4_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_5_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_6_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_1489_itm : STD_LOGIC;
  SIGNAL mux_1531_itm : STD_LOGIC;
  SIGNAL mux_1536_itm : STD_LOGIC;
  SIGNAL mux_1538_itm : STD_LOGIC;
  SIGNAL mux_1543_itm : STD_LOGIC;
  SIGNAL z_out : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL and_dcpl_334 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL and_dcpl_347 : STD_LOGIC;
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_dcpl_353 : STD_LOGIC;
  SIGNAL and_dcpl_365 : STD_LOGIC;
  SIGNAL and_dcpl_372 : STD_LOGIC;
  SIGNAL and_dcpl_419 : STD_LOGIC;
  SIGNAL and_dcpl_420 : STD_LOGIC;
  SIGNAL and_dcpl_422 : STD_LOGIC;
  SIGNAL and_dcpl_423 : STD_LOGIC;
  SIGNAL and_dcpl_425 : STD_LOGIC;
  SIGNAL and_dcpl_428 : STD_LOGIC;
  SIGNAL and_dcpl_429 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL and_dcpl_434 : STD_LOGIC;
  SIGNAL and_dcpl_435 : STD_LOGIC;
  SIGNAL and_dcpl_436 : STD_LOGIC;
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_448 : STD_LOGIC;
  SIGNAL and_dcpl_452 : STD_LOGIC;
  SIGNAL and_dcpl_456 : STD_LOGIC;
  SIGNAL and_dcpl_458 : STD_LOGIC;
  SIGNAL and_dcpl_461 : STD_LOGIC;
  SIGNAL and_dcpl_465 : STD_LOGIC;
  SIGNAL and_dcpl_468 : STD_LOGIC;
  SIGNAL and_dcpl_472 : STD_LOGIC;
  SIGNAL z_out_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_dcpl_479 : STD_LOGIC;
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_acc_cse_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tmp_21_sva_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_11 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_13 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_14 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_15 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_17 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_18 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_19 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_21 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_22 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_23 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_25 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_26 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_27 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_29 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_30 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_31 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_18_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_20_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_21_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_22_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_23_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_24_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_25_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_26_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_27_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_28_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_29_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_30_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_126_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_128_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_129_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_130_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_132_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_133_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_134_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_136_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_141_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_142_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_144_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_126_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_127_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_157_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_129_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_159_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_160_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_161_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_133_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_163_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_164_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_165_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_166_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_167_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_168_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_169_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_171_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_172_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_173_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_174_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_175_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_176_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_177_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_178_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_179_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_180_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_181_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_182_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_183_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_184_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_185_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_3_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_226_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_227_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_281_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_229_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_283_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_284_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_285_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_233_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_287_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_288_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_289_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_290_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_291_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_292_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_293_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_240_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_295_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_296_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_297_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_298_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_299_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_300_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_301_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_302_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_303_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_304_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_305_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_306_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_307_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_308_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_309_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_26_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_28_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_31_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_377_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_326_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_327_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_405_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_329_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_407_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_408_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_409_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_333_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_411_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_412_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_413_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_414_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_415_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_416_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_417_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_340_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_419_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_420_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_421_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_422_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_423_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_424_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_425_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_426_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_427_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_428_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_429_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_430_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_431_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_432_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_433_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_17_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_426_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_427_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_529_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_429_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_531_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_532_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_533_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_433_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_535_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_536_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_537_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_538_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_539_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_540_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_541_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_440_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_543_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_544_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_545_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_546_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_547_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_548_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_549_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_550_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_551_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_552_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_553_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_554_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_555_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_556_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_557_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_625_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_21_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_526_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_527_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_653_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_529_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_655_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_656_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_657_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_533_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_659_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_660_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_661_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_662_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_663_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_664_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_665_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_540_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_667_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_668_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_669_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_670_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_671_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_672_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_673_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_674_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_675_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_676_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_677_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_678_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_679_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_680_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_681_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_25_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_626_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_627_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_777_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_629_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_779_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_780_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_781_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_633_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_783_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_784_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_785_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_786_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_787_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_788_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_789_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_640_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_791_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_792_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_793_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_794_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_795_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_796_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_797_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_798_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_799_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_800_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_801_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_802_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_803_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_804_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_805_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_29_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_726_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_727_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_901_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_729_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_903_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_904_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_905_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_733_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_907_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_908_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_909_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_910_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_911_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_912_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_913_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_740_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_915_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_916_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_917_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_918_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_919_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_920_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_921_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_922_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_923_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_924_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_925_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_926_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_927_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_928_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_929_itm : STD_LOGIC;
  SIGNAL STAGE_LOOP_i_3_0_sva_mx0c1 : STD_LOGIC;
  SIGNAL VEC_LOOP_j_10_0_sva_9_0_mx0c0 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_itm_mx0c0 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_itm_mx0c1 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_itm_mx0c2 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_itm_mx0c3 : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_8_itm_mx0c4 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_165 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 : STD_LOGIC;
  SIGNAL COMP_LOOP_3_tmp_mul_idiv_sva_3_0 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_or_59_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_27_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_29_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_30_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_32_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_33_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_34_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_1_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_41_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_101_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_105_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_35_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_39_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_78_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_79_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_81_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_42_cse : STD_LOGIC;
  SIGNAL nor_489_cse : STD_LOGIC;
  SIGNAL nor_480_cse : STD_LOGIC;
  SIGNAL nor_479_cse : STD_LOGIC;
  SIGNAL nor_461_cse : STD_LOGIC;
  SIGNAL nor_460_cse : STD_LOGIC;
  SIGNAL nor_450_cse : STD_LOGIC;
  SIGNAL nor_441_cse : STD_LOGIC;
  SIGNAL nor_440_cse : STD_LOGIC;
  SIGNAL nor_422_cse : STD_LOGIC;
  SIGNAL nor_421_cse : STD_LOGIC;
  SIGNAL nor_411_cse : STD_LOGIC;
  SIGNAL nor_402_cse : STD_LOGIC;
  SIGNAL nor_401_cse : STD_LOGIC;
  SIGNAL nor_383_cse : STD_LOGIC;
  SIGNAL nor_382_cse : STD_LOGIC;
  SIGNAL nor_372_cse : STD_LOGIC;
  SIGNAL nor_363_cse : STD_LOGIC;
  SIGNAL nor_362_cse : STD_LOGIC;
  SIGNAL nor_347_cse : STD_LOGIC;
  SIGNAL and_325_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse : STD_LOGIC;
  SIGNAL and_628_cse : STD_LOGIC;
  SIGNAL and_605_cse : STD_LOGIC;
  SIGNAL and_609_cse : STD_LOGIC;
  SIGNAL and_614_cse : STD_LOGIC;
  SIGNAL and_617_cse : STD_LOGIC;
  SIGNAL and_621_cse : STD_LOGIC;
  SIGNAL and_624_cse : STD_LOGIC;
  SIGNAL or_tmp_2098 : STD_LOGIC;
  SIGNAL mux_tmp_1564 : STD_LOGIC;
  SIGNAL COMP_LOOP_or_36_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_33_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_71_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_2_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_3_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_4_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_5_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_6_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_7_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_8_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_or_54_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_385_cse : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_135_cse : STD_LOGIC;

  SIGNAL nor_1019_nl : STD_LOGIC;
  SIGNAL mux_320_nl : STD_LOGIC;
  SIGNAL mux_347_nl : STD_LOGIC;
  SIGNAL nand_11_nl : STD_LOGIC;
  SIGNAL nand_22_nl : STD_LOGIC;
  SIGNAL mux_409_nl : STD_LOGIC;
  SIGNAL mux_471_nl : STD_LOGIC;
  SIGNAL nand_33_nl : STD_LOGIC;
  SIGNAL nand_44_nl : STD_LOGIC;
  SIGNAL mux_533_nl : STD_LOGIC;
  SIGNAL mux_595_nl : STD_LOGIC;
  SIGNAL nand_55_nl : STD_LOGIC;
  SIGNAL nand_66_nl : STD_LOGIC;
  SIGNAL mux_657_nl : STD_LOGIC;
  SIGNAL mux_719_nl : STD_LOGIC;
  SIGNAL nand_77_nl : STD_LOGIC;
  SIGNAL nand_88_nl : STD_LOGIC;
  SIGNAL mux_781_nl : STD_LOGIC;
  SIGNAL or_1066_nl : STD_LOGIC;
  SIGNAL or_1064_nl : STD_LOGIC;
  SIGNAL mux_843_nl : STD_LOGIC;
  SIGNAL nand_99_nl : STD_LOGIC;
  SIGNAL nor_730_nl : STD_LOGIC;
  SIGNAL nor_731_nl : STD_LOGIC;
  SIGNAL nand_110_nl : STD_LOGIC;
  SIGNAL mux_905_nl : STD_LOGIC;
  SIGNAL or_1274_nl : STD_LOGIC;
  SIGNAL or_1272_nl : STD_LOGIC;
  SIGNAL mux_967_nl : STD_LOGIC;
  SIGNAL nand_121_nl : STD_LOGIC;
  SIGNAL nor_662_nl : STD_LOGIC;
  SIGNAL nor_663_nl : STD_LOGIC;
  SIGNAL nand_132_nl : STD_LOGIC;
  SIGNAL mux_1029_nl : STD_LOGIC;
  SIGNAL or_1481_nl : STD_LOGIC;
  SIGNAL or_1480_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL nand_143_nl : STD_LOGIC;
  SIGNAL nor_595_nl : STD_LOGIC;
  SIGNAL nor_596_nl : STD_LOGIC;
  SIGNAL nand_154_nl : STD_LOGIC;
  SIGNAL mux_1153_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL nand_165_nl : STD_LOGIC;
  SIGNAL nand_176_nl : STD_LOGIC;
  SIGNAL mux_1277_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_j_not_1_nl : STD_LOGIC;
  SIGNAL nor_1160_nl : STD_LOGIC;
  SIGNAL and_nl : STD_LOGIC;
  SIGNAL nand_nl : STD_LOGIC;
  SIGNAL mux_312_nl : STD_LOGIC;
  SIGNAL nor_1021_nl : STD_LOGIC;
  SIGNAL and_451_nl : STD_LOGIC;
  SIGNAL mux_1604_nl : STD_LOGIC;
  SIGNAL or_2285_nl : STD_LOGIC;
  SIGNAL mux_1603_nl : STD_LOGIC;
  SIGNAL or_2284_nl : STD_LOGIC;
  SIGNAL mux_1602_nl : STD_LOGIC;
  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL or_nl : STD_LOGIC;
  SIGNAL mux_1492_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL mux_1499_nl : STD_LOGIC;
  SIGNAL mux_1498_nl : STD_LOGIC;
  SIGNAL and_260_nl : STD_LOGIC;
  SIGNAL mux_1500_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_3_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL and_310_nl : STD_LOGIC;
  SIGNAL mux_1505_nl : STD_LOGIC;
  SIGNAL mux_1504_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL mux_1506_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_12_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_5_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_1513_nl : STD_LOGIC;
  SIGNAL mux_1512_nl : STD_LOGIC;
  SIGNAL mux_1518_nl : STD_LOGIC;
  SIGNAL mux_1520_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_6_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_1523_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_7_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_1528_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL or_162_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_15_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL and_305_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL and_304_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_33_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_35_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_36_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_37_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_39_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_40_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_41_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_42_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_43_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_44_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_45_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_47_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_48_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_49_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_50_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_51_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_52_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_53_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_54_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_55_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_56_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_57_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_58_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_59_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_60_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_61_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_33_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_40_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_17_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_mux_2_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_or_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_23_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_24_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_25_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_28_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_30_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_31_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_127_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_128_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_129_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_130_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_131_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_132_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_133_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_134_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_135_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_136_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_137_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_138_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_139_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_140_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_141_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_142_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_143_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_144_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_145_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_146_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_147_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_148_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_149_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_150_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_151_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_152_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_153_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_154_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_155_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_115_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_116_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_117_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_118_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_119_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_120_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_121_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_122_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_123_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_124_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_125_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_126_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_83_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_84_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_85_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_86_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_87_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_88_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_89_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_90_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_91_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_92_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_93_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_94_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_95_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_96_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_97_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_98_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_99_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_100_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_101_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_102_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_103_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_104_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_105_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_106_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_107_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_108_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_109_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_110_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_111_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_112_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_113_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_114_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_78_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_79_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_80_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_81_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_82_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_47_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_48_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_49_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_50_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_51_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_52_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_53_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_54_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_55_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_56_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_57_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_58_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_59_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_60_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_61_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_62_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_63_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_64_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_65_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_66_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_67_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_68_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_69_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_70_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_71_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_72_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_73_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_74_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_75_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_76_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_77_nl : STD_LOGIC;
  SIGNAL mux_1585_nl : STD_LOGIC;
  SIGNAL mux_1584_nl : STD_LOGIC;
  SIGNAL mux_1583_nl : STD_LOGIC;
  SIGNAL nor_337_nl : STD_LOGIC;
  SIGNAL mux_1582_nl : STD_LOGIC;
  SIGNAL mux_1591_nl : STD_LOGIC;
  SIGNAL mux_1590_nl : STD_LOGIC;
  SIGNAL mux_1589_nl : STD_LOGIC;
  SIGNAL mux_1588_nl : STD_LOGIC;
  SIGNAL mux_1587_nl : STD_LOGIC;
  SIGNAL mux_1586_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_23_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_24_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_25_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_28_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_30_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_31_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_32_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_33_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_34_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_35_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_36_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_37_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_38_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_39_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_40_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_41_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_42_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_43_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_44_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_45_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_46_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_14_nl : STD_LOGIC;
  SIGNAL mux_1597_nl : STD_LOGIC;
  SIGNAL mux_1596_nl : STD_LOGIC;
  SIGNAL mux_1595_nl : STD_LOGIC;
  SIGNAL mux_1594_nl : STD_LOGIC;
  SIGNAL mux_217_nl : STD_LOGIC;
  SIGNAL and_478_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_2_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_3_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_4_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_5_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_6_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_7_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_8_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL or_238_nl : STD_LOGIC;
  SIGNAL or_236_nl : STD_LOGIC;
  SIGNAL or_284_nl : STD_LOGIC;
  SIGNAL or_282_nl : STD_LOGIC;
  SIGNAL nor_1001_nl : STD_LOGIC;
  SIGNAL nor_1002_nl : STD_LOGIC;
  SIGNAL or_388_nl : STD_LOGIC;
  SIGNAL or_386_nl : STD_LOGIC;
  SIGNAL or_446_nl : STD_LOGIC;
  SIGNAL or_444_nl : STD_LOGIC;
  SIGNAL or_492_nl : STD_LOGIC;
  SIGNAL or_490_nl : STD_LOGIC;
  SIGNAL nor_933_nl : STD_LOGIC;
  SIGNAL nor_934_nl : STD_LOGIC;
  SIGNAL or_596_nl : STD_LOGIC;
  SIGNAL or_594_nl : STD_LOGIC;
  SIGNAL or_654_nl : STD_LOGIC;
  SIGNAL or_652_nl : STD_LOGIC;
  SIGNAL or_700_nl : STD_LOGIC;
  SIGNAL or_698_nl : STD_LOGIC;
  SIGNAL nor_865_nl : STD_LOGIC;
  SIGNAL nor_866_nl : STD_LOGIC;
  SIGNAL or_804_nl : STD_LOGIC;
  SIGNAL or_802_nl : STD_LOGIC;
  SIGNAL nand_518_nl : STD_LOGIC;
  SIGNAL or_860_nl : STD_LOGIC;
  SIGNAL or_908_nl : STD_LOGIC;
  SIGNAL or_906_nl : STD_LOGIC;
  SIGNAL and_532_nl : STD_LOGIC;
  SIGNAL nor_798_nl : STD_LOGIC;
  SIGNAL nand_472_nl : STD_LOGIC;
  SIGNAL or_1009_nl : STD_LOGIC;
  SIGNAL or_1112_nl : STD_LOGIC;
  SIGNAL or_1110_nl : STD_LOGIC;
  SIGNAL or_1216_nl : STD_LOGIC;
  SIGNAL or_1214_nl : STD_LOGIC;
  SIGNAL or_1320_nl : STD_LOGIC;
  SIGNAL or_1318_nl : STD_LOGIC;
  SIGNAL nand_469_nl : STD_LOGIC;
  SIGNAL or_1422_nl : STD_LOGIC;
  SIGNAL or_1527_nl : STD_LOGIC;
  SIGNAL or_1525_nl : STD_LOGIC;
  SIGNAL nand_466_nl : STD_LOGIC;
  SIGNAL or_1627_nl : STD_LOGIC;
  SIGNAL nand_268_nl : STD_LOGIC;
  SIGNAL nand_269_nl : STD_LOGIC;
  SIGNAL nand_463_nl : STD_LOGIC;
  SIGNAL or_1727_nl : STD_LOGIC;
  SIGNAL and_353_nl : STD_LOGIC;
  SIGNAL and_354_nl : STD_LOGIC;
  SIGNAL nand_459_nl : STD_LOGIC;
  SIGNAL nand_236_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL mux_240_nl : STD_LOGIC;
  SIGNAL or_2109_nl : STD_LOGIC;
  SIGNAL mux_1488_nl : STD_LOGIC;
  SIGNAL mux_1486_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL and_448_nl : STD_LOGIC;
  SIGNAL mux_1606_nl : STD_LOGIC;
  SIGNAL nor_340_nl : STD_LOGIC;
  SIGNAL and_511_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL nand_188_nl : STD_LOGIC;
  SIGNAL mux_1515_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL mux_1599_nl : STD_LOGIC;
  SIGNAL and_446_nl : STD_LOGIC;
  SIGNAL mux_1526_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL mux_1535_nl : STD_LOGIC;
  SIGNAL and_306_nl : STD_LOGIC;
  SIGNAL mux_1537_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL mux_1551_nl : STD_LOGIC;
  SIGNAL nor_1128_nl : STD_LOGIC;
  SIGNAL nor_1129_nl : STD_LOGIC;
  SIGNAL mux_1555_nl : STD_LOGIC;
  SIGNAL mux_1554_nl : STD_LOGIC;
  SIGNAL mux_1553_nl : STD_LOGIC;
  SIGNAL nand_185_nl : STD_LOGIC;
  SIGNAL mux_1552_nl : STD_LOGIC;
  SIGNAL nand_473_nl : STD_LOGIC;
  SIGNAL or_2171_nl : STD_LOGIC;
  SIGNAL mux_1575_nl : STD_LOGIC;
  SIGNAL mux_1574_nl : STD_LOGIC;
  SIGNAL or_229_nl : STD_LOGIC;
  SIGNAL mux_1573_nl : STD_LOGIC;
  SIGNAL mux_1579_nl : STD_LOGIC;
  SIGNAL mux_1578_nl : STD_LOGIC;
  SIGNAL mux_1577_nl : STD_LOGIC;
  SIGNAL mux_1576_nl : STD_LOGIC;
  SIGNAL nor_1059_nl : STD_LOGIC;
  SIGNAL mux_1581_nl : STD_LOGIC;
  SIGNAL mux_1580_nl : STD_LOGIC;
  SIGNAL nor_1062_nl : STD_LOGIC;
  SIGNAL nor_1063_nl : STD_LOGIC;
  SIGNAL and_520_nl : STD_LOGIC;
  SIGNAL and_54_nl : STD_LOGIC;
  SIGNAL and_64_nl : STD_LOGIC;
  SIGNAL and_68_nl : STD_LOGIC;
  SIGNAL and_74_nl : STD_LOGIC;
  SIGNAL and_78_nl : STD_LOGIC;
  SIGNAL and_84_nl : STD_LOGIC;
  SIGNAL and_88_nl : STD_LOGIC;
  SIGNAL and_92_nl : STD_LOGIC;
  SIGNAL and_95_nl : STD_LOGIC;
  SIGNAL and_97_nl : STD_LOGIC;
  SIGNAL and_98_nl : STD_LOGIC;
  SIGNAL and_99_nl : STD_LOGIC;
  SIGNAL and_101_nl : STD_LOGIC;
  SIGNAL and_103_nl : STD_LOGIC;
  SIGNAL and_104_nl : STD_LOGIC;
  SIGNAL and_105_nl : STD_LOGIC;
  SIGNAL and_107_nl : STD_LOGIC;
  SIGNAL and_109_nl : STD_LOGIC;
  SIGNAL and_110_nl : STD_LOGIC;
  SIGNAL and_111_nl : STD_LOGIC;
  SIGNAL and_112_nl : STD_LOGIC;
  SIGNAL and_114_nl : STD_LOGIC;
  SIGNAL and_116_nl : STD_LOGIC;
  SIGNAL and_117_nl : STD_LOGIC;
  SIGNAL mux_336_nl : STD_LOGIC;
  SIGNAL nand_506_nl : STD_LOGIC;
  SIGNAL mux_335_nl : STD_LOGIC;
  SIGNAL and_443_nl : STD_LOGIC;
  SIGNAL mux_334_nl : STD_LOGIC;
  SIGNAL mux_333_nl : STD_LOGIC;
  SIGNAL nor_1010_nl : STD_LOGIC;
  SIGNAL nor_1011_nl : STD_LOGIC;
  SIGNAL mux_332_nl : STD_LOGIC;
  SIGNAL nor_1012_nl : STD_LOGIC;
  SIGNAL nor_1013_nl : STD_LOGIC;
  SIGNAL nor_1014_nl : STD_LOGIC;
  SIGNAL mux_331_nl : STD_LOGIC;
  SIGNAL mux_330_nl : STD_LOGIC;
  SIGNAL or_257_nl : STD_LOGIC;
  SIGNAL or_255_nl : STD_LOGIC;
  SIGNAL mux_329_nl : STD_LOGIC;
  SIGNAL or_254_nl : STD_LOGIC;
  SIGNAL or_252_nl : STD_LOGIC;
  SIGNAL or_2280_nl : STD_LOGIC;
  SIGNAL mux_328_nl : STD_LOGIC;
  SIGNAL nand_8_nl : STD_LOGIC;
  SIGNAL mux_327_nl : STD_LOGIC;
  SIGNAL mux_326_nl : STD_LOGIC;
  SIGNAL nor_1016_nl : STD_LOGIC;
  SIGNAL nor_1017_nl : STD_LOGIC;
  SIGNAL nor_1018_nl : STD_LOGIC;
  SIGNAL mux_325_nl : STD_LOGIC;
  SIGNAL or_246_nl : STD_LOGIC;
  SIGNAL or_244_nl : STD_LOGIC;
  SIGNAL or_243_nl : STD_LOGIC;
  SIGNAL mux_324_nl : STD_LOGIC;
  SIGNAL mux_323_nl : STD_LOGIC;
  SIGNAL or_242_nl : STD_LOGIC;
  SIGNAL or_240_nl : STD_LOGIC;
  SIGNAL or_239_nl : STD_LOGIC;
  SIGNAL mux_352_nl : STD_LOGIC;
  SIGNAL mux_351_nl : STD_LOGIC;
  SIGNAL mux_350_nl : STD_LOGIC;
  SIGNAL nor_1003_nl : STD_LOGIC;
  SIGNAL nor_1004_nl : STD_LOGIC;
  SIGNAL mux_349_nl : STD_LOGIC;
  SIGNAL nor_1005_nl : STD_LOGIC;
  SIGNAL mux_345_nl : STD_LOGIC;
  SIGNAL nor_1006_nl : STD_LOGIC;
  SIGNAL mux_344_nl : STD_LOGIC;
  SIGNAL nor_1007_nl : STD_LOGIC;
  SIGNAL nor_1008_nl : STD_LOGIC;
  SIGNAL nor_1009_nl : STD_LOGIC;
  SIGNAL mux_343_nl : STD_LOGIC;
  SIGNAL mux_342_nl : STD_LOGIC;
  SIGNAL mux_341_nl : STD_LOGIC;
  SIGNAL or_276_nl : STD_LOGIC;
  SIGNAL or_274_nl : STD_LOGIC;
  SIGNAL mux_340_nl : STD_LOGIC;
  SIGNAL or_273_nl : STD_LOGIC;
  SIGNAL or_271_nl : STD_LOGIC;
  SIGNAL mux_339_nl : STD_LOGIC;
  SIGNAL mux_338_nl : STD_LOGIC;
  SIGNAL or_270_nl : STD_LOGIC;
  SIGNAL or_268_nl : STD_LOGIC;
  SIGNAL mux_337_nl : STD_LOGIC;
  SIGNAL or_267_nl : STD_LOGIC;
  SIGNAL or_265_nl : STD_LOGIC;
  SIGNAL mux_367_nl : STD_LOGIC;
  SIGNAL nand_505_nl : STD_LOGIC;
  SIGNAL mux_366_nl : STD_LOGIC;
  SIGNAL and_440_nl : STD_LOGIC;
  SIGNAL mux_365_nl : STD_LOGIC;
  SIGNAL mux_364_nl : STD_LOGIC;
  SIGNAL nor_991_nl : STD_LOGIC;
  SIGNAL nor_992_nl : STD_LOGIC;
  SIGNAL mux_363_nl : STD_LOGIC;
  SIGNAL nor_993_nl : STD_LOGIC;
  SIGNAL nor_994_nl : STD_LOGIC;
  SIGNAL nor_995_nl : STD_LOGIC;
  SIGNAL mux_362_nl : STD_LOGIC;
  SIGNAL mux_361_nl : STD_LOGIC;
  SIGNAL or_308_nl : STD_LOGIC;
  SIGNAL or_306_nl : STD_LOGIC;
  SIGNAL mux_360_nl : STD_LOGIC;
  SIGNAL or_305_nl : STD_LOGIC;
  SIGNAL or_303_nl : STD_LOGIC;
  SIGNAL or_2279_nl : STD_LOGIC;
  SIGNAL mux_359_nl : STD_LOGIC;
  SIGNAL nand_14_nl : STD_LOGIC;
  SIGNAL mux_358_nl : STD_LOGIC;
  SIGNAL mux_357_nl : STD_LOGIC;
  SIGNAL nor_997_nl : STD_LOGIC;
  SIGNAL nor_998_nl : STD_LOGIC;
  SIGNAL and_441_nl : STD_LOGIC;
  SIGNAL mux_356_nl : STD_LOGIC;
  SIGNAL nor_999_nl : STD_LOGIC;
  SIGNAL nor_1000_nl : STD_LOGIC;
  SIGNAL or_295_nl : STD_LOGIC;
  SIGNAL mux_355_nl : STD_LOGIC;
  SIGNAL mux_354_nl : STD_LOGIC;
  SIGNAL or_294_nl : STD_LOGIC;
  SIGNAL or_292_nl : STD_LOGIC;
  SIGNAL nand_12_nl : STD_LOGIC;
  SIGNAL mux_383_nl : STD_LOGIC;
  SIGNAL mux_382_nl : STD_LOGIC;
  SIGNAL mux_381_nl : STD_LOGIC;
  SIGNAL nor_985_nl : STD_LOGIC;
  SIGNAL nor_986_nl : STD_LOGIC;
  SIGNAL mux_380_nl : STD_LOGIC;
  SIGNAL and_438_nl : STD_LOGIC;
  SIGNAL mux_376_nl : STD_LOGIC;
  SIGNAL nor_987_nl : STD_LOGIC;
  SIGNAL mux_375_nl : STD_LOGIC;
  SIGNAL nor_988_nl : STD_LOGIC;
  SIGNAL nor_989_nl : STD_LOGIC;
  SIGNAL nor_990_nl : STD_LOGIC;
  SIGNAL mux_374_nl : STD_LOGIC;
  SIGNAL mux_373_nl : STD_LOGIC;
  SIGNAL mux_372_nl : STD_LOGIC;
  SIGNAL or_327_nl : STD_LOGIC;
  SIGNAL or_325_nl : STD_LOGIC;
  SIGNAL mux_371_nl : STD_LOGIC;
  SIGNAL or_324_nl : STD_LOGIC;
  SIGNAL or_322_nl : STD_LOGIC;
  SIGNAL mux_370_nl : STD_LOGIC;
  SIGNAL mux_369_nl : STD_LOGIC;
  SIGNAL or_321_nl : STD_LOGIC;
  SIGNAL or_319_nl : STD_LOGIC;
  SIGNAL mux_368_nl : STD_LOGIC;
  SIGNAL or_318_nl : STD_LOGIC;
  SIGNAL or_316_nl : STD_LOGIC;
  SIGNAL mux_398_nl : STD_LOGIC;
  SIGNAL nand_504_nl : STD_LOGIC;
  SIGNAL mux_397_nl : STD_LOGIC;
  SIGNAL and_437_nl : STD_LOGIC;
  SIGNAL mux_396_nl : STD_LOGIC;
  SIGNAL mux_395_nl : STD_LOGIC;
  SIGNAL nor_976_nl : STD_LOGIC;
  SIGNAL nor_977_nl : STD_LOGIC;
  SIGNAL mux_394_nl : STD_LOGIC;
  SIGNAL nor_978_nl : STD_LOGIC;
  SIGNAL nor_979_nl : STD_LOGIC;
  SIGNAL nor_980_nl : STD_LOGIC;
  SIGNAL mux_393_nl : STD_LOGIC;
  SIGNAL mux_392_nl : STD_LOGIC;
  SIGNAL or_361_nl : STD_LOGIC;
  SIGNAL or_359_nl : STD_LOGIC;
  SIGNAL mux_391_nl : STD_LOGIC;
  SIGNAL or_358_nl : STD_LOGIC;
  SIGNAL or_356_nl : STD_LOGIC;
  SIGNAL or_2278_nl : STD_LOGIC;
  SIGNAL mux_390_nl : STD_LOGIC;
  SIGNAL nand_19_nl : STD_LOGIC;
  SIGNAL mux_389_nl : STD_LOGIC;
  SIGNAL mux_388_nl : STD_LOGIC;
  SIGNAL nor_982_nl : STD_LOGIC;
  SIGNAL nor_983_nl : STD_LOGIC;
  SIGNAL nor_984_nl : STD_LOGIC;
  SIGNAL mux_387_nl : STD_LOGIC;
  SIGNAL or_350_nl : STD_LOGIC;
  SIGNAL or_348_nl : STD_LOGIC;
  SIGNAL or_347_nl : STD_LOGIC;
  SIGNAL mux_386_nl : STD_LOGIC;
  SIGNAL mux_385_nl : STD_LOGIC;
  SIGNAL or_346_nl : STD_LOGIC;
  SIGNAL or_344_nl : STD_LOGIC;
  SIGNAL or_343_nl : STD_LOGIC;
  SIGNAL mux_414_nl : STD_LOGIC;
  SIGNAL mux_413_nl : STD_LOGIC;
  SIGNAL mux_412_nl : STD_LOGIC;
  SIGNAL nor_969_nl : STD_LOGIC;
  SIGNAL nor_970_nl : STD_LOGIC;
  SIGNAL mux_411_nl : STD_LOGIC;
  SIGNAL nor_971_nl : STD_LOGIC;
  SIGNAL mux_407_nl : STD_LOGIC;
  SIGNAL nor_972_nl : STD_LOGIC;
  SIGNAL mux_406_nl : STD_LOGIC;
  SIGNAL nor_973_nl : STD_LOGIC;
  SIGNAL nor_974_nl : STD_LOGIC;
  SIGNAL nor_975_nl : STD_LOGIC;
  SIGNAL mux_405_nl : STD_LOGIC;
  SIGNAL mux_404_nl : STD_LOGIC;
  SIGNAL mux_403_nl : STD_LOGIC;
  SIGNAL or_380_nl : STD_LOGIC;
  SIGNAL or_378_nl : STD_LOGIC;
  SIGNAL mux_402_nl : STD_LOGIC;
  SIGNAL or_377_nl : STD_LOGIC;
  SIGNAL or_375_nl : STD_LOGIC;
  SIGNAL mux_401_nl : STD_LOGIC;
  SIGNAL mux_400_nl : STD_LOGIC;
  SIGNAL or_374_nl : STD_LOGIC;
  SIGNAL or_372_nl : STD_LOGIC;
  SIGNAL mux_399_nl : STD_LOGIC;
  SIGNAL or_371_nl : STD_LOGIC;
  SIGNAL or_369_nl : STD_LOGIC;
  SIGNAL mux_429_nl : STD_LOGIC;
  SIGNAL nand_503_nl : STD_LOGIC;
  SIGNAL mux_428_nl : STD_LOGIC;
  SIGNAL and_434_nl : STD_LOGIC;
  SIGNAL mux_427_nl : STD_LOGIC;
  SIGNAL mux_426_nl : STD_LOGIC;
  SIGNAL nor_957_nl : STD_LOGIC;
  SIGNAL nor_958_nl : STD_LOGIC;
  SIGNAL mux_425_nl : STD_LOGIC;
  SIGNAL nor_959_nl : STD_LOGIC;
  SIGNAL nor_960_nl : STD_LOGIC;
  SIGNAL nor_961_nl : STD_LOGIC;
  SIGNAL mux_424_nl : STD_LOGIC;
  SIGNAL mux_423_nl : STD_LOGIC;
  SIGNAL or_412_nl : STD_LOGIC;
  SIGNAL or_410_nl : STD_LOGIC;
  SIGNAL mux_422_nl : STD_LOGIC;
  SIGNAL or_409_nl : STD_LOGIC;
  SIGNAL or_407_nl : STD_LOGIC;
  SIGNAL or_2277_nl : STD_LOGIC;
  SIGNAL mux_421_nl : STD_LOGIC;
  SIGNAL nand_25_nl : STD_LOGIC;
  SIGNAL mux_420_nl : STD_LOGIC;
  SIGNAL mux_419_nl : STD_LOGIC;
  SIGNAL nor_963_nl : STD_LOGIC;
  SIGNAL nor_964_nl : STD_LOGIC;
  SIGNAL and_435_nl : STD_LOGIC;
  SIGNAL mux_418_nl : STD_LOGIC;
  SIGNAL nor_965_nl : STD_LOGIC;
  SIGNAL nor_966_nl : STD_LOGIC;
  SIGNAL or_399_nl : STD_LOGIC;
  SIGNAL mux_417_nl : STD_LOGIC;
  SIGNAL mux_416_nl : STD_LOGIC;
  SIGNAL or_398_nl : STD_LOGIC;
  SIGNAL or_396_nl : STD_LOGIC;
  SIGNAL nand_23_nl : STD_LOGIC;
  SIGNAL mux_445_nl : STD_LOGIC;
  SIGNAL mux_444_nl : STD_LOGIC;
  SIGNAL mux_443_nl : STD_LOGIC;
  SIGNAL nor_951_nl : STD_LOGIC;
  SIGNAL nor_952_nl : STD_LOGIC;
  SIGNAL mux_442_nl : STD_LOGIC;
  SIGNAL and_432_nl : STD_LOGIC;
  SIGNAL mux_438_nl : STD_LOGIC;
  SIGNAL nor_953_nl : STD_LOGIC;
  SIGNAL mux_437_nl : STD_LOGIC;
  SIGNAL nor_954_nl : STD_LOGIC;
  SIGNAL nor_955_nl : STD_LOGIC;
  SIGNAL nor_956_nl : STD_LOGIC;
  SIGNAL mux_436_nl : STD_LOGIC;
  SIGNAL mux_435_nl : STD_LOGIC;
  SIGNAL mux_434_nl : STD_LOGIC;
  SIGNAL or_431_nl : STD_LOGIC;
  SIGNAL or_429_nl : STD_LOGIC;
  SIGNAL mux_433_nl : STD_LOGIC;
  SIGNAL or_428_nl : STD_LOGIC;
  SIGNAL or_426_nl : STD_LOGIC;
  SIGNAL mux_432_nl : STD_LOGIC;
  SIGNAL mux_431_nl : STD_LOGIC;
  SIGNAL or_425_nl : STD_LOGIC;
  SIGNAL or_423_nl : STD_LOGIC;
  SIGNAL mux_430_nl : STD_LOGIC;
  SIGNAL or_422_nl : STD_LOGIC;
  SIGNAL or_420_nl : STD_LOGIC;
  SIGNAL mux_460_nl : STD_LOGIC;
  SIGNAL nand_502_nl : STD_LOGIC;
  SIGNAL mux_459_nl : STD_LOGIC;
  SIGNAL and_431_nl : STD_LOGIC;
  SIGNAL mux_458_nl : STD_LOGIC;
  SIGNAL mux_457_nl : STD_LOGIC;
  SIGNAL nor_942_nl : STD_LOGIC;
  SIGNAL nor_943_nl : STD_LOGIC;
  SIGNAL mux_456_nl : STD_LOGIC;
  SIGNAL nor_944_nl : STD_LOGIC;
  SIGNAL nor_945_nl : STD_LOGIC;
  SIGNAL nor_946_nl : STD_LOGIC;
  SIGNAL mux_455_nl : STD_LOGIC;
  SIGNAL mux_454_nl : STD_LOGIC;
  SIGNAL or_465_nl : STD_LOGIC;
  SIGNAL or_463_nl : STD_LOGIC;
  SIGNAL mux_453_nl : STD_LOGIC;
  SIGNAL or_462_nl : STD_LOGIC;
  SIGNAL or_460_nl : STD_LOGIC;
  SIGNAL or_2276_nl : STD_LOGIC;
  SIGNAL mux_452_nl : STD_LOGIC;
  SIGNAL nand_30_nl : STD_LOGIC;
  SIGNAL mux_451_nl : STD_LOGIC;
  SIGNAL mux_450_nl : STD_LOGIC;
  SIGNAL nor_948_nl : STD_LOGIC;
  SIGNAL nor_949_nl : STD_LOGIC;
  SIGNAL nor_950_nl : STD_LOGIC;
  SIGNAL mux_449_nl : STD_LOGIC;
  SIGNAL or_454_nl : STD_LOGIC;
  SIGNAL or_452_nl : STD_LOGIC;
  SIGNAL or_451_nl : STD_LOGIC;
  SIGNAL mux_448_nl : STD_LOGIC;
  SIGNAL mux_447_nl : STD_LOGIC;
  SIGNAL or_450_nl : STD_LOGIC;
  SIGNAL or_448_nl : STD_LOGIC;
  SIGNAL or_447_nl : STD_LOGIC;
  SIGNAL mux_476_nl : STD_LOGIC;
  SIGNAL mux_475_nl : STD_LOGIC;
  SIGNAL mux_474_nl : STD_LOGIC;
  SIGNAL nor_935_nl : STD_LOGIC;
  SIGNAL nor_936_nl : STD_LOGIC;
  SIGNAL mux_473_nl : STD_LOGIC;
  SIGNAL nor_937_nl : STD_LOGIC;
  SIGNAL mux_469_nl : STD_LOGIC;
  SIGNAL nor_938_nl : STD_LOGIC;
  SIGNAL mux_468_nl : STD_LOGIC;
  SIGNAL nor_939_nl : STD_LOGIC;
  SIGNAL nor_940_nl : STD_LOGIC;
  SIGNAL nor_941_nl : STD_LOGIC;
  SIGNAL mux_467_nl : STD_LOGIC;
  SIGNAL mux_466_nl : STD_LOGIC;
  SIGNAL mux_465_nl : STD_LOGIC;
  SIGNAL or_484_nl : STD_LOGIC;
  SIGNAL or_482_nl : STD_LOGIC;
  SIGNAL mux_464_nl : STD_LOGIC;
  SIGNAL or_481_nl : STD_LOGIC;
  SIGNAL or_479_nl : STD_LOGIC;
  SIGNAL mux_463_nl : STD_LOGIC;
  SIGNAL mux_462_nl : STD_LOGIC;
  SIGNAL or_478_nl : STD_LOGIC;
  SIGNAL or_476_nl : STD_LOGIC;
  SIGNAL mux_461_nl : STD_LOGIC;
  SIGNAL or_475_nl : STD_LOGIC;
  SIGNAL or_473_nl : STD_LOGIC;
  SIGNAL mux_491_nl : STD_LOGIC;
  SIGNAL nand_501_nl : STD_LOGIC;
  SIGNAL mux_490_nl : STD_LOGIC;
  SIGNAL and_428_nl : STD_LOGIC;
  SIGNAL mux_489_nl : STD_LOGIC;
  SIGNAL mux_488_nl : STD_LOGIC;
  SIGNAL nor_923_nl : STD_LOGIC;
  SIGNAL nor_924_nl : STD_LOGIC;
  SIGNAL mux_487_nl : STD_LOGIC;
  SIGNAL nor_925_nl : STD_LOGIC;
  SIGNAL nor_926_nl : STD_LOGIC;
  SIGNAL nor_927_nl : STD_LOGIC;
  SIGNAL mux_486_nl : STD_LOGIC;
  SIGNAL mux_485_nl : STD_LOGIC;
  SIGNAL or_516_nl : STD_LOGIC;
  SIGNAL or_514_nl : STD_LOGIC;
  SIGNAL mux_484_nl : STD_LOGIC;
  SIGNAL or_513_nl : STD_LOGIC;
  SIGNAL or_511_nl : STD_LOGIC;
  SIGNAL or_2275_nl : STD_LOGIC;
  SIGNAL mux_483_nl : STD_LOGIC;
  SIGNAL nand_36_nl : STD_LOGIC;
  SIGNAL mux_482_nl : STD_LOGIC;
  SIGNAL mux_481_nl : STD_LOGIC;
  SIGNAL nor_929_nl : STD_LOGIC;
  SIGNAL nor_930_nl : STD_LOGIC;
  SIGNAL and_429_nl : STD_LOGIC;
  SIGNAL mux_480_nl : STD_LOGIC;
  SIGNAL nor_931_nl : STD_LOGIC;
  SIGNAL nor_932_nl : STD_LOGIC;
  SIGNAL or_503_nl : STD_LOGIC;
  SIGNAL mux_479_nl : STD_LOGIC;
  SIGNAL mux_478_nl : STD_LOGIC;
  SIGNAL or_502_nl : STD_LOGIC;
  SIGNAL or_500_nl : STD_LOGIC;
  SIGNAL nand_34_nl : STD_LOGIC;
  SIGNAL mux_507_nl : STD_LOGIC;
  SIGNAL mux_506_nl : STD_LOGIC;
  SIGNAL mux_505_nl : STD_LOGIC;
  SIGNAL nor_917_nl : STD_LOGIC;
  SIGNAL nor_918_nl : STD_LOGIC;
  SIGNAL mux_504_nl : STD_LOGIC;
  SIGNAL and_426_nl : STD_LOGIC;
  SIGNAL mux_500_nl : STD_LOGIC;
  SIGNAL nor_919_nl : STD_LOGIC;
  SIGNAL mux_499_nl : STD_LOGIC;
  SIGNAL nor_920_nl : STD_LOGIC;
  SIGNAL nor_921_nl : STD_LOGIC;
  SIGNAL nor_922_nl : STD_LOGIC;
  SIGNAL mux_498_nl : STD_LOGIC;
  SIGNAL mux_497_nl : STD_LOGIC;
  SIGNAL mux_496_nl : STD_LOGIC;
  SIGNAL or_535_nl : STD_LOGIC;
  SIGNAL or_533_nl : STD_LOGIC;
  SIGNAL mux_495_nl : STD_LOGIC;
  SIGNAL or_532_nl : STD_LOGIC;
  SIGNAL or_530_nl : STD_LOGIC;
  SIGNAL mux_494_nl : STD_LOGIC;
  SIGNAL mux_493_nl : STD_LOGIC;
  SIGNAL or_529_nl : STD_LOGIC;
  SIGNAL or_527_nl : STD_LOGIC;
  SIGNAL mux_492_nl : STD_LOGIC;
  SIGNAL or_526_nl : STD_LOGIC;
  SIGNAL or_524_nl : STD_LOGIC;
  SIGNAL mux_522_nl : STD_LOGIC;
  SIGNAL nand_500_nl : STD_LOGIC;
  SIGNAL mux_521_nl : STD_LOGIC;
  SIGNAL and_425_nl : STD_LOGIC;
  SIGNAL mux_520_nl : STD_LOGIC;
  SIGNAL mux_519_nl : STD_LOGIC;
  SIGNAL nor_908_nl : STD_LOGIC;
  SIGNAL nor_909_nl : STD_LOGIC;
  SIGNAL mux_518_nl : STD_LOGIC;
  SIGNAL nor_910_nl : STD_LOGIC;
  SIGNAL nor_911_nl : STD_LOGIC;
  SIGNAL nor_912_nl : STD_LOGIC;
  SIGNAL mux_517_nl : STD_LOGIC;
  SIGNAL mux_516_nl : STD_LOGIC;
  SIGNAL or_569_nl : STD_LOGIC;
  SIGNAL or_567_nl : STD_LOGIC;
  SIGNAL mux_515_nl : STD_LOGIC;
  SIGNAL or_566_nl : STD_LOGIC;
  SIGNAL or_564_nl : STD_LOGIC;
  SIGNAL or_2274_nl : STD_LOGIC;
  SIGNAL mux_514_nl : STD_LOGIC;
  SIGNAL nand_41_nl : STD_LOGIC;
  SIGNAL mux_513_nl : STD_LOGIC;
  SIGNAL mux_512_nl : STD_LOGIC;
  SIGNAL nor_914_nl : STD_LOGIC;
  SIGNAL nor_915_nl : STD_LOGIC;
  SIGNAL nor_916_nl : STD_LOGIC;
  SIGNAL mux_511_nl : STD_LOGIC;
  SIGNAL or_558_nl : STD_LOGIC;
  SIGNAL or_556_nl : STD_LOGIC;
  SIGNAL or_555_nl : STD_LOGIC;
  SIGNAL mux_510_nl : STD_LOGIC;
  SIGNAL mux_509_nl : STD_LOGIC;
  SIGNAL or_554_nl : STD_LOGIC;
  SIGNAL or_552_nl : STD_LOGIC;
  SIGNAL or_551_nl : STD_LOGIC;
  SIGNAL mux_538_nl : STD_LOGIC;
  SIGNAL mux_537_nl : STD_LOGIC;
  SIGNAL mux_536_nl : STD_LOGIC;
  SIGNAL nor_901_nl : STD_LOGIC;
  SIGNAL nor_902_nl : STD_LOGIC;
  SIGNAL mux_535_nl : STD_LOGIC;
  SIGNAL nor_903_nl : STD_LOGIC;
  SIGNAL mux_531_nl : STD_LOGIC;
  SIGNAL nor_904_nl : STD_LOGIC;
  SIGNAL mux_530_nl : STD_LOGIC;
  SIGNAL nor_905_nl : STD_LOGIC;
  SIGNAL nor_906_nl : STD_LOGIC;
  SIGNAL nor_907_nl : STD_LOGIC;
  SIGNAL mux_529_nl : STD_LOGIC;
  SIGNAL mux_528_nl : STD_LOGIC;
  SIGNAL mux_527_nl : STD_LOGIC;
  SIGNAL or_588_nl : STD_LOGIC;
  SIGNAL or_586_nl : STD_LOGIC;
  SIGNAL mux_526_nl : STD_LOGIC;
  SIGNAL or_585_nl : STD_LOGIC;
  SIGNAL or_583_nl : STD_LOGIC;
  SIGNAL mux_525_nl : STD_LOGIC;
  SIGNAL mux_524_nl : STD_LOGIC;
  SIGNAL or_582_nl : STD_LOGIC;
  SIGNAL or_580_nl : STD_LOGIC;
  SIGNAL mux_523_nl : STD_LOGIC;
  SIGNAL or_579_nl : STD_LOGIC;
  SIGNAL or_577_nl : STD_LOGIC;
  SIGNAL mux_553_nl : STD_LOGIC;
  SIGNAL nand_499_nl : STD_LOGIC;
  SIGNAL mux_552_nl : STD_LOGIC;
  SIGNAL and_422_nl : STD_LOGIC;
  SIGNAL mux_551_nl : STD_LOGIC;
  SIGNAL mux_550_nl : STD_LOGIC;
  SIGNAL nor_889_nl : STD_LOGIC;
  SIGNAL nor_890_nl : STD_LOGIC;
  SIGNAL mux_549_nl : STD_LOGIC;
  SIGNAL nor_891_nl : STD_LOGIC;
  SIGNAL nor_892_nl : STD_LOGIC;
  SIGNAL nor_893_nl : STD_LOGIC;
  SIGNAL mux_548_nl : STD_LOGIC;
  SIGNAL mux_547_nl : STD_LOGIC;
  SIGNAL or_620_nl : STD_LOGIC;
  SIGNAL or_618_nl : STD_LOGIC;
  SIGNAL mux_546_nl : STD_LOGIC;
  SIGNAL or_617_nl : STD_LOGIC;
  SIGNAL or_615_nl : STD_LOGIC;
  SIGNAL or_2273_nl : STD_LOGIC;
  SIGNAL mux_545_nl : STD_LOGIC;
  SIGNAL nand_47_nl : STD_LOGIC;
  SIGNAL mux_544_nl : STD_LOGIC;
  SIGNAL mux_543_nl : STD_LOGIC;
  SIGNAL nor_895_nl : STD_LOGIC;
  SIGNAL nor_896_nl : STD_LOGIC;
  SIGNAL and_423_nl : STD_LOGIC;
  SIGNAL mux_542_nl : STD_LOGIC;
  SIGNAL nor_897_nl : STD_LOGIC;
  SIGNAL nor_898_nl : STD_LOGIC;
  SIGNAL or_607_nl : STD_LOGIC;
  SIGNAL mux_541_nl : STD_LOGIC;
  SIGNAL mux_540_nl : STD_LOGIC;
  SIGNAL or_606_nl : STD_LOGIC;
  SIGNAL or_604_nl : STD_LOGIC;
  SIGNAL nand_45_nl : STD_LOGIC;
  SIGNAL mux_569_nl : STD_LOGIC;
  SIGNAL mux_568_nl : STD_LOGIC;
  SIGNAL mux_567_nl : STD_LOGIC;
  SIGNAL nor_883_nl : STD_LOGIC;
  SIGNAL nor_884_nl : STD_LOGIC;
  SIGNAL mux_566_nl : STD_LOGIC;
  SIGNAL and_420_nl : STD_LOGIC;
  SIGNAL mux_562_nl : STD_LOGIC;
  SIGNAL nor_885_nl : STD_LOGIC;
  SIGNAL mux_561_nl : STD_LOGIC;
  SIGNAL nor_886_nl : STD_LOGIC;
  SIGNAL nor_887_nl : STD_LOGIC;
  SIGNAL nor_888_nl : STD_LOGIC;
  SIGNAL mux_560_nl : STD_LOGIC;
  SIGNAL mux_559_nl : STD_LOGIC;
  SIGNAL mux_558_nl : STD_LOGIC;
  SIGNAL or_639_nl : STD_LOGIC;
  SIGNAL or_637_nl : STD_LOGIC;
  SIGNAL mux_557_nl : STD_LOGIC;
  SIGNAL or_636_nl : STD_LOGIC;
  SIGNAL or_634_nl : STD_LOGIC;
  SIGNAL mux_556_nl : STD_LOGIC;
  SIGNAL mux_555_nl : STD_LOGIC;
  SIGNAL or_633_nl : STD_LOGIC;
  SIGNAL or_631_nl : STD_LOGIC;
  SIGNAL mux_554_nl : STD_LOGIC;
  SIGNAL or_630_nl : STD_LOGIC;
  SIGNAL or_628_nl : STD_LOGIC;
  SIGNAL mux_584_nl : STD_LOGIC;
  SIGNAL nand_498_nl : STD_LOGIC;
  SIGNAL mux_583_nl : STD_LOGIC;
  SIGNAL and_419_nl : STD_LOGIC;
  SIGNAL mux_582_nl : STD_LOGIC;
  SIGNAL mux_581_nl : STD_LOGIC;
  SIGNAL nor_874_nl : STD_LOGIC;
  SIGNAL nor_875_nl : STD_LOGIC;
  SIGNAL mux_580_nl : STD_LOGIC;
  SIGNAL nor_876_nl : STD_LOGIC;
  SIGNAL nor_877_nl : STD_LOGIC;
  SIGNAL nor_878_nl : STD_LOGIC;
  SIGNAL mux_579_nl : STD_LOGIC;
  SIGNAL mux_578_nl : STD_LOGIC;
  SIGNAL or_673_nl : STD_LOGIC;
  SIGNAL or_671_nl : STD_LOGIC;
  SIGNAL mux_577_nl : STD_LOGIC;
  SIGNAL or_670_nl : STD_LOGIC;
  SIGNAL or_668_nl : STD_LOGIC;
  SIGNAL or_2272_nl : STD_LOGIC;
  SIGNAL mux_576_nl : STD_LOGIC;
  SIGNAL nand_52_nl : STD_LOGIC;
  SIGNAL mux_575_nl : STD_LOGIC;
  SIGNAL mux_574_nl : STD_LOGIC;
  SIGNAL nor_880_nl : STD_LOGIC;
  SIGNAL nor_881_nl : STD_LOGIC;
  SIGNAL nor_882_nl : STD_LOGIC;
  SIGNAL mux_573_nl : STD_LOGIC;
  SIGNAL or_662_nl : STD_LOGIC;
  SIGNAL or_660_nl : STD_LOGIC;
  SIGNAL or_659_nl : STD_LOGIC;
  SIGNAL mux_572_nl : STD_LOGIC;
  SIGNAL mux_571_nl : STD_LOGIC;
  SIGNAL or_658_nl : STD_LOGIC;
  SIGNAL or_656_nl : STD_LOGIC;
  SIGNAL or_655_nl : STD_LOGIC;
  SIGNAL mux_600_nl : STD_LOGIC;
  SIGNAL mux_599_nl : STD_LOGIC;
  SIGNAL mux_598_nl : STD_LOGIC;
  SIGNAL nor_867_nl : STD_LOGIC;
  SIGNAL nor_868_nl : STD_LOGIC;
  SIGNAL mux_597_nl : STD_LOGIC;
  SIGNAL nor_869_nl : STD_LOGIC;
  SIGNAL mux_593_nl : STD_LOGIC;
  SIGNAL nor_870_nl : STD_LOGIC;
  SIGNAL mux_592_nl : STD_LOGIC;
  SIGNAL nor_871_nl : STD_LOGIC;
  SIGNAL nor_872_nl : STD_LOGIC;
  SIGNAL nor_873_nl : STD_LOGIC;
  SIGNAL mux_591_nl : STD_LOGIC;
  SIGNAL mux_590_nl : STD_LOGIC;
  SIGNAL mux_589_nl : STD_LOGIC;
  SIGNAL or_692_nl : STD_LOGIC;
  SIGNAL or_690_nl : STD_LOGIC;
  SIGNAL mux_588_nl : STD_LOGIC;
  SIGNAL or_689_nl : STD_LOGIC;
  SIGNAL or_687_nl : STD_LOGIC;
  SIGNAL mux_587_nl : STD_LOGIC;
  SIGNAL mux_586_nl : STD_LOGIC;
  SIGNAL or_686_nl : STD_LOGIC;
  SIGNAL or_684_nl : STD_LOGIC;
  SIGNAL mux_585_nl : STD_LOGIC;
  SIGNAL or_683_nl : STD_LOGIC;
  SIGNAL or_681_nl : STD_LOGIC;
  SIGNAL mux_615_nl : STD_LOGIC;
  SIGNAL nand_497_nl : STD_LOGIC;
  SIGNAL mux_614_nl : STD_LOGIC;
  SIGNAL and_416_nl : STD_LOGIC;
  SIGNAL mux_613_nl : STD_LOGIC;
  SIGNAL mux_612_nl : STD_LOGIC;
  SIGNAL nor_855_nl : STD_LOGIC;
  SIGNAL nor_856_nl : STD_LOGIC;
  SIGNAL mux_611_nl : STD_LOGIC;
  SIGNAL nor_857_nl : STD_LOGIC;
  SIGNAL nor_858_nl : STD_LOGIC;
  SIGNAL nor_859_nl : STD_LOGIC;
  SIGNAL mux_610_nl : STD_LOGIC;
  SIGNAL mux_609_nl : STD_LOGIC;
  SIGNAL or_724_nl : STD_LOGIC;
  SIGNAL or_722_nl : STD_LOGIC;
  SIGNAL mux_608_nl : STD_LOGIC;
  SIGNAL or_721_nl : STD_LOGIC;
  SIGNAL or_719_nl : STD_LOGIC;
  SIGNAL or_2271_nl : STD_LOGIC;
  SIGNAL mux_607_nl : STD_LOGIC;
  SIGNAL nand_58_nl : STD_LOGIC;
  SIGNAL mux_606_nl : STD_LOGIC;
  SIGNAL mux_605_nl : STD_LOGIC;
  SIGNAL nor_861_nl : STD_LOGIC;
  SIGNAL nor_862_nl : STD_LOGIC;
  SIGNAL and_417_nl : STD_LOGIC;
  SIGNAL mux_604_nl : STD_LOGIC;
  SIGNAL nor_863_nl : STD_LOGIC;
  SIGNAL nor_864_nl : STD_LOGIC;
  SIGNAL or_711_nl : STD_LOGIC;
  SIGNAL mux_603_nl : STD_LOGIC;
  SIGNAL mux_602_nl : STD_LOGIC;
  SIGNAL or_710_nl : STD_LOGIC;
  SIGNAL or_708_nl : STD_LOGIC;
  SIGNAL nand_56_nl : STD_LOGIC;
  SIGNAL mux_631_nl : STD_LOGIC;
  SIGNAL mux_630_nl : STD_LOGIC;
  SIGNAL mux_629_nl : STD_LOGIC;
  SIGNAL nor_849_nl : STD_LOGIC;
  SIGNAL nor_850_nl : STD_LOGIC;
  SIGNAL mux_628_nl : STD_LOGIC;
  SIGNAL and_414_nl : STD_LOGIC;
  SIGNAL mux_624_nl : STD_LOGIC;
  SIGNAL nor_851_nl : STD_LOGIC;
  SIGNAL mux_623_nl : STD_LOGIC;
  SIGNAL nor_852_nl : STD_LOGIC;
  SIGNAL nor_853_nl : STD_LOGIC;
  SIGNAL nor_854_nl : STD_LOGIC;
  SIGNAL mux_622_nl : STD_LOGIC;
  SIGNAL mux_621_nl : STD_LOGIC;
  SIGNAL mux_620_nl : STD_LOGIC;
  SIGNAL or_743_nl : STD_LOGIC;
  SIGNAL or_741_nl : STD_LOGIC;
  SIGNAL mux_619_nl : STD_LOGIC;
  SIGNAL or_740_nl : STD_LOGIC;
  SIGNAL or_738_nl : STD_LOGIC;
  SIGNAL mux_618_nl : STD_LOGIC;
  SIGNAL mux_617_nl : STD_LOGIC;
  SIGNAL or_737_nl : STD_LOGIC;
  SIGNAL or_735_nl : STD_LOGIC;
  SIGNAL mux_616_nl : STD_LOGIC;
  SIGNAL or_734_nl : STD_LOGIC;
  SIGNAL or_732_nl : STD_LOGIC;
  SIGNAL mux_646_nl : STD_LOGIC;
  SIGNAL nand_496_nl : STD_LOGIC;
  SIGNAL mux_645_nl : STD_LOGIC;
  SIGNAL and_413_nl : STD_LOGIC;
  SIGNAL mux_644_nl : STD_LOGIC;
  SIGNAL mux_643_nl : STD_LOGIC;
  SIGNAL nor_840_nl : STD_LOGIC;
  SIGNAL nor_841_nl : STD_LOGIC;
  SIGNAL mux_642_nl : STD_LOGIC;
  SIGNAL nor_842_nl : STD_LOGIC;
  SIGNAL nor_843_nl : STD_LOGIC;
  SIGNAL nor_844_nl : STD_LOGIC;
  SIGNAL mux_641_nl : STD_LOGIC;
  SIGNAL mux_640_nl : STD_LOGIC;
  SIGNAL or_777_nl : STD_LOGIC;
  SIGNAL or_775_nl : STD_LOGIC;
  SIGNAL mux_639_nl : STD_LOGIC;
  SIGNAL or_774_nl : STD_LOGIC;
  SIGNAL or_772_nl : STD_LOGIC;
  SIGNAL or_2270_nl : STD_LOGIC;
  SIGNAL mux_638_nl : STD_LOGIC;
  SIGNAL nand_63_nl : STD_LOGIC;
  SIGNAL mux_637_nl : STD_LOGIC;
  SIGNAL mux_636_nl : STD_LOGIC;
  SIGNAL nor_846_nl : STD_LOGIC;
  SIGNAL nor_847_nl : STD_LOGIC;
  SIGNAL nor_848_nl : STD_LOGIC;
  SIGNAL mux_635_nl : STD_LOGIC;
  SIGNAL or_766_nl : STD_LOGIC;
  SIGNAL or_764_nl : STD_LOGIC;
  SIGNAL or_763_nl : STD_LOGIC;
  SIGNAL mux_634_nl : STD_LOGIC;
  SIGNAL mux_633_nl : STD_LOGIC;
  SIGNAL or_762_nl : STD_LOGIC;
  SIGNAL or_760_nl : STD_LOGIC;
  SIGNAL or_759_nl : STD_LOGIC;
  SIGNAL mux_662_nl : STD_LOGIC;
  SIGNAL mux_661_nl : STD_LOGIC;
  SIGNAL mux_660_nl : STD_LOGIC;
  SIGNAL nor_833_nl : STD_LOGIC;
  SIGNAL nor_834_nl : STD_LOGIC;
  SIGNAL mux_659_nl : STD_LOGIC;
  SIGNAL nor_835_nl : STD_LOGIC;
  SIGNAL mux_655_nl : STD_LOGIC;
  SIGNAL nor_836_nl : STD_LOGIC;
  SIGNAL mux_654_nl : STD_LOGIC;
  SIGNAL nor_837_nl : STD_LOGIC;
  SIGNAL nor_838_nl : STD_LOGIC;
  SIGNAL nor_839_nl : STD_LOGIC;
  SIGNAL mux_653_nl : STD_LOGIC;
  SIGNAL mux_652_nl : STD_LOGIC;
  SIGNAL mux_651_nl : STD_LOGIC;
  SIGNAL or_796_nl : STD_LOGIC;
  SIGNAL or_794_nl : STD_LOGIC;
  SIGNAL mux_650_nl : STD_LOGIC;
  SIGNAL or_793_nl : STD_LOGIC;
  SIGNAL or_791_nl : STD_LOGIC;
  SIGNAL mux_649_nl : STD_LOGIC;
  SIGNAL mux_648_nl : STD_LOGIC;
  SIGNAL or_790_nl : STD_LOGIC;
  SIGNAL or_788_nl : STD_LOGIC;
  SIGNAL mux_647_nl : STD_LOGIC;
  SIGNAL or_787_nl : STD_LOGIC;
  SIGNAL or_785_nl : STD_LOGIC;
  SIGNAL mux_677_nl : STD_LOGIC;
  SIGNAL nand_495_nl : STD_LOGIC;
  SIGNAL mux_676_nl : STD_LOGIC;
  SIGNAL and_410_nl : STD_LOGIC;
  SIGNAL mux_675_nl : STD_LOGIC;
  SIGNAL mux_674_nl : STD_LOGIC;
  SIGNAL nor_821_nl : STD_LOGIC;
  SIGNAL nor_822_nl : STD_LOGIC;
  SIGNAL mux_673_nl : STD_LOGIC;
  SIGNAL nor_823_nl : STD_LOGIC;
  SIGNAL nor_824_nl : STD_LOGIC;
  SIGNAL nor_825_nl : STD_LOGIC;
  SIGNAL mux_672_nl : STD_LOGIC;
  SIGNAL mux_671_nl : STD_LOGIC;
  SIGNAL or_828_nl : STD_LOGIC;
  SIGNAL or_826_nl : STD_LOGIC;
  SIGNAL mux_670_nl : STD_LOGIC;
  SIGNAL or_825_nl : STD_LOGIC;
  SIGNAL or_823_nl : STD_LOGIC;
  SIGNAL or_2269_nl : STD_LOGIC;
  SIGNAL mux_669_nl : STD_LOGIC;
  SIGNAL nand_69_nl : STD_LOGIC;
  SIGNAL mux_668_nl : STD_LOGIC;
  SIGNAL mux_667_nl : STD_LOGIC;
  SIGNAL nor_827_nl : STD_LOGIC;
  SIGNAL nor_828_nl : STD_LOGIC;
  SIGNAL and_411_nl : STD_LOGIC;
  SIGNAL mux_666_nl : STD_LOGIC;
  SIGNAL nor_829_nl : STD_LOGIC;
  SIGNAL nor_830_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL mux_665_nl : STD_LOGIC;
  SIGNAL mux_664_nl : STD_LOGIC;
  SIGNAL or_814_nl : STD_LOGIC;
  SIGNAL or_812_nl : STD_LOGIC;
  SIGNAL nand_67_nl : STD_LOGIC;
  SIGNAL mux_693_nl : STD_LOGIC;
  SIGNAL mux_692_nl : STD_LOGIC;
  SIGNAL mux_691_nl : STD_LOGIC;
  SIGNAL nor_815_nl : STD_LOGIC;
  SIGNAL nor_816_nl : STD_LOGIC;
  SIGNAL mux_690_nl : STD_LOGIC;
  SIGNAL and_408_nl : STD_LOGIC;
  SIGNAL mux_686_nl : STD_LOGIC;
  SIGNAL nor_817_nl : STD_LOGIC;
  SIGNAL mux_685_nl : STD_LOGIC;
  SIGNAL nor_818_nl : STD_LOGIC;
  SIGNAL nor_819_nl : STD_LOGIC;
  SIGNAL nor_820_nl : STD_LOGIC;
  SIGNAL mux_684_nl : STD_LOGIC;
  SIGNAL mux_683_nl : STD_LOGIC;
  SIGNAL mux_682_nl : STD_LOGIC;
  SIGNAL or_847_nl : STD_LOGIC;
  SIGNAL or_845_nl : STD_LOGIC;
  SIGNAL mux_681_nl : STD_LOGIC;
  SIGNAL or_844_nl : STD_LOGIC;
  SIGNAL or_842_nl : STD_LOGIC;
  SIGNAL mux_680_nl : STD_LOGIC;
  SIGNAL mux_679_nl : STD_LOGIC;
  SIGNAL or_841_nl : STD_LOGIC;
  SIGNAL or_839_nl : STD_LOGIC;
  SIGNAL mux_678_nl : STD_LOGIC;
  SIGNAL or_838_nl : STD_LOGIC;
  SIGNAL or_836_nl : STD_LOGIC;
  SIGNAL mux_708_nl : STD_LOGIC;
  SIGNAL nand_494_nl : STD_LOGIC;
  SIGNAL mux_707_nl : STD_LOGIC;
  SIGNAL and_407_nl : STD_LOGIC;
  SIGNAL mux_706_nl : STD_LOGIC;
  SIGNAL mux_705_nl : STD_LOGIC;
  SIGNAL nor_806_nl : STD_LOGIC;
  SIGNAL nor_807_nl : STD_LOGIC;
  SIGNAL mux_704_nl : STD_LOGIC;
  SIGNAL nor_808_nl : STD_LOGIC;
  SIGNAL nor_809_nl : STD_LOGIC;
  SIGNAL nor_810_nl : STD_LOGIC;
  SIGNAL mux_703_nl : STD_LOGIC;
  SIGNAL mux_702_nl : STD_LOGIC;
  SIGNAL or_881_nl : STD_LOGIC;
  SIGNAL or_879_nl : STD_LOGIC;
  SIGNAL mux_701_nl : STD_LOGIC;
  SIGNAL or_878_nl : STD_LOGIC;
  SIGNAL or_876_nl : STD_LOGIC;
  SIGNAL or_2268_nl : STD_LOGIC;
  SIGNAL mux_700_nl : STD_LOGIC;
  SIGNAL nand_74_nl : STD_LOGIC;
  SIGNAL mux_699_nl : STD_LOGIC;
  SIGNAL mux_698_nl : STD_LOGIC;
  SIGNAL nor_812_nl : STD_LOGIC;
  SIGNAL nor_813_nl : STD_LOGIC;
  SIGNAL nor_814_nl : STD_LOGIC;
  SIGNAL mux_697_nl : STD_LOGIC;
  SIGNAL or_870_nl : STD_LOGIC;
  SIGNAL or_868_nl : STD_LOGIC;
  SIGNAL or_867_nl : STD_LOGIC;
  SIGNAL mux_696_nl : STD_LOGIC;
  SIGNAL mux_695_nl : STD_LOGIC;
  SIGNAL or_866_nl : STD_LOGIC;
  SIGNAL or_864_nl : STD_LOGIC;
  SIGNAL or_863_nl : STD_LOGIC;
  SIGNAL mux_724_nl : STD_LOGIC;
  SIGNAL mux_723_nl : STD_LOGIC;
  SIGNAL mux_722_nl : STD_LOGIC;
  SIGNAL nor_799_nl : STD_LOGIC;
  SIGNAL nor_800_nl : STD_LOGIC;
  SIGNAL mux_721_nl : STD_LOGIC;
  SIGNAL nor_801_nl : STD_LOGIC;
  SIGNAL mux_717_nl : STD_LOGIC;
  SIGNAL nor_802_nl : STD_LOGIC;
  SIGNAL mux_716_nl : STD_LOGIC;
  SIGNAL nor_803_nl : STD_LOGIC;
  SIGNAL nor_804_nl : STD_LOGIC;
  SIGNAL nor_805_nl : STD_LOGIC;
  SIGNAL mux_715_nl : STD_LOGIC;
  SIGNAL mux_714_nl : STD_LOGIC;
  SIGNAL mux_713_nl : STD_LOGIC;
  SIGNAL or_900_nl : STD_LOGIC;
  SIGNAL or_898_nl : STD_LOGIC;
  SIGNAL mux_712_nl : STD_LOGIC;
  SIGNAL or_897_nl : STD_LOGIC;
  SIGNAL or_895_nl : STD_LOGIC;
  SIGNAL mux_711_nl : STD_LOGIC;
  SIGNAL mux_710_nl : STD_LOGIC;
  SIGNAL or_894_nl : STD_LOGIC;
  SIGNAL or_892_nl : STD_LOGIC;
  SIGNAL mux_709_nl : STD_LOGIC;
  SIGNAL or_891_nl : STD_LOGIC;
  SIGNAL or_889_nl : STD_LOGIC;
  SIGNAL mux_739_nl : STD_LOGIC;
  SIGNAL nand_493_nl : STD_LOGIC;
  SIGNAL mux_738_nl : STD_LOGIC;
  SIGNAL and_404_nl : STD_LOGIC;
  SIGNAL mux_737_nl : STD_LOGIC;
  SIGNAL mux_736_nl : STD_LOGIC;
  SIGNAL nor_787_nl : STD_LOGIC;
  SIGNAL nor_788_nl : STD_LOGIC;
  SIGNAL mux_735_nl : STD_LOGIC;
  SIGNAL nor_789_nl : STD_LOGIC;
  SIGNAL nor_790_nl : STD_LOGIC;
  SIGNAL nor_791_nl : STD_LOGIC;
  SIGNAL mux_734_nl : STD_LOGIC;
  SIGNAL mux_733_nl : STD_LOGIC;
  SIGNAL or_932_nl : STD_LOGIC;
  SIGNAL or_930_nl : STD_LOGIC;
  SIGNAL mux_732_nl : STD_LOGIC;
  SIGNAL or_929_nl : STD_LOGIC;
  SIGNAL or_927_nl : STD_LOGIC;
  SIGNAL or_2267_nl : STD_LOGIC;
  SIGNAL mux_731_nl : STD_LOGIC;
  SIGNAL nand_80_nl : STD_LOGIC;
  SIGNAL mux_730_nl : STD_LOGIC;
  SIGNAL mux_729_nl : STD_LOGIC;
  SIGNAL nor_793_nl : STD_LOGIC;
  SIGNAL nor_794_nl : STD_LOGIC;
  SIGNAL and_405_nl : STD_LOGIC;
  SIGNAL mux_728_nl : STD_LOGIC;
  SIGNAL nor_795_nl : STD_LOGIC;
  SIGNAL nor_796_nl : STD_LOGIC;
  SIGNAL or_919_nl : STD_LOGIC;
  SIGNAL mux_727_nl : STD_LOGIC;
  SIGNAL mux_726_nl : STD_LOGIC;
  SIGNAL or_918_nl : STD_LOGIC;
  SIGNAL or_916_nl : STD_LOGIC;
  SIGNAL nand_78_nl : STD_LOGIC;
  SIGNAL mux_755_nl : STD_LOGIC;
  SIGNAL mux_754_nl : STD_LOGIC;
  SIGNAL mux_753_nl : STD_LOGIC;
  SIGNAL nor_781_nl : STD_LOGIC;
  SIGNAL nor_782_nl : STD_LOGIC;
  SIGNAL mux_752_nl : STD_LOGIC;
  SIGNAL and_402_nl : STD_LOGIC;
  SIGNAL mux_748_nl : STD_LOGIC;
  SIGNAL nor_783_nl : STD_LOGIC;
  SIGNAL mux_747_nl : STD_LOGIC;
  SIGNAL nor_784_nl : STD_LOGIC;
  SIGNAL nor_785_nl : STD_LOGIC;
  SIGNAL nor_786_nl : STD_LOGIC;
  SIGNAL mux_746_nl : STD_LOGIC;
  SIGNAL mux_745_nl : STD_LOGIC;
  SIGNAL mux_744_nl : STD_LOGIC;
  SIGNAL or_951_nl : STD_LOGIC;
  SIGNAL or_949_nl : STD_LOGIC;
  SIGNAL mux_743_nl : STD_LOGIC;
  SIGNAL or_948_nl : STD_LOGIC;
  SIGNAL or_946_nl : STD_LOGIC;
  SIGNAL mux_742_nl : STD_LOGIC;
  SIGNAL mux_741_nl : STD_LOGIC;
  SIGNAL or_945_nl : STD_LOGIC;
  SIGNAL or_943_nl : STD_LOGIC;
  SIGNAL mux_740_nl : STD_LOGIC;
  SIGNAL or_942_nl : STD_LOGIC;
  SIGNAL or_940_nl : STD_LOGIC;
  SIGNAL mux_770_nl : STD_LOGIC;
  SIGNAL nand_492_nl : STD_LOGIC;
  SIGNAL mux_769_nl : STD_LOGIC;
  SIGNAL and_401_nl : STD_LOGIC;
  SIGNAL mux_768_nl : STD_LOGIC;
  SIGNAL mux_767_nl : STD_LOGIC;
  SIGNAL nor_772_nl : STD_LOGIC;
  SIGNAL nor_773_nl : STD_LOGIC;
  SIGNAL mux_766_nl : STD_LOGIC;
  SIGNAL nor_774_nl : STD_LOGIC;
  SIGNAL nor_775_nl : STD_LOGIC;
  SIGNAL nor_776_nl : STD_LOGIC;
  SIGNAL mux_765_nl : STD_LOGIC;
  SIGNAL mux_764_nl : STD_LOGIC;
  SIGNAL or_984_nl : STD_LOGIC;
  SIGNAL or_982_nl : STD_LOGIC;
  SIGNAL mux_763_nl : STD_LOGIC;
  SIGNAL or_981_nl : STD_LOGIC;
  SIGNAL or_979_nl : STD_LOGIC;
  SIGNAL or_2266_nl : STD_LOGIC;
  SIGNAL mux_762_nl : STD_LOGIC;
  SIGNAL nand_85_nl : STD_LOGIC;
  SIGNAL mux_761_nl : STD_LOGIC;
  SIGNAL mux_760_nl : STD_LOGIC;
  SIGNAL nor_778_nl : STD_LOGIC;
  SIGNAL nor_779_nl : STD_LOGIC;
  SIGNAL nor_780_nl : STD_LOGIC;
  SIGNAL mux_759_nl : STD_LOGIC;
  SIGNAL or_973_nl : STD_LOGIC;
  SIGNAL or_972_nl : STD_LOGIC;
  SIGNAL or_971_nl : STD_LOGIC;
  SIGNAL mux_758_nl : STD_LOGIC;
  SIGNAL mux_757_nl : STD_LOGIC;
  SIGNAL or_970_nl : STD_LOGIC;
  SIGNAL or_968_nl : STD_LOGIC;
  SIGNAL or_967_nl : STD_LOGIC;
  SIGNAL mux_786_nl : STD_LOGIC;
  SIGNAL mux_785_nl : STD_LOGIC;
  SIGNAL mux_784_nl : STD_LOGIC;
  SIGNAL nor_765_nl : STD_LOGIC;
  SIGNAL nor_766_nl : STD_LOGIC;
  SIGNAL mux_783_nl : STD_LOGIC;
  SIGNAL nor_767_nl : STD_LOGIC;
  SIGNAL mux_779_nl : STD_LOGIC;
  SIGNAL nor_768_nl : STD_LOGIC;
  SIGNAL mux_778_nl : STD_LOGIC;
  SIGNAL nor_769_nl : STD_LOGIC;
  SIGNAL nor_770_nl : STD_LOGIC;
  SIGNAL nor_771_nl : STD_LOGIC;
  SIGNAL mux_777_nl : STD_LOGIC;
  SIGNAL mux_776_nl : STD_LOGIC;
  SIGNAL mux_775_nl : STD_LOGIC;
  SIGNAL or_1003_nl : STD_LOGIC;
  SIGNAL or_1001_nl : STD_LOGIC;
  SIGNAL mux_774_nl : STD_LOGIC;
  SIGNAL or_1000_nl : STD_LOGIC;
  SIGNAL or_998_nl : STD_LOGIC;
  SIGNAL mux_773_nl : STD_LOGIC;
  SIGNAL mux_772_nl : STD_LOGIC;
  SIGNAL or_997_nl : STD_LOGIC;
  SIGNAL or_995_nl : STD_LOGIC;
  SIGNAL mux_771_nl : STD_LOGIC;
  SIGNAL or_994_nl : STD_LOGIC;
  SIGNAL or_992_nl : STD_LOGIC;
  SIGNAL mux_801_nl : STD_LOGIC;
  SIGNAL nand_491_nl : STD_LOGIC;
  SIGNAL mux_800_nl : STD_LOGIC;
  SIGNAL and_398_nl : STD_LOGIC;
  SIGNAL mux_799_nl : STD_LOGIC;
  SIGNAL mux_798_nl : STD_LOGIC;
  SIGNAL nor_753_nl : STD_LOGIC;
  SIGNAL nor_754_nl : STD_LOGIC;
  SIGNAL mux_797_nl : STD_LOGIC;
  SIGNAL nor_755_nl : STD_LOGIC;
  SIGNAL nor_756_nl : STD_LOGIC;
  SIGNAL nor_757_nl : STD_LOGIC;
  SIGNAL mux_796_nl : STD_LOGIC;
  SIGNAL mux_795_nl : STD_LOGIC;
  SIGNAL nand_516_nl : STD_LOGIC;
  SIGNAL or_1031_nl : STD_LOGIC;
  SIGNAL mux_794_nl : STD_LOGIC;
  SIGNAL or_1030_nl : STD_LOGIC;
  SIGNAL or_1028_nl : STD_LOGIC;
  SIGNAL or_2265_nl : STD_LOGIC;
  SIGNAL mux_793_nl : STD_LOGIC;
  SIGNAL nand_91_nl : STD_LOGIC;
  SIGNAL mux_792_nl : STD_LOGIC;
  SIGNAL mux_791_nl : STD_LOGIC;
  SIGNAL nor_759_nl : STD_LOGIC;
  SIGNAL nor_760_nl : STD_LOGIC;
  SIGNAL and_399_nl : STD_LOGIC;
  SIGNAL mux_790_nl : STD_LOGIC;
  SIGNAL nor_761_nl : STD_LOGIC;
  SIGNAL nor_762_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL mux_789_nl : STD_LOGIC;
  SIGNAL mux_788_nl : STD_LOGIC;
  SIGNAL or_1021_nl : STD_LOGIC;
  SIGNAL or_1019_nl : STD_LOGIC;
  SIGNAL nand_89_nl : STD_LOGIC;
  SIGNAL mux_817_nl : STD_LOGIC;
  SIGNAL mux_816_nl : STD_LOGIC;
  SIGNAL mux_815_nl : STD_LOGIC;
  SIGNAL nor_748_nl : STD_LOGIC;
  SIGNAL nor_749_nl : STD_LOGIC;
  SIGNAL mux_814_nl : STD_LOGIC;
  SIGNAL and_395_nl : STD_LOGIC;
  SIGNAL mux_810_nl : STD_LOGIC;
  SIGNAL and_396_nl : STD_LOGIC;
  SIGNAL mux_809_nl : STD_LOGIC;
  SIGNAL and_527_nl : STD_LOGIC;
  SIGNAL nor_751_nl : STD_LOGIC;
  SIGNAL nor_752_nl : STD_LOGIC;
  SIGNAL mux_808_nl : STD_LOGIC;
  SIGNAL mux_807_nl : STD_LOGIC;
  SIGNAL mux_806_nl : STD_LOGIC;
  SIGNAL or_1051_nl : STD_LOGIC;
  SIGNAL nand_369_nl : STD_LOGIC;
  SIGNAL mux_805_nl : STD_LOGIC;
  SIGNAL nand_515_nl : STD_LOGIC;
  SIGNAL or_1046_nl : STD_LOGIC;
  SIGNAL mux_804_nl : STD_LOGIC;
  SIGNAL mux_803_nl : STD_LOGIC;
  SIGNAL or_1045_nl : STD_LOGIC;
  SIGNAL nand_373_nl : STD_LOGIC;
  SIGNAL mux_802_nl : STD_LOGIC;
  SIGNAL nand_471_nl : STD_LOGIC;
  SIGNAL or_1040_nl : STD_LOGIC;
  SIGNAL mux_832_nl : STD_LOGIC;
  SIGNAL nand_490_nl : STD_LOGIC;
  SIGNAL mux_831_nl : STD_LOGIC;
  SIGNAL and_394_nl : STD_LOGIC;
  SIGNAL mux_830_nl : STD_LOGIC;
  SIGNAL mux_829_nl : STD_LOGIC;
  SIGNAL nor_739_nl : STD_LOGIC;
  SIGNAL nor_740_nl : STD_LOGIC;
  SIGNAL mux_828_nl : STD_LOGIC;
  SIGNAL nor_741_nl : STD_LOGIC;
  SIGNAL nor_742_nl : STD_LOGIC;
  SIGNAL nor_743_nl : STD_LOGIC;
  SIGNAL mux_827_nl : STD_LOGIC;
  SIGNAL mux_826_nl : STD_LOGIC;
  SIGNAL or_1085_nl : STD_LOGIC;
  SIGNAL or_1083_nl : STD_LOGIC;
  SIGNAL mux_825_nl : STD_LOGIC;
  SIGNAL or_1082_nl : STD_LOGIC;
  SIGNAL or_1080_nl : STD_LOGIC;
  SIGNAL or_2264_nl : STD_LOGIC;
  SIGNAL mux_824_nl : STD_LOGIC;
  SIGNAL nand_96_nl : STD_LOGIC;
  SIGNAL mux_823_nl : STD_LOGIC;
  SIGNAL mux_822_nl : STD_LOGIC;
  SIGNAL nor_745_nl : STD_LOGIC;
  SIGNAL nor_746_nl : STD_LOGIC;
  SIGNAL nor_747_nl : STD_LOGIC;
  SIGNAL mux_821_nl : STD_LOGIC;
  SIGNAL or_1074_nl : STD_LOGIC;
  SIGNAL or_1072_nl : STD_LOGIC;
  SIGNAL or_1071_nl : STD_LOGIC;
  SIGNAL mux_820_nl : STD_LOGIC;
  SIGNAL mux_819_nl : STD_LOGIC;
  SIGNAL or_1070_nl : STD_LOGIC;
  SIGNAL or_1068_nl : STD_LOGIC;
  SIGNAL or_1067_nl : STD_LOGIC;
  SIGNAL mux_848_nl : STD_LOGIC;
  SIGNAL mux_847_nl : STD_LOGIC;
  SIGNAL mux_846_nl : STD_LOGIC;
  SIGNAL nor_732_nl : STD_LOGIC;
  SIGNAL nor_733_nl : STD_LOGIC;
  SIGNAL mux_845_nl : STD_LOGIC;
  SIGNAL nor_734_nl : STD_LOGIC;
  SIGNAL mux_841_nl : STD_LOGIC;
  SIGNAL nor_735_nl : STD_LOGIC;
  SIGNAL mux_840_nl : STD_LOGIC;
  SIGNAL nor_736_nl : STD_LOGIC;
  SIGNAL nor_737_nl : STD_LOGIC;
  SIGNAL nor_738_nl : STD_LOGIC;
  SIGNAL mux_839_nl : STD_LOGIC;
  SIGNAL mux_838_nl : STD_LOGIC;
  SIGNAL mux_837_nl : STD_LOGIC;
  SIGNAL or_1104_nl : STD_LOGIC;
  SIGNAL or_1102_nl : STD_LOGIC;
  SIGNAL mux_836_nl : STD_LOGIC;
  SIGNAL or_1101_nl : STD_LOGIC;
  SIGNAL or_1099_nl : STD_LOGIC;
  SIGNAL mux_835_nl : STD_LOGIC;
  SIGNAL mux_834_nl : STD_LOGIC;
  SIGNAL or_1098_nl : STD_LOGIC;
  SIGNAL or_1096_nl : STD_LOGIC;
  SIGNAL mux_833_nl : STD_LOGIC;
  SIGNAL or_1095_nl : STD_LOGIC;
  SIGNAL or_1093_nl : STD_LOGIC;
  SIGNAL mux_863_nl : STD_LOGIC;
  SIGNAL nand_489_nl : STD_LOGIC;
  SIGNAL mux_862_nl : STD_LOGIC;
  SIGNAL and_391_nl : STD_LOGIC;
  SIGNAL mux_861_nl : STD_LOGIC;
  SIGNAL mux_860_nl : STD_LOGIC;
  SIGNAL nor_720_nl : STD_LOGIC;
  SIGNAL nor_721_nl : STD_LOGIC;
  SIGNAL mux_859_nl : STD_LOGIC;
  SIGNAL nor_722_nl : STD_LOGIC;
  SIGNAL nor_723_nl : STD_LOGIC;
  SIGNAL nor_724_nl : STD_LOGIC;
  SIGNAL mux_858_nl : STD_LOGIC;
  SIGNAL mux_857_nl : STD_LOGIC;
  SIGNAL or_1136_nl : STD_LOGIC;
  SIGNAL or_1134_nl : STD_LOGIC;
  SIGNAL mux_856_nl : STD_LOGIC;
  SIGNAL or_1133_nl : STD_LOGIC;
  SIGNAL or_1131_nl : STD_LOGIC;
  SIGNAL or_2263_nl : STD_LOGIC;
  SIGNAL mux_855_nl : STD_LOGIC;
  SIGNAL nand_102_nl : STD_LOGIC;
  SIGNAL mux_854_nl : STD_LOGIC;
  SIGNAL mux_853_nl : STD_LOGIC;
  SIGNAL nor_726_nl : STD_LOGIC;
  SIGNAL nor_727_nl : STD_LOGIC;
  SIGNAL and_392_nl : STD_LOGIC;
  SIGNAL mux_852_nl : STD_LOGIC;
  SIGNAL nor_728_nl : STD_LOGIC;
  SIGNAL nor_729_nl : STD_LOGIC;
  SIGNAL or_1123_nl : STD_LOGIC;
  SIGNAL mux_851_nl : STD_LOGIC;
  SIGNAL mux_850_nl : STD_LOGIC;
  SIGNAL or_1122_nl : STD_LOGIC;
  SIGNAL or_1120_nl : STD_LOGIC;
  SIGNAL nand_100_nl : STD_LOGIC;
  SIGNAL mux_879_nl : STD_LOGIC;
  SIGNAL mux_878_nl : STD_LOGIC;
  SIGNAL mux_877_nl : STD_LOGIC;
  SIGNAL nor_714_nl : STD_LOGIC;
  SIGNAL nor_715_nl : STD_LOGIC;
  SIGNAL mux_876_nl : STD_LOGIC;
  SIGNAL and_389_nl : STD_LOGIC;
  SIGNAL mux_872_nl : STD_LOGIC;
  SIGNAL nor_716_nl : STD_LOGIC;
  SIGNAL mux_871_nl : STD_LOGIC;
  SIGNAL nor_717_nl : STD_LOGIC;
  SIGNAL nor_718_nl : STD_LOGIC;
  SIGNAL nor_719_nl : STD_LOGIC;
  SIGNAL mux_870_nl : STD_LOGIC;
  SIGNAL mux_869_nl : STD_LOGIC;
  SIGNAL mux_868_nl : STD_LOGIC;
  SIGNAL or_1155_nl : STD_LOGIC;
  SIGNAL or_1153_nl : STD_LOGIC;
  SIGNAL mux_867_nl : STD_LOGIC;
  SIGNAL or_1152_nl : STD_LOGIC;
  SIGNAL or_1150_nl : STD_LOGIC;
  SIGNAL mux_866_nl : STD_LOGIC;
  SIGNAL mux_865_nl : STD_LOGIC;
  SIGNAL or_1149_nl : STD_LOGIC;
  SIGNAL or_1147_nl : STD_LOGIC;
  SIGNAL mux_864_nl : STD_LOGIC;
  SIGNAL or_1146_nl : STD_LOGIC;
  SIGNAL or_1144_nl : STD_LOGIC;
  SIGNAL mux_894_nl : STD_LOGIC;
  SIGNAL nand_488_nl : STD_LOGIC;
  SIGNAL mux_893_nl : STD_LOGIC;
  SIGNAL and_388_nl : STD_LOGIC;
  SIGNAL mux_892_nl : STD_LOGIC;
  SIGNAL mux_891_nl : STD_LOGIC;
  SIGNAL nor_705_nl : STD_LOGIC;
  SIGNAL nor_706_nl : STD_LOGIC;
  SIGNAL mux_890_nl : STD_LOGIC;
  SIGNAL nor_707_nl : STD_LOGIC;
  SIGNAL nor_708_nl : STD_LOGIC;
  SIGNAL nor_709_nl : STD_LOGIC;
  SIGNAL mux_889_nl : STD_LOGIC;
  SIGNAL mux_888_nl : STD_LOGIC;
  SIGNAL or_1189_nl : STD_LOGIC;
  SIGNAL or_1187_nl : STD_LOGIC;
  SIGNAL mux_887_nl : STD_LOGIC;
  SIGNAL or_1186_nl : STD_LOGIC;
  SIGNAL or_1184_nl : STD_LOGIC;
  SIGNAL or_2262_nl : STD_LOGIC;
  SIGNAL mux_886_nl : STD_LOGIC;
  SIGNAL nand_107_nl : STD_LOGIC;
  SIGNAL mux_885_nl : STD_LOGIC;
  SIGNAL mux_884_nl : STD_LOGIC;
  SIGNAL nor_711_nl : STD_LOGIC;
  SIGNAL nor_712_nl : STD_LOGIC;
  SIGNAL nor_713_nl : STD_LOGIC;
  SIGNAL mux_883_nl : STD_LOGIC;
  SIGNAL or_1178_nl : STD_LOGIC;
  SIGNAL or_1176_nl : STD_LOGIC;
  SIGNAL or_1175_nl : STD_LOGIC;
  SIGNAL mux_882_nl : STD_LOGIC;
  SIGNAL mux_881_nl : STD_LOGIC;
  SIGNAL or_1174_nl : STD_LOGIC;
  SIGNAL or_1172_nl : STD_LOGIC;
  SIGNAL or_1171_nl : STD_LOGIC;
  SIGNAL mux_910_nl : STD_LOGIC;
  SIGNAL mux_909_nl : STD_LOGIC;
  SIGNAL mux_908_nl : STD_LOGIC;
  SIGNAL nor_698_nl : STD_LOGIC;
  SIGNAL nor_699_nl : STD_LOGIC;
  SIGNAL mux_907_nl : STD_LOGIC;
  SIGNAL nor_700_nl : STD_LOGIC;
  SIGNAL mux_903_nl : STD_LOGIC;
  SIGNAL nor_701_nl : STD_LOGIC;
  SIGNAL mux_902_nl : STD_LOGIC;
  SIGNAL nor_702_nl : STD_LOGIC;
  SIGNAL nor_703_nl : STD_LOGIC;
  SIGNAL nor_704_nl : STD_LOGIC;
  SIGNAL mux_901_nl : STD_LOGIC;
  SIGNAL mux_900_nl : STD_LOGIC;
  SIGNAL mux_899_nl : STD_LOGIC;
  SIGNAL or_1208_nl : STD_LOGIC;
  SIGNAL or_1206_nl : STD_LOGIC;
  SIGNAL mux_898_nl : STD_LOGIC;
  SIGNAL or_1205_nl : STD_LOGIC;
  SIGNAL or_1203_nl : STD_LOGIC;
  SIGNAL mux_897_nl : STD_LOGIC;
  SIGNAL mux_896_nl : STD_LOGIC;
  SIGNAL or_1202_nl : STD_LOGIC;
  SIGNAL or_1200_nl : STD_LOGIC;
  SIGNAL mux_895_nl : STD_LOGIC;
  SIGNAL or_1199_nl : STD_LOGIC;
  SIGNAL or_1197_nl : STD_LOGIC;
  SIGNAL mux_925_nl : STD_LOGIC;
  SIGNAL nand_487_nl : STD_LOGIC;
  SIGNAL mux_924_nl : STD_LOGIC;
  SIGNAL and_385_nl : STD_LOGIC;
  SIGNAL mux_923_nl : STD_LOGIC;
  SIGNAL mux_922_nl : STD_LOGIC;
  SIGNAL nor_686_nl : STD_LOGIC;
  SIGNAL nor_687_nl : STD_LOGIC;
  SIGNAL mux_921_nl : STD_LOGIC;
  SIGNAL nor_688_nl : STD_LOGIC;
  SIGNAL nor_689_nl : STD_LOGIC;
  SIGNAL nor_690_nl : STD_LOGIC;
  SIGNAL mux_920_nl : STD_LOGIC;
  SIGNAL mux_919_nl : STD_LOGIC;
  SIGNAL or_1240_nl : STD_LOGIC;
  SIGNAL or_1238_nl : STD_LOGIC;
  SIGNAL mux_918_nl : STD_LOGIC;
  SIGNAL or_1237_nl : STD_LOGIC;
  SIGNAL or_1235_nl : STD_LOGIC;
  SIGNAL or_2261_nl : STD_LOGIC;
  SIGNAL mux_917_nl : STD_LOGIC;
  SIGNAL nand_113_nl : STD_LOGIC;
  SIGNAL mux_916_nl : STD_LOGIC;
  SIGNAL mux_915_nl : STD_LOGIC;
  SIGNAL nor_692_nl : STD_LOGIC;
  SIGNAL nor_693_nl : STD_LOGIC;
  SIGNAL and_386_nl : STD_LOGIC;
  SIGNAL mux_914_nl : STD_LOGIC;
  SIGNAL nor_694_nl : STD_LOGIC;
  SIGNAL nor_695_nl : STD_LOGIC;
  SIGNAL or_1227_nl : STD_LOGIC;
  SIGNAL mux_913_nl : STD_LOGIC;
  SIGNAL mux_912_nl : STD_LOGIC;
  SIGNAL or_1226_nl : STD_LOGIC;
  SIGNAL or_1224_nl : STD_LOGIC;
  SIGNAL nand_111_nl : STD_LOGIC;
  SIGNAL mux_941_nl : STD_LOGIC;
  SIGNAL mux_940_nl : STD_LOGIC;
  SIGNAL mux_939_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL mux_938_nl : STD_LOGIC;
  SIGNAL and_383_nl : STD_LOGIC;
  SIGNAL mux_934_nl : STD_LOGIC;
  SIGNAL nor_682_nl : STD_LOGIC;
  SIGNAL mux_933_nl : STD_LOGIC;
  SIGNAL nor_683_nl : STD_LOGIC;
  SIGNAL nor_684_nl : STD_LOGIC;
  SIGNAL nor_685_nl : STD_LOGIC;
  SIGNAL mux_932_nl : STD_LOGIC;
  SIGNAL mux_931_nl : STD_LOGIC;
  SIGNAL mux_930_nl : STD_LOGIC;
  SIGNAL or_1259_nl : STD_LOGIC;
  SIGNAL or_1257_nl : STD_LOGIC;
  SIGNAL mux_929_nl : STD_LOGIC;
  SIGNAL or_1256_nl : STD_LOGIC;
  SIGNAL or_1254_nl : STD_LOGIC;
  SIGNAL mux_928_nl : STD_LOGIC;
  SIGNAL mux_927_nl : STD_LOGIC;
  SIGNAL or_1253_nl : STD_LOGIC;
  SIGNAL or_1251_nl : STD_LOGIC;
  SIGNAL mux_926_nl : STD_LOGIC;
  SIGNAL or_1250_nl : STD_LOGIC;
  SIGNAL or_1248_nl : STD_LOGIC;
  SIGNAL mux_956_nl : STD_LOGIC;
  SIGNAL nand_486_nl : STD_LOGIC;
  SIGNAL mux_955_nl : STD_LOGIC;
  SIGNAL and_382_nl : STD_LOGIC;
  SIGNAL mux_954_nl : STD_LOGIC;
  SIGNAL mux_953_nl : STD_LOGIC;
  SIGNAL nor_671_nl : STD_LOGIC;
  SIGNAL nor_672_nl : STD_LOGIC;
  SIGNAL mux_952_nl : STD_LOGIC;
  SIGNAL nor_673_nl : STD_LOGIC;
  SIGNAL nor_674_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL mux_951_nl : STD_LOGIC;
  SIGNAL mux_950_nl : STD_LOGIC;
  SIGNAL or_1293_nl : STD_LOGIC;
  SIGNAL or_1291_nl : STD_LOGIC;
  SIGNAL mux_949_nl : STD_LOGIC;
  SIGNAL or_1290_nl : STD_LOGIC;
  SIGNAL or_1288_nl : STD_LOGIC;
  SIGNAL or_2260_nl : STD_LOGIC;
  SIGNAL mux_948_nl : STD_LOGIC;
  SIGNAL nand_118_nl : STD_LOGIC;
  SIGNAL mux_947_nl : STD_LOGIC;
  SIGNAL mux_946_nl : STD_LOGIC;
  SIGNAL nor_677_nl : STD_LOGIC;
  SIGNAL nor_678_nl : STD_LOGIC;
  SIGNAL nor_679_nl : STD_LOGIC;
  SIGNAL mux_945_nl : STD_LOGIC;
  SIGNAL or_1282_nl : STD_LOGIC;
  SIGNAL or_1280_nl : STD_LOGIC;
  SIGNAL or_1279_nl : STD_LOGIC;
  SIGNAL mux_944_nl : STD_LOGIC;
  SIGNAL mux_943_nl : STD_LOGIC;
  SIGNAL or_1278_nl : STD_LOGIC;
  SIGNAL or_1276_nl : STD_LOGIC;
  SIGNAL or_1275_nl : STD_LOGIC;
  SIGNAL mux_972_nl : STD_LOGIC;
  SIGNAL mux_971_nl : STD_LOGIC;
  SIGNAL mux_970_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL nor_665_nl : STD_LOGIC;
  SIGNAL mux_969_nl : STD_LOGIC;
  SIGNAL nor_666_nl : STD_LOGIC;
  SIGNAL mux_965_nl : STD_LOGIC;
  SIGNAL nor_667_nl : STD_LOGIC;
  SIGNAL mux_964_nl : STD_LOGIC;
  SIGNAL nor_668_nl : STD_LOGIC;
  SIGNAL nor_669_nl : STD_LOGIC;
  SIGNAL nor_670_nl : STD_LOGIC;
  SIGNAL mux_963_nl : STD_LOGIC;
  SIGNAL mux_962_nl : STD_LOGIC;
  SIGNAL mux_961_nl : STD_LOGIC;
  SIGNAL or_1312_nl : STD_LOGIC;
  SIGNAL or_1310_nl : STD_LOGIC;
  SIGNAL mux_960_nl : STD_LOGIC;
  SIGNAL or_1309_nl : STD_LOGIC;
  SIGNAL or_1307_nl : STD_LOGIC;
  SIGNAL mux_959_nl : STD_LOGIC;
  SIGNAL mux_958_nl : STD_LOGIC;
  SIGNAL or_1306_nl : STD_LOGIC;
  SIGNAL or_1304_nl : STD_LOGIC;
  SIGNAL mux_957_nl : STD_LOGIC;
  SIGNAL or_1303_nl : STD_LOGIC;
  SIGNAL or_1301_nl : STD_LOGIC;
  SIGNAL mux_987_nl : STD_LOGIC;
  SIGNAL nand_485_nl : STD_LOGIC;
  SIGNAL mux_986_nl : STD_LOGIC;
  SIGNAL and_379_nl : STD_LOGIC;
  SIGNAL mux_985_nl : STD_LOGIC;
  SIGNAL mux_984_nl : STD_LOGIC;
  SIGNAL nor_652_nl : STD_LOGIC;
  SIGNAL nor_653_nl : STD_LOGIC;
  SIGNAL mux_983_nl : STD_LOGIC;
  SIGNAL nor_654_nl : STD_LOGIC;
  SIGNAL nor_655_nl : STD_LOGIC;
  SIGNAL nor_656_nl : STD_LOGIC;
  SIGNAL mux_982_nl : STD_LOGIC;
  SIGNAL mux_981_nl : STD_LOGIC;
  SIGNAL or_1344_nl : STD_LOGIC;
  SIGNAL or_1342_nl : STD_LOGIC;
  SIGNAL mux_980_nl : STD_LOGIC;
  SIGNAL or_1341_nl : STD_LOGIC;
  SIGNAL or_1339_nl : STD_LOGIC;
  SIGNAL or_2259_nl : STD_LOGIC;
  SIGNAL mux_979_nl : STD_LOGIC;
  SIGNAL nand_124_nl : STD_LOGIC;
  SIGNAL mux_978_nl : STD_LOGIC;
  SIGNAL mux_977_nl : STD_LOGIC;
  SIGNAL nor_658_nl : STD_LOGIC;
  SIGNAL nor_659_nl : STD_LOGIC;
  SIGNAL and_380_nl : STD_LOGIC;
  SIGNAL mux_976_nl : STD_LOGIC;
  SIGNAL nor_660_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL or_1331_nl : STD_LOGIC;
  SIGNAL mux_975_nl : STD_LOGIC;
  SIGNAL mux_974_nl : STD_LOGIC;
  SIGNAL or_1330_nl : STD_LOGIC;
  SIGNAL or_1328_nl : STD_LOGIC;
  SIGNAL nand_122_nl : STD_LOGIC;
  SIGNAL mux_1003_nl : STD_LOGIC;
  SIGNAL mux_1002_nl : STD_LOGIC;
  SIGNAL mux_1001_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL nor_647_nl : STD_LOGIC;
  SIGNAL mux_1000_nl : STD_LOGIC;
  SIGNAL and_377_nl : STD_LOGIC;
  SIGNAL mux_996_nl : STD_LOGIC;
  SIGNAL nor_648_nl : STD_LOGIC;
  SIGNAL mux_995_nl : STD_LOGIC;
  SIGNAL nor_649_nl : STD_LOGIC;
  SIGNAL nor_650_nl : STD_LOGIC;
  SIGNAL nor_651_nl : STD_LOGIC;
  SIGNAL mux_994_nl : STD_LOGIC;
  SIGNAL mux_993_nl : STD_LOGIC;
  SIGNAL mux_992_nl : STD_LOGIC;
  SIGNAL or_1363_nl : STD_LOGIC;
  SIGNAL or_1361_nl : STD_LOGIC;
  SIGNAL mux_991_nl : STD_LOGIC;
  SIGNAL or_1360_nl : STD_LOGIC;
  SIGNAL or_1358_nl : STD_LOGIC;
  SIGNAL mux_990_nl : STD_LOGIC;
  SIGNAL mux_989_nl : STD_LOGIC;
  SIGNAL or_1357_nl : STD_LOGIC;
  SIGNAL or_1355_nl : STD_LOGIC;
  SIGNAL mux_988_nl : STD_LOGIC;
  SIGNAL or_1354_nl : STD_LOGIC;
  SIGNAL or_1352_nl : STD_LOGIC;
  SIGNAL mux_1018_nl : STD_LOGIC;
  SIGNAL nand_484_nl : STD_LOGIC;
  SIGNAL mux_1017_nl : STD_LOGIC;
  SIGNAL and_376_nl : STD_LOGIC;
  SIGNAL mux_1016_nl : STD_LOGIC;
  SIGNAL mux_1015_nl : STD_LOGIC;
  SIGNAL nor_637_nl : STD_LOGIC;
  SIGNAL nor_638_nl : STD_LOGIC;
  SIGNAL mux_1014_nl : STD_LOGIC;
  SIGNAL nor_639_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL nor_641_nl : STD_LOGIC;
  SIGNAL mux_1013_nl : STD_LOGIC;
  SIGNAL mux_1012_nl : STD_LOGIC;
  SIGNAL or_1397_nl : STD_LOGIC;
  SIGNAL or_1395_nl : STD_LOGIC;
  SIGNAL mux_1011_nl : STD_LOGIC;
  SIGNAL or_1394_nl : STD_LOGIC;
  SIGNAL or_1392_nl : STD_LOGIC;
  SIGNAL or_2258_nl : STD_LOGIC;
  SIGNAL mux_1010_nl : STD_LOGIC;
  SIGNAL nand_129_nl : STD_LOGIC;
  SIGNAL mux_1009_nl : STD_LOGIC;
  SIGNAL mux_1008_nl : STD_LOGIC;
  SIGNAL nor_643_nl : STD_LOGIC;
  SIGNAL nor_644_nl : STD_LOGIC;
  SIGNAL nor_645_nl : STD_LOGIC;
  SIGNAL mux_1007_nl : STD_LOGIC;
  SIGNAL or_1386_nl : STD_LOGIC;
  SIGNAL or_1384_nl : STD_LOGIC;
  SIGNAL or_1383_nl : STD_LOGIC;
  SIGNAL mux_1006_nl : STD_LOGIC;
  SIGNAL mux_1005_nl : STD_LOGIC;
  SIGNAL or_1382_nl : STD_LOGIC;
  SIGNAL or_1380_nl : STD_LOGIC;
  SIGNAL or_1379_nl : STD_LOGIC;
  SIGNAL mux_1034_nl : STD_LOGIC;
  SIGNAL mux_1033_nl : STD_LOGIC;
  SIGNAL mux_1032_nl : STD_LOGIC;
  SIGNAL nor_630_nl : STD_LOGIC;
  SIGNAL nor_631_nl : STD_LOGIC;
  SIGNAL mux_1031_nl : STD_LOGIC;
  SIGNAL nor_632_nl : STD_LOGIC;
  SIGNAL mux_1027_nl : STD_LOGIC;
  SIGNAL nor_633_nl : STD_LOGIC;
  SIGNAL mux_1026_nl : STD_LOGIC;
  SIGNAL nor_634_nl : STD_LOGIC;
  SIGNAL nor_635_nl : STD_LOGIC;
  SIGNAL nor_636_nl : STD_LOGIC;
  SIGNAL mux_1025_nl : STD_LOGIC;
  SIGNAL mux_1024_nl : STD_LOGIC;
  SIGNAL mux_1023_nl : STD_LOGIC;
  SIGNAL or_1416_nl : STD_LOGIC;
  SIGNAL or_1414_nl : STD_LOGIC;
  SIGNAL mux_1022_nl : STD_LOGIC;
  SIGNAL or_1413_nl : STD_LOGIC;
  SIGNAL or_1411_nl : STD_LOGIC;
  SIGNAL mux_1021_nl : STD_LOGIC;
  SIGNAL mux_1020_nl : STD_LOGIC;
  SIGNAL or_1410_nl : STD_LOGIC;
  SIGNAL or_1408_nl : STD_LOGIC;
  SIGNAL mux_1019_nl : STD_LOGIC;
  SIGNAL or_1407_nl : STD_LOGIC;
  SIGNAL or_1405_nl : STD_LOGIC;
  SIGNAL mux_1049_nl : STD_LOGIC;
  SIGNAL nand_483_nl : STD_LOGIC;
  SIGNAL mux_1048_nl : STD_LOGIC;
  SIGNAL and_373_nl : STD_LOGIC;
  SIGNAL mux_1047_nl : STD_LOGIC;
  SIGNAL mux_1046_nl : STD_LOGIC;
  SIGNAL nor_618_nl : STD_LOGIC;
  SIGNAL nor_619_nl : STD_LOGIC;
  SIGNAL mux_1045_nl : STD_LOGIC;
  SIGNAL nor_620_nl : STD_LOGIC;
  SIGNAL nor_621_nl : STD_LOGIC;
  SIGNAL nor_622_nl : STD_LOGIC;
  SIGNAL mux_1044_nl : STD_LOGIC;
  SIGNAL mux_1043_nl : STD_LOGIC;
  SIGNAL or_1448_nl : STD_LOGIC;
  SIGNAL or_1446_nl : STD_LOGIC;
  SIGNAL mux_1042_nl : STD_LOGIC;
  SIGNAL or_1445_nl : STD_LOGIC;
  SIGNAL or_1443_nl : STD_LOGIC;
  SIGNAL or_2257_nl : STD_LOGIC;
  SIGNAL mux_1041_nl : STD_LOGIC;
  SIGNAL nand_135_nl : STD_LOGIC;
  SIGNAL mux_1040_nl : STD_LOGIC;
  SIGNAL mux_1039_nl : STD_LOGIC;
  SIGNAL nor_624_nl : STD_LOGIC;
  SIGNAL nor_625_nl : STD_LOGIC;
  SIGNAL and_374_nl : STD_LOGIC;
  SIGNAL mux_1038_nl : STD_LOGIC;
  SIGNAL nor_626_nl : STD_LOGIC;
  SIGNAL nor_627_nl : STD_LOGIC;
  SIGNAL or_1435_nl : STD_LOGIC;
  SIGNAL mux_1037_nl : STD_LOGIC;
  SIGNAL mux_1036_nl : STD_LOGIC;
  SIGNAL or_1434_nl : STD_LOGIC;
  SIGNAL or_1432_nl : STD_LOGIC;
  SIGNAL nand_133_nl : STD_LOGIC;
  SIGNAL mux_1065_nl : STD_LOGIC;
  SIGNAL mux_1064_nl : STD_LOGIC;
  SIGNAL mux_1063_nl : STD_LOGIC;
  SIGNAL nor_613_nl : STD_LOGIC;
  SIGNAL nor_614_nl : STD_LOGIC;
  SIGNAL mux_1062_nl : STD_LOGIC;
  SIGNAL and_370_nl : STD_LOGIC;
  SIGNAL mux_1058_nl : STD_LOGIC;
  SIGNAL and_371_nl : STD_LOGIC;
  SIGNAL mux_1057_nl : STD_LOGIC;
  SIGNAL and_526_nl : STD_LOGIC;
  SIGNAL nor_616_nl : STD_LOGIC;
  SIGNAL nor_617_nl : STD_LOGIC;
  SIGNAL mux_1056_nl : STD_LOGIC;
  SIGNAL mux_1055_nl : STD_LOGIC;
  SIGNAL mux_1054_nl : STD_LOGIC;
  SIGNAL or_1467_nl : STD_LOGIC;
  SIGNAL nand_307_nl : STD_LOGIC;
  SIGNAL mux_1053_nl : STD_LOGIC;
  SIGNAL nand_514_nl : STD_LOGIC;
  SIGNAL or_1462_nl : STD_LOGIC;
  SIGNAL mux_1052_nl : STD_LOGIC;
  SIGNAL mux_1051_nl : STD_LOGIC;
  SIGNAL or_1461_nl : STD_LOGIC;
  SIGNAL nand_310_nl : STD_LOGIC;
  SIGNAL mux_1050_nl : STD_LOGIC;
  SIGNAL nand_468_nl : STD_LOGIC;
  SIGNAL or_1456_nl : STD_LOGIC;
  SIGNAL mux_1080_nl : STD_LOGIC;
  SIGNAL nand_482_nl : STD_LOGIC;
  SIGNAL mux_1079_nl : STD_LOGIC;
  SIGNAL and_369_nl : STD_LOGIC;
  SIGNAL mux_1078_nl : STD_LOGIC;
  SIGNAL mux_1077_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL nor_605_nl : STD_LOGIC;
  SIGNAL mux_1076_nl : STD_LOGIC;
  SIGNAL nor_606_nl : STD_LOGIC;
  SIGNAL nor_607_nl : STD_LOGIC;
  SIGNAL nor_608_nl : STD_LOGIC;
  SIGNAL mux_1075_nl : STD_LOGIC;
  SIGNAL mux_1074_nl : STD_LOGIC;
  SIGNAL or_1500_nl : STD_LOGIC;
  SIGNAL or_1498_nl : STD_LOGIC;
  SIGNAL mux_1073_nl : STD_LOGIC;
  SIGNAL or_1497_nl : STD_LOGIC;
  SIGNAL or_1495_nl : STD_LOGIC;
  SIGNAL or_2256_nl : STD_LOGIC;
  SIGNAL mux_1072_nl : STD_LOGIC;
  SIGNAL nand_140_nl : STD_LOGIC;
  SIGNAL mux_1071_nl : STD_LOGIC;
  SIGNAL mux_1070_nl : STD_LOGIC;
  SIGNAL nor_610_nl : STD_LOGIC;
  SIGNAL nor_611_nl : STD_LOGIC;
  SIGNAL nor_612_nl : STD_LOGIC;
  SIGNAL mux_1069_nl : STD_LOGIC;
  SIGNAL or_1489_nl : STD_LOGIC;
  SIGNAL or_1487_nl : STD_LOGIC;
  SIGNAL or_1486_nl : STD_LOGIC;
  SIGNAL mux_1068_nl : STD_LOGIC;
  SIGNAL mux_1067_nl : STD_LOGIC;
  SIGNAL or_1485_nl : STD_LOGIC;
  SIGNAL or_1483_nl : STD_LOGIC;
  SIGNAL or_1482_nl : STD_LOGIC;
  SIGNAL mux_1096_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL mux_1094_nl : STD_LOGIC;
  SIGNAL nor_597_nl : STD_LOGIC;
  SIGNAL nor_598_nl : STD_LOGIC;
  SIGNAL mux_1093_nl : STD_LOGIC;
  SIGNAL nor_599_nl : STD_LOGIC;
  SIGNAL mux_1089_nl : STD_LOGIC;
  SIGNAL nor_600_nl : STD_LOGIC;
  SIGNAL mux_1088_nl : STD_LOGIC;
  SIGNAL nor_601_nl : STD_LOGIC;
  SIGNAL nor_602_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL mux_1087_nl : STD_LOGIC;
  SIGNAL mux_1086_nl : STD_LOGIC;
  SIGNAL mux_1085_nl : STD_LOGIC;
  SIGNAL or_1519_nl : STD_LOGIC;
  SIGNAL or_1517_nl : STD_LOGIC;
  SIGNAL mux_1084_nl : STD_LOGIC;
  SIGNAL or_1516_nl : STD_LOGIC;
  SIGNAL or_1514_nl : STD_LOGIC;
  SIGNAL mux_1083_nl : STD_LOGIC;
  SIGNAL mux_1082_nl : STD_LOGIC;
  SIGNAL or_1513_nl : STD_LOGIC;
  SIGNAL or_1511_nl : STD_LOGIC;
  SIGNAL mux_1081_nl : STD_LOGIC;
  SIGNAL or_1510_nl : STD_LOGIC;
  SIGNAL or_1508_nl : STD_LOGIC;
  SIGNAL mux_1111_nl : STD_LOGIC;
  SIGNAL nand_481_nl : STD_LOGIC;
  SIGNAL mux_1110_nl : STD_LOGIC;
  SIGNAL and_366_nl : STD_LOGIC;
  SIGNAL mux_1109_nl : STD_LOGIC;
  SIGNAL mux_1108_nl : STD_LOGIC;
  SIGNAL nor_585_nl : STD_LOGIC;
  SIGNAL nor_586_nl : STD_LOGIC;
  SIGNAL mux_1107_nl : STD_LOGIC;
  SIGNAL nor_587_nl : STD_LOGIC;
  SIGNAL nor_588_nl : STD_LOGIC;
  SIGNAL nor_589_nl : STD_LOGIC;
  SIGNAL mux_1106_nl : STD_LOGIC;
  SIGNAL mux_1105_nl : STD_LOGIC;
  SIGNAL or_1550_nl : STD_LOGIC;
  SIGNAL or_1548_nl : STD_LOGIC;
  SIGNAL mux_1104_nl : STD_LOGIC;
  SIGNAL or_1547_nl : STD_LOGIC;
  SIGNAL or_1545_nl : STD_LOGIC;
  SIGNAL or_2255_nl : STD_LOGIC;
  SIGNAL mux_1103_nl : STD_LOGIC;
  SIGNAL nand_146_nl : STD_LOGIC;
  SIGNAL mux_1102_nl : STD_LOGIC;
  SIGNAL mux_1101_nl : STD_LOGIC;
  SIGNAL nor_591_nl : STD_LOGIC;
  SIGNAL nor_592_nl : STD_LOGIC;
  SIGNAL and_367_nl : STD_LOGIC;
  SIGNAL mux_1100_nl : STD_LOGIC;
  SIGNAL nor_593_nl : STD_LOGIC;
  SIGNAL nor_594_nl : STD_LOGIC;
  SIGNAL or_1537_nl : STD_LOGIC;
  SIGNAL mux_1099_nl : STD_LOGIC;
  SIGNAL mux_1098_nl : STD_LOGIC;
  SIGNAL or_1536_nl : STD_LOGIC;
  SIGNAL or_1534_nl : STD_LOGIC;
  SIGNAL nand_144_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL mux_1125_nl : STD_LOGIC;
  SIGNAL nor_579_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL mux_1124_nl : STD_LOGIC;
  SIGNAL and_364_nl : STD_LOGIC;
  SIGNAL mux_1120_nl : STD_LOGIC;
  SIGNAL nor_581_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL nor_582_nl : STD_LOGIC;
  SIGNAL nor_583_nl : STD_LOGIC;
  SIGNAL nor_584_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL mux_1116_nl : STD_LOGIC;
  SIGNAL or_1569_nl : STD_LOGIC;
  SIGNAL or_1567_nl : STD_LOGIC;
  SIGNAL mux_1115_nl : STD_LOGIC;
  SIGNAL or_1566_nl : STD_LOGIC;
  SIGNAL or_1564_nl : STD_LOGIC;
  SIGNAL mux_1114_nl : STD_LOGIC;
  SIGNAL mux_1113_nl : STD_LOGIC;
  SIGNAL or_1563_nl : STD_LOGIC;
  SIGNAL or_1561_nl : STD_LOGIC;
  SIGNAL mux_1112_nl : STD_LOGIC;
  SIGNAL or_1560_nl : STD_LOGIC;
  SIGNAL or_1558_nl : STD_LOGIC;
  SIGNAL mux_1142_nl : STD_LOGIC;
  SIGNAL nand_480_nl : STD_LOGIC;
  SIGNAL mux_1141_nl : STD_LOGIC;
  SIGNAL and_363_nl : STD_LOGIC;
  SIGNAL mux_1140_nl : STD_LOGIC;
  SIGNAL mux_1139_nl : STD_LOGIC;
  SIGNAL nor_570_nl : STD_LOGIC;
  SIGNAL nor_571_nl : STD_LOGIC;
  SIGNAL mux_1138_nl : STD_LOGIC;
  SIGNAL nor_572_nl : STD_LOGIC;
  SIGNAL nor_573_nl : STD_LOGIC;
  SIGNAL nor_574_nl : STD_LOGIC;
  SIGNAL mux_1137_nl : STD_LOGIC;
  SIGNAL mux_1136_nl : STD_LOGIC;
  SIGNAL or_1602_nl : STD_LOGIC;
  SIGNAL or_1600_nl : STD_LOGIC;
  SIGNAL mux_1135_nl : STD_LOGIC;
  SIGNAL or_1599_nl : STD_LOGIC;
  SIGNAL or_1597_nl : STD_LOGIC;
  SIGNAL or_2254_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL nand_151_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL mux_1132_nl : STD_LOGIC;
  SIGNAL nor_576_nl : STD_LOGIC;
  SIGNAL nor_577_nl : STD_LOGIC;
  SIGNAL nor_578_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL or_1591_nl : STD_LOGIC;
  SIGNAL or_1589_nl : STD_LOGIC;
  SIGNAL or_1588_nl : STD_LOGIC;
  SIGNAL mux_1130_nl : STD_LOGIC;
  SIGNAL mux_1129_nl : STD_LOGIC;
  SIGNAL or_1587_nl : STD_LOGIC;
  SIGNAL or_1585_nl : STD_LOGIC;
  SIGNAL or_1584_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL mux_1157_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL nor_563_nl : STD_LOGIC;
  SIGNAL nor_564_nl : STD_LOGIC;
  SIGNAL mux_1155_nl : STD_LOGIC;
  SIGNAL nor_565_nl : STD_LOGIC;
  SIGNAL mux_1151_nl : STD_LOGIC;
  SIGNAL nor_566_nl : STD_LOGIC;
  SIGNAL mux_1150_nl : STD_LOGIC;
  SIGNAL nor_567_nl : STD_LOGIC;
  SIGNAL nor_568_nl : STD_LOGIC;
  SIGNAL nor_569_nl : STD_LOGIC;
  SIGNAL mux_1149_nl : STD_LOGIC;
  SIGNAL mux_1148_nl : STD_LOGIC;
  SIGNAL mux_1147_nl : STD_LOGIC;
  SIGNAL or_1621_nl : STD_LOGIC;
  SIGNAL or_1619_nl : STD_LOGIC;
  SIGNAL mux_1146_nl : STD_LOGIC;
  SIGNAL or_1618_nl : STD_LOGIC;
  SIGNAL or_1616_nl : STD_LOGIC;
  SIGNAL mux_1145_nl : STD_LOGIC;
  SIGNAL mux_1144_nl : STD_LOGIC;
  SIGNAL or_1615_nl : STD_LOGIC;
  SIGNAL or_1613_nl : STD_LOGIC;
  SIGNAL mux_1143_nl : STD_LOGIC;
  SIGNAL or_1612_nl : STD_LOGIC;
  SIGNAL or_1610_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL nand_479_nl : STD_LOGIC;
  SIGNAL mux_1172_nl : STD_LOGIC;
  SIGNAL and_360_nl : STD_LOGIC;
  SIGNAL mux_1171_nl : STD_LOGIC;
  SIGNAL mux_1170_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL mux_1169_nl : STD_LOGIC;
  SIGNAL nor_553_nl : STD_LOGIC;
  SIGNAL nor_554_nl : STD_LOGIC;
  SIGNAL nor_555_nl : STD_LOGIC;
  SIGNAL mux_1168_nl : STD_LOGIC;
  SIGNAL mux_1167_nl : STD_LOGIC;
  SIGNAL or_1651_nl : STD_LOGIC;
  SIGNAL or_1649_nl : STD_LOGIC;
  SIGNAL mux_1166_nl : STD_LOGIC;
  SIGNAL or_1648_nl : STD_LOGIC;
  SIGNAL or_1647_nl : STD_LOGIC;
  SIGNAL or_2253_nl : STD_LOGIC;
  SIGNAL mux_1165_nl : STD_LOGIC;
  SIGNAL nand_157_nl : STD_LOGIC;
  SIGNAL mux_1164_nl : STD_LOGIC;
  SIGNAL mux_1163_nl : STD_LOGIC;
  SIGNAL nor_557_nl : STD_LOGIC;
  SIGNAL nor_558_nl : STD_LOGIC;
  SIGNAL and_361_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL nor_559_nl : STD_LOGIC;
  SIGNAL nor_560_nl : STD_LOGIC;
  SIGNAL or_1639_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL or_1638_nl : STD_LOGIC;
  SIGNAL or_1636_nl : STD_LOGIC;
  SIGNAL nand_155_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL nor_546_nl : STD_LOGIC;
  SIGNAL nor_547_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL and_357_nl : STD_LOGIC;
  SIGNAL mux_1182_nl : STD_LOGIC;
  SIGNAL and_358_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL and_525_nl : STD_LOGIC;
  SIGNAL nor_549_nl : STD_LOGIC;
  SIGNAL nor_550_nl : STD_LOGIC;
  SIGNAL mux_1180_nl : STD_LOGIC;
  SIGNAL mux_1179_nl : STD_LOGIC;
  SIGNAL mux_1178_nl : STD_LOGIC;
  SIGNAL or_1670_nl : STD_LOGIC;
  SIGNAL nand_273_nl : STD_LOGIC;
  SIGNAL mux_1177_nl : STD_LOGIC;
  SIGNAL nand_513_nl : STD_LOGIC;
  SIGNAL or_1665_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL mux_1175_nl : STD_LOGIC;
  SIGNAL or_1664_nl : STD_LOGIC;
  SIGNAL nand_276_nl : STD_LOGIC;
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL nand_465_nl : STD_LOGIC;
  SIGNAL or_1659_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL nand_478_nl : STD_LOGIC;
  SIGNAL mux_1203_nl : STD_LOGIC;
  SIGNAL and_356_nl : STD_LOGIC;
  SIGNAL mux_1202_nl : STD_LOGIC;
  SIGNAL mux_1201_nl : STD_LOGIC;
  SIGNAL nor_537_nl : STD_LOGIC;
  SIGNAL nor_538_nl : STD_LOGIC;
  SIGNAL mux_1200_nl : STD_LOGIC;
  SIGNAL nor_539_nl : STD_LOGIC;
  SIGNAL nor_540_nl : STD_LOGIC;
  SIGNAL nor_541_nl : STD_LOGIC;
  SIGNAL mux_1199_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL or_1702_nl : STD_LOGIC;
  SIGNAL or_1700_nl : STD_LOGIC;
  SIGNAL mux_1197_nl : STD_LOGIC;
  SIGNAL or_1699_nl : STD_LOGIC;
  SIGNAL or_1697_nl : STD_LOGIC;
  SIGNAL or_2252_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL nand_162_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL nor_543_nl : STD_LOGIC;
  SIGNAL nor_544_nl : STD_LOGIC;
  SIGNAL nor_545_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL nand_519_nl : STD_LOGIC;
  SIGNAL or_1689_nl : STD_LOGIC;
  SIGNAL or_1688_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL or_1687_nl : STD_LOGIC;
  SIGNAL or_1685_nl : STD_LOGIC;
  SIGNAL or_1684_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL mux_1219_nl : STD_LOGIC;
  SIGNAL mux_1218_nl : STD_LOGIC;
  SIGNAL nor_530_nl : STD_LOGIC;
  SIGNAL nor_531_nl : STD_LOGIC;
  SIGNAL mux_1217_nl : STD_LOGIC;
  SIGNAL nor_532_nl : STD_LOGIC;
  SIGNAL mux_1213_nl : STD_LOGIC;
  SIGNAL nor_533_nl : STD_LOGIC;
  SIGNAL mux_1212_nl : STD_LOGIC;
  SIGNAL nor_534_nl : STD_LOGIC;
  SIGNAL nor_535_nl : STD_LOGIC;
  SIGNAL nor_536_nl : STD_LOGIC;
  SIGNAL mux_1211_nl : STD_LOGIC;
  SIGNAL mux_1210_nl : STD_LOGIC;
  SIGNAL mux_1209_nl : STD_LOGIC;
  SIGNAL or_1721_nl : STD_LOGIC;
  SIGNAL or_1719_nl : STD_LOGIC;
  SIGNAL mux_1208_nl : STD_LOGIC;
  SIGNAL or_1718_nl : STD_LOGIC;
  SIGNAL or_1716_nl : STD_LOGIC;
  SIGNAL mux_1207_nl : STD_LOGIC;
  SIGNAL mux_1206_nl : STD_LOGIC;
  SIGNAL or_1715_nl : STD_LOGIC;
  SIGNAL or_1713_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL or_1712_nl : STD_LOGIC;
  SIGNAL or_1710_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL nand_477_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL and_351_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL mux_1232_nl : STD_LOGIC;
  SIGNAL nor_520_nl : STD_LOGIC;
  SIGNAL nor_521_nl : STD_LOGIC;
  SIGNAL mux_1231_nl : STD_LOGIC;
  SIGNAL nor_522_nl : STD_LOGIC;
  SIGNAL nor_523_nl : STD_LOGIC;
  SIGNAL nor_524_nl : STD_LOGIC;
  SIGNAL mux_1230_nl : STD_LOGIC;
  SIGNAL mux_1229_nl : STD_LOGIC;
  SIGNAL or_1751_nl : STD_LOGIC;
  SIGNAL or_1749_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL or_1748_nl : STD_LOGIC;
  SIGNAL or_1746_nl : STD_LOGIC;
  SIGNAL or_2251_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL nand_168_nl : STD_LOGIC;
  SIGNAL mux_1226_nl : STD_LOGIC;
  SIGNAL mux_1225_nl : STD_LOGIC;
  SIGNAL nor_526_nl : STD_LOGIC;
  SIGNAL nor_527_nl : STD_LOGIC;
  SIGNAL and_352_nl : STD_LOGIC;
  SIGNAL mux_1224_nl : STD_LOGIC;
  SIGNAL and_524_nl : STD_LOGIC;
  SIGNAL nor_529_nl : STD_LOGIC;
  SIGNAL or_1738_nl : STD_LOGIC;
  SIGNAL mux_1223_nl : STD_LOGIC;
  SIGNAL mux_1222_nl : STD_LOGIC;
  SIGNAL nand_512_nl : STD_LOGIC;
  SIGNAL or_1735_nl : STD_LOGIC;
  SIGNAL nand_166_nl : STD_LOGIC;
  SIGNAL mux_1251_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL mux_1248_nl : STD_LOGIC;
  SIGNAL and_348_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL and_349_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL and_523_nl : STD_LOGIC;
  SIGNAL nor_518_nl : STD_LOGIC;
  SIGNAL nor_519_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL or_1768_nl : STD_LOGIC;
  SIGNAL nand_251_nl : STD_LOGIC;
  SIGNAL mux_1239_nl : STD_LOGIC;
  SIGNAL nand_511_nl : STD_LOGIC;
  SIGNAL or_1763_nl : STD_LOGIC;
  SIGNAL mux_1238_nl : STD_LOGIC;
  SIGNAL mux_1237_nl : STD_LOGIC;
  SIGNAL or_1762_nl : STD_LOGIC;
  SIGNAL nand_254_nl : STD_LOGIC;
  SIGNAL mux_1236_nl : STD_LOGIC;
  SIGNAL nand_462_nl : STD_LOGIC;
  SIGNAL or_1758_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL nand_476_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL and_347_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL and_529_nl : STD_LOGIC;
  SIGNAL nor_507_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL and_530_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL or_1796_nl : STD_LOGIC;
  SIGNAL or_1795_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL nand_510_nl : STD_LOGIC;
  SIGNAL or_1792_nl : STD_LOGIC;
  SIGNAL or_2250_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL nand_173_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL and_531_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL nand_243_nl : STD_LOGIC;
  SIGNAL nand_244_nl : STD_LOGIC;
  SIGNAL or_1785_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL or_1784_nl : STD_LOGIC;
  SIGNAL or_1783_nl : STD_LOGIC;
  SIGNAL or_1782_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL mux_1281_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL nor_501_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL and_345_nl : STD_LOGIC;
  SIGNAL mux_1274_nl : STD_LOGIC;
  SIGNAL and_522_nl : STD_LOGIC;
  SIGNAL nor_504_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL mux_1273_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL or_1815_nl : STD_LOGIC;
  SIGNAL nand_231_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL nand_509_nl : STD_LOGIC;
  SIGNAL or_1810_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL or_1809_nl : STD_LOGIC;
  SIGNAL nand_234_nl : STD_LOGIC;
  SIGNAL mux_1267_nl : STD_LOGIC;
  SIGNAL nand_460_nl : STD_LOGIC;
  SIGNAL or_1804_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL nand_475_nl : STD_LOGIC;
  SIGNAL mux_1296_nl : STD_LOGIC;
  SIGNAL and_333_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL mux_1294_nl : STD_LOGIC;
  SIGNAL and_334_nl : STD_LOGIC;
  SIGNAL and_335_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL and_336_nl : STD_LOGIC;
  SIGNAL and_337_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL mux_1292_nl : STD_LOGIC;
  SIGNAL mux_1291_nl : STD_LOGIC;
  SIGNAL nand_223_nl : STD_LOGIC;
  SIGNAL nand_224_nl : STD_LOGIC;
  SIGNAL mux_1290_nl : STD_LOGIC;
  SIGNAL nand_225_nl : STD_LOGIC;
  SIGNAL nand_226_nl : STD_LOGIC;
  SIGNAL or_2249_nl : STD_LOGIC;
  SIGNAL mux_1289_nl : STD_LOGIC;
  SIGNAL nand_179_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL mux_1287_nl : STD_LOGIC;
  SIGNAL and_338_nl : STD_LOGIC;
  SIGNAL and_339_nl : STD_LOGIC;
  SIGNAL and_340_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL and_341_nl : STD_LOGIC;
  SIGNAL and_342_nl : STD_LOGIC;
  SIGNAL or_1830_nl : STD_LOGIC;
  SIGNAL mux_1285_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL nand_227_nl : STD_LOGIC;
  SIGNAL nand_228_nl : STD_LOGIC;
  SIGNAL nand_177_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL nor_495_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL and_329_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL and_330_nl : STD_LOGIC;
  SIGNAL mux_1305_nl : STD_LOGIC;
  SIGNAL and_521_nl : STD_LOGIC;
  SIGNAL and_331_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL mux_1303_nl : STD_LOGIC;
  SIGNAL mux_1302_nl : STD_LOGIC;
  SIGNAL or_1848_nl : STD_LOGIC;
  SIGNAL nand_214_nl : STD_LOGIC;
  SIGNAL mux_1301_nl : STD_LOGIC;
  SIGNAL nand_508_nl : STD_LOGIC;
  SIGNAL nand_216_nl : STD_LOGIC;
  SIGNAL mux_1300_nl : STD_LOGIC;
  SIGNAL mux_1299_nl : STD_LOGIC;
  SIGNAL nand_217_nl : STD_LOGIC;
  SIGNAL nand_218_nl : STD_LOGIC;
  SIGNAL mux_1298_nl : STD_LOGIC;
  SIGNAL nand_458_nl : STD_LOGIC;
  SIGNAL nand_220_nl : STD_LOGIC;
  SIGNAL mux_1320_nl : STD_LOGIC;
  SIGNAL mux_1319_nl : STD_LOGIC;
  SIGNAL mux_1318_nl : STD_LOGIC;
  SIGNAL nor_486_nl : STD_LOGIC;
  SIGNAL nor_487_nl : STD_LOGIC;
  SIGNAL mux_1317_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL mux_1316_nl : STD_LOGIC;
  SIGNAL mux_1315_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL nor_492_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL nor_483_nl : STD_LOGIC;
  SIGNAL nor_484_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL or_1872_nl : STD_LOGIC;
  SIGNAL or_1870_nl : STD_LOGIC;
  SIGNAL mux_1328_nl : STD_LOGIC;
  SIGNAL mux_1327_nl : STD_LOGIC;
  SIGNAL nor_477_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL mux_1326_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL mux_1331_nl : STD_LOGIC;
  SIGNAL mux_1330_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL nor_476_nl : STD_LOGIC;
  SIGNAL mux_1329_nl : STD_LOGIC;
  SIGNAL or_1886_nl : STD_LOGIC;
  SIGNAL or_1884_nl : STD_LOGIC;
  SIGNAL mux_1337_nl : STD_LOGIC;
  SIGNAL mux_1336_nl : STD_LOGIC;
  SIGNAL mux_1335_nl : STD_LOGIC;
  SIGNAL nor_467_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL mux_1334_nl : STD_LOGIC;
  SIGNAL mux_1333_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL nor_471_nl : STD_LOGIC;
  SIGNAL mux_1332_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL nor_473_nl : STD_LOGIC;
  SIGNAL mux_1340_nl : STD_LOGIC;
  SIGNAL mux_1339_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL nor_465_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL mux_1338_nl : STD_LOGIC;
  SIGNAL or_1902_nl : STD_LOGIC;
  SIGNAL or_1900_nl : STD_LOGIC;
  SIGNAL mux_1345_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL nor_459_nl : STD_LOGIC;
  SIGNAL mux_1343_nl : STD_LOGIC;
  SIGNAL mux_1342_nl : STD_LOGIC;
  SIGNAL mux_1341_nl : STD_LOGIC;
  SIGNAL mux_1348_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL nor_457_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL or_1916_nl : STD_LOGIC;
  SIGNAL or_1914_nl : STD_LOGIC;
  SIGNAL mux_1355_nl : STD_LOGIC;
  SIGNAL mux_1354_nl : STD_LOGIC;
  SIGNAL mux_1353_nl : STD_LOGIC;
  SIGNAL nor_447_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL mux_1352_nl : STD_LOGIC;
  SIGNAL nor_449_nl : STD_LOGIC;
  SIGNAL mux_1351_nl : STD_LOGIC;
  SIGNAL mux_1350_nl : STD_LOGIC;
  SIGNAL nor_451_nl : STD_LOGIC;
  SIGNAL mux_1349_nl : STD_LOGIC;
  SIGNAL nor_453_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL mux_1358_nl : STD_LOGIC;
  SIGNAL mux_1357_nl : STD_LOGIC;
  SIGNAL nor_444_nl : STD_LOGIC;
  SIGNAL nor_445_nl : STD_LOGIC;
  SIGNAL nor_446_nl : STD_LOGIC;
  SIGNAL mux_1356_nl : STD_LOGIC;
  SIGNAL or_1933_nl : STD_LOGIC;
  SIGNAL or_1931_nl : STD_LOGIC;
  SIGNAL mux_1363_nl : STD_LOGIC;
  SIGNAL mux_1362_nl : STD_LOGIC;
  SIGNAL nor_438_nl : STD_LOGIC;
  SIGNAL nor_439_nl : STD_LOGIC;
  SIGNAL mux_1361_nl : STD_LOGIC;
  SIGNAL mux_1360_nl : STD_LOGIC;
  SIGNAL mux_1359_nl : STD_LOGIC;
  SIGNAL mux_1366_nl : STD_LOGIC;
  SIGNAL mux_1365_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL nor_436_nl : STD_LOGIC;
  SIGNAL nor_437_nl : STD_LOGIC;
  SIGNAL mux_1364_nl : STD_LOGIC;
  SIGNAL or_1947_nl : STD_LOGIC;
  SIGNAL or_1945_nl : STD_LOGIC;
  SIGNAL mux_1372_nl : STD_LOGIC;
  SIGNAL mux_1371_nl : STD_LOGIC;
  SIGNAL mux_1370_nl : STD_LOGIC;
  SIGNAL nor_428_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL mux_1369_nl : STD_LOGIC;
  SIGNAL mux_1368_nl : STD_LOGIC;
  SIGNAL nor_431_nl : STD_LOGIC;
  SIGNAL nor_432_nl : STD_LOGIC;
  SIGNAL mux_1367_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL nor_434_nl : STD_LOGIC;
  SIGNAL mux_1375_nl : STD_LOGIC;
  SIGNAL mux_1374_nl : STD_LOGIC;
  SIGNAL nor_425_nl : STD_LOGIC;
  SIGNAL nor_426_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL mux_1373_nl : STD_LOGIC;
  SIGNAL or_1963_nl : STD_LOGIC;
  SIGNAL or_1961_nl : STD_LOGIC;
  SIGNAL mux_1380_nl : STD_LOGIC;
  SIGNAL mux_1379_nl : STD_LOGIC;
  SIGNAL nor_419_nl : STD_LOGIC;
  SIGNAL nor_420_nl : STD_LOGIC;
  SIGNAL mux_1378_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL mux_1376_nl : STD_LOGIC;
  SIGNAL mux_1383_nl : STD_LOGIC;
  SIGNAL mux_1382_nl : STD_LOGIC;
  SIGNAL nor_416_nl : STD_LOGIC;
  SIGNAL nor_417_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL mux_1381_nl : STD_LOGIC;
  SIGNAL or_1977_nl : STD_LOGIC;
  SIGNAL or_1975_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL mux_1389_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL nor_408_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL mux_1387_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL mux_1386_nl : STD_LOGIC;
  SIGNAL mux_1385_nl : STD_LOGIC;
  SIGNAL nor_412_nl : STD_LOGIC;
  SIGNAL mux_1384_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL nor_415_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL nor_406_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL or_1994_nl : STD_LOGIC;
  SIGNAL or_1992_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL mux_1397_nl : STD_LOGIC;
  SIGNAL nor_399_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL nor_396_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL nor_398_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL or_2008_nl : STD_LOGIC;
  SIGNAL or_2006_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL nor_389_nl : STD_LOGIC;
  SIGNAL nor_390_nl : STD_LOGIC;
  SIGNAL nor_391_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL nor_392_nl : STD_LOGIC;
  SIGNAL nor_393_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL nor_394_nl : STD_LOGIC;
  SIGNAL nor_395_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL nor_387_nl : STD_LOGIC;
  SIGNAL nor_388_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL or_2024_nl : STD_LOGIC;
  SIGNAL or_2022_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL mux_1414_nl : STD_LOGIC;
  SIGNAL nor_380_nl : STD_LOGIC;
  SIGNAL nor_381_nl : STD_LOGIC;
  SIGNAL mux_1413_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL mux_1418_nl : STD_LOGIC;
  SIGNAL mux_1417_nl : STD_LOGIC;
  SIGNAL nor_377_nl : STD_LOGIC;
  SIGNAL nor_378_nl : STD_LOGIC;
  SIGNAL nor_379_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL or_2038_nl : STD_LOGIC;
  SIGNAL or_2036_nl : STD_LOGIC;
  SIGNAL mux_1425_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL nor_369_nl : STD_LOGIC;
  SIGNAL nor_370_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL nor_371_nl : STD_LOGIC;
  SIGNAL mux_1421_nl : STD_LOGIC;
  SIGNAL mux_1420_nl : STD_LOGIC;
  SIGNAL nor_373_nl : STD_LOGIC;
  SIGNAL mux_1419_nl : STD_LOGIC;
  SIGNAL nor_375_nl : STD_LOGIC;
  SIGNAL nor_376_nl : STD_LOGIC;
  SIGNAL mux_1428_nl : STD_LOGIC;
  SIGNAL mux_1427_nl : STD_LOGIC;
  SIGNAL nor_366_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL nor_368_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL or_2054_nl : STD_LOGIC;
  SIGNAL or_2052_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL nor_360_nl : STD_LOGIC;
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL mux_1436_nl : STD_LOGIC;
  SIGNAL mux_1435_nl : STD_LOGIC;
  SIGNAL nor_357_nl : STD_LOGIC;
  SIGNAL nor_358_nl : STD_LOGIC;
  SIGNAL nor_359_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL or_2067_nl : STD_LOGIC;
  SIGNAL or_2066_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL mux_1441_nl : STD_LOGIC;
  SIGNAL mux_1440_nl : STD_LOGIC;
  SIGNAL nor_351_nl : STD_LOGIC;
  SIGNAL nor_352_nl : STD_LOGIC;
  SIGNAL nor_353_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL nor_354_nl : STD_LOGIC;
  SIGNAL nor_355_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL and_328_nl : STD_LOGIC;
  SIGNAL nor_356_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL and_327_nl : STD_LOGIC;
  SIGNAL nor_349_nl : STD_LOGIC;
  SIGNAL nor_350_nl : STD_LOGIC;
  SIGNAL mux_1443_nl : STD_LOGIC;
  SIGNAL nand_474_nl : STD_LOGIC;
  SIGNAL or_2080_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL and_323_nl : STD_LOGIC;
  SIGNAL and_324_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL and_321_nl : STD_LOGIC;
  SIGNAL and_322_nl : STD_LOGIC;
  SIGNAL nor_346_nl : STD_LOGIC;
  SIGNAL mux_1451_nl : STD_LOGIC;
  SIGNAL nand_192_nl : STD_LOGIC;
  SIGNAL nand_193_nl : STD_LOGIC;
  SIGNAL nand_520_nl : STD_LOGIC;
  SIGNAL mux_1600_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_382_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL and_755_nl : STD_LOGIC;
  SIGNAL acc_1_nl : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_383_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nand_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_384_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL STAGE_LOOP_mux_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_94_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_or_76_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_161_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_95_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_or_77_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_78_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_mux_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_96_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_756_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux_22_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_or_79_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_657_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_658_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_930_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_931_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_932_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_933_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_934_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_935_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_936_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_659_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_937_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_938_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_939_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_940_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_941_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_942_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_943_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_660_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_661_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_944_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_945_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_946_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_947_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_948_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_949_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_950_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_662_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_663_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_664_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_665_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_951_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_952_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_953_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_954_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_955_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_956_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_957_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_666_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_667_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_668_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_669_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_670_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_671_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_672_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_673_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_958_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_959_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_960_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_961_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_962_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_963_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_964_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_674_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_675_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_676_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_677_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_678_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_679_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_680_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_681_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_682_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_683_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_684_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_685_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_686_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_687_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_688_nl : STD_LOGIC;
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT modulo_dev
    PORT (
      base_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1 : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat : STD_LOGIC;

  SIGNAL COMP_LOOP_5_tmp_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL COMP_LOOP_5_tmp_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_5_tmp_lshift_rg_z : STD_LOGIC_VECTOR (10 DOWNTO 0);

  SIGNAL COMP_LOOP_1_tmp_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_lshift_rg_z : STD_LOGIC_VECTOR (9 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_core_wait_dp
    PORT(
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      COMP_LOOP_C_28_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_56_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_84_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_112_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_140_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_168_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_196_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_224_tr0 : IN STD_LOGIC;
      VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_1_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_5_2(input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_8_2(input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_16_2(input_15 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_6_2(input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_7_2(input_6 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_16_2(input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_32_2(input_31 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(31 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_33_2(input_32 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(32 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
      tmp := (OTHERS=>sel( 32));
      result := result or ( input_32 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_36_2(input_35 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_34 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_33 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_32 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(35 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
      tmp := (OTHERS=>sel( 32));
      result := result or ( input_32 and tmp);
      tmp := (OTHERS=>sel( 33));
      result := result or ( input_33 and tmp);
      tmp := (OTHERS=>sel( 34));
      result := result or ( input_34 and tmp);
      tmp := (OTHERS=>sel( 35));
      result := result or ( input_35 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_3_2(input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_4_2(input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_8_2(input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_9_2(input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_3_2(input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_9_4_2(input_3 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_11_2_2(input_0 : STD_LOGIC_VECTOR(10 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(10 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(10 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_9_2_2(input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION minimum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1<arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION maximum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1>arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION READSLICE_64_65(input_val:STD_LOGIC_VECTOR(64 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC_VECTOR IS
    CONSTANT min_sat_index:INTEGER:= maximum( index, 0 );
    CONSTANT sat_index:INTEGER:= minimum( min_sat_index, 1);
  BEGIN
    RETURN input_val(sat_index+63 DOWNTO sat_index);
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 5,
      width => 64
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  vec_rsc_triosy_0_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_31_lz
    );
  vec_rsc_triosy_0_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_30_lz
    );
  vec_rsc_triosy_0_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_29_lz
    );
  vec_rsc_triosy_0_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_28_lz
    );
  vec_rsc_triosy_0_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_27_lz
    );
  vec_rsc_triosy_0_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_26_lz
    );
  vec_rsc_triosy_0_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_25_lz
    );
  vec_rsc_triosy_0_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_24_lz
    );
  vec_rsc_triosy_0_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_23_lz
    );
  vec_rsc_triosy_0_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_22_lz
    );
  vec_rsc_triosy_0_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_21_lz
    );
  vec_rsc_triosy_0_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_20_lz
    );
  vec_rsc_triosy_0_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_19_lz
    );
  vec_rsc_triosy_0_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_18_lz
    );
  vec_rsc_triosy_0_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_17_lz
    );
  vec_rsc_triosy_0_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_16_lz
    );
  vec_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_15_lz
    );
  vec_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_14_lz
    );
  vec_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_13_lz
    );
  vec_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_12_lz
    );
  vec_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_11_lz
    );
  vec_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_10_lz
    );
  vec_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_9_lz
    );
  vec_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_8_lz
    );
  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_7_lz
    );
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_6_lz
    );
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_5_lz
    );
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_4_lz
    );
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_3_lz
    );
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_2_lz
    );
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_1_lz
    );
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => vec_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  twiddle_rsc_triosy_0_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_31_lz
    );
  twiddle_rsc_triosy_0_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_30_lz
    );
  twiddle_rsc_triosy_0_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_29_lz
    );
  twiddle_rsc_triosy_0_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_28_lz
    );
  twiddle_rsc_triosy_0_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_27_lz
    );
  twiddle_rsc_triosy_0_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_26_lz
    );
  twiddle_rsc_triosy_0_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_25_lz
    );
  twiddle_rsc_triosy_0_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_24_lz
    );
  twiddle_rsc_triosy_0_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_23_lz
    );
  twiddle_rsc_triosy_0_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_22_lz
    );
  twiddle_rsc_triosy_0_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_21_lz
    );
  twiddle_rsc_triosy_0_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_20_lz
    );
  twiddle_rsc_triosy_0_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_19_lz
    );
  twiddle_rsc_triosy_0_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_18_lz
    );
  twiddle_rsc_triosy_0_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_17_lz
    );
  twiddle_rsc_triosy_0_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_16_lz
    );
  twiddle_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_15_lz
    );
  twiddle_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_14_lz
    );
  twiddle_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_13_lz
    );
  twiddle_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_12_lz
    );
  twiddle_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_11_lz
    );
  twiddle_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_10_lz
    );
  twiddle_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_9_lz
    );
  twiddle_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_8_lz
    );
  twiddle_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_7_lz
    );
  twiddle_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_6_lz
    );
  twiddle_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_5_lz
    );
  twiddle_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_4_lz
    );
  twiddle_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_3_lz
    );
  twiddle_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_2_lz
    );
  twiddle_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_1_lz
    );
  twiddle_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_31_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_0_lz
    );
  COMP_LOOP_1_modulo_dev_cmp : modulo_dev
    PORT MAP(
      base_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat,
      m_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat,
      return_rsc_z => COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1,
      ccs_ccore_start_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => clk,
      ccs_ccore_srst => rst,
      ccs_ccore_en => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
    );
  COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat <= MUX1HOT_v_64_3_2((READSLICE_64_65(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_385_cse
      & '1') + UNSIGNED((MUX_v_64_2_2((NOT COMP_LOOP_1_acc_8_itm), (NOT z_out_9),
      COMP_LOOP_or_33_itm)) & '1'), 65)), 1)), COMP_LOOP_1_acc_8_itm, z_out_8, STD_LOGIC_VECTOR'(
      COMP_LOOP_or_36_itm & ((NOT (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((NOT and_449_cse),
      mux_tmp_1430, fsm_output(4))), or_tmp_2025, fsm_output(2))), (MUX_s_1_2_2(or_tmp_2025,
      (MUX_s_1_2_2(((NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7)))),
      mux_tmp_1423, fsm_output(4))), fsm_output(2))), fsm_output(5)))) AND and_dcpl_40)
      & ((and_dcpl_33 AND and_dcpl_220) OR (and_dcpl_33 AND and_dcpl_223) OR (and_dcpl_89
      AND and_dcpl_175) OR (and_dcpl_89 AND and_dcpl_36) OR (and_dcpl_95 AND and_dcpl_30)
      OR (and_dcpl_95 AND and_dcpl_52) OR (and_dcpl_95 AND and_dcpl_56) OR (and_dcpl_38
      AND and_dcpl_60))));
  COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat <= p_sva;
  COMP_LOOP_1_modulo_dev_cmp_return_rsc_z <= COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1;
  COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat <= NOT((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(((fsm_output(3))
      OR (NOT (MUX_s_1_2_2(or_145_cse, and_490_cse, fsm_output(0))))), nand_tmp_184,
      fsm_output(6))), ((fsm_output(6)) OR mux_tmp_1437), fsm_output(5))), (MUX_s_1_2_2((MUX_s_1_2_2(mux_tmp_1437,
      ((fsm_output(3)) OR (fsm_output(0)) OR (NOT and_490_cse)), fsm_output(6))),
      (MUX_s_1_2_2(nand_tmp_184, ((fsm_output(3)) OR (NOT((NOT (fsm_output(0))) OR
      (fsm_output(4)))) OR (fsm_output(7))), fsm_output(6))), fsm_output(5))), fsm_output(2)))
      OR (fsm_output(1)));

  COMP_LOOP_5_tmp_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 11
      )
    PORT MAP(
      a => COMP_LOOP_5_tmp_lshift_rg_a,
      s => COMP_LOOP_5_tmp_lshift_rg_s,
      z => COMP_LOOP_5_tmp_lshift_rg_z
    );
  COMP_LOOP_5_tmp_lshift_rg_a(0) <= '1';
  COMP_LOOP_5_tmp_lshift_rg_s <= MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, z_out_4, CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("00000010")));
  z_out <= COMP_LOOP_5_tmp_lshift_rg_z;

  COMP_LOOP_1_tmp_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 10
      )
    PORT MAP(
      a => COMP_LOOP_1_tmp_lshift_rg_a,
      s => COMP_LOOP_1_tmp_lshift_rg_s,
      z => COMP_LOOP_1_tmp_lshift_rg_z
    );
  COMP_LOOP_1_tmp_lshift_rg_a(0) <= '1';
  COMP_LOOP_1_tmp_lshift_rg_s <= MUX_v_4_2_2(z_out_4, COMP_LOOP_1_tmp_acc_cse_sva,
      (nor_1025_cse AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND and_dcpl_29 AND (NOT (fsm_output(2))) AND (NOT (fsm_output(5)))) OR (nor_1025_cse
      AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("00")) AND and_dcpl_29
      AND (fsm_output(2)) AND (NOT (fsm_output(5)))));
  z_out_1 <= COMP_LOOP_1_tmp_lshift_rg_z;

  inPlaceNTT_DIF_core_wait_dp_inst : inPlaceNTT_DIF_core_wait_dp
    PORT MAP(
      ensig_cgo_iro => mux_1462_rmff,
      ensig_cgo => reg_ensig_cgo_cse,
      COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
    );
  inPlaceNTT_DIF_core_core_fsm_inst : inPlaceNTT_DIF_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => inPlaceNTT_DIF_core_core_fsm_inst_fsm_output,
      COMP_LOOP_C_28_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0,
      COMP_LOOP_C_56_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0,
      COMP_LOOP_C_84_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0,
      COMP_LOOP_C_112_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0,
      COMP_LOOP_C_140_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0,
      COMP_LOOP_C_168_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0,
      COMP_LOOP_C_196_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0,
      COMP_LOOP_C_224_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0,
      VEC_LOOP_C_0_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_1_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0
    );
  fsm_output <= inPlaceNTT_DIF_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0 <= NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0 <= NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0 <= NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0 <= NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0 <= NOT COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 <= z_out_3(10);
  inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 <= NOT (z_out_2(4));

  and_449_cse <= (fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(7));
  or_285_cse <= (NOT (fsm_output(4))) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_347_nl <= MUX_s_1_2_2(or_285_cse, mux_tmp_311, fsm_output(3));
  nand_11_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_311));
  mux_348_cse <= MUX_s_1_2_2(mux_347_nl, nand_11_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_443_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")));
  nand_444_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(0)) AND CONV_SL_1_1(fsm_output(7
      DOWNTO 6)=STD_LOGIC_VECTOR'("11")));
  nand_22_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_373));
  mux_409_nl <= MUX_s_1_2_2(or_285_cse, mux_tmp_373, fsm_output(3));
  mux_410_cse <= MUX_s_1_2_2(nand_22_nl, mux_409_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  or_493_cse <= (NOT (fsm_output(4))) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_471_nl <= MUX_s_1_2_2(or_493_cse, mux_tmp_435, fsm_output(3));
  nand_33_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_435));
  mux_472_cse <= MUX_s_1_2_2(mux_471_nl, nand_33_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_44_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_497));
  mux_533_nl <= MUX_s_1_2_2(or_493_cse, mux_tmp_497, fsm_output(3));
  mux_534_cse <= MUX_s_1_2_2(nand_44_nl, mux_533_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  or_701_cse <= (NOT (fsm_output(4))) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_595_nl <= MUX_s_1_2_2(or_701_cse, mux_tmp_559, fsm_output(3));
  nand_55_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_559));
  mux_596_cse <= MUX_s_1_2_2(mux_595_nl, nand_55_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_66_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_621));
  mux_657_nl <= MUX_s_1_2_2(or_701_cse, mux_tmp_621, fsm_output(3));
  mux_658_cse <= MUX_s_1_2_2(nand_66_nl, mux_657_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_394_cse <= NOT((fsm_output(4)) AND CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("011")) AND COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_719_nl <= MUX_s_1_2_2(nand_394_cse, mux_tmp_683, fsm_output(3));
  nand_77_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_683));
  mux_720_cse <= MUX_s_1_2_2(mux_719_nl, nand_77_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_88_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_745));
  mux_781_nl <= MUX_s_1_2_2(nand_394_cse, mux_tmp_745, fsm_output(3));
  mux_782_cse <= MUX_s_1_2_2(nand_88_nl, mux_781_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_371_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)=STD_LOGIC_VECTOR'("0111")));
  or_1066_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_365_cse;
  or_1064_nl <= (COMP_LOOP_acc_psp_sva(0)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR (NOT
      (COMP_LOOP_acc_psp_sva(1))) OR (fsm_output(7));
  mux_818_cse <= MUX_s_1_2_2(or_1066_nl, or_1064_nl, fsm_output(4));
  or_1113_cse <= (NOT (fsm_output(4))) OR CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_843_nl <= MUX_s_1_2_2(or_1113_cse, mux_tmp_807, fsm_output(3));
  nand_99_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_807));
  mux_844_cse <= MUX_s_1_2_2(mux_843_nl, nand_99_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nor_730_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_365_cse);
  nor_731_nl <= NOT((COMP_LOOP_acc_psp_sva(0)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR
      (NOT (COMP_LOOP_acc_psp_sva(1))) OR (fsm_output(7)));
  mux_849_cse <= MUX_s_1_2_2(nor_730_nl, nor_731_nl, fsm_output(4));
  nand_356_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_sva(0))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")));
  nand_110_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_869));
  mux_905_nl <= MUX_s_1_2_2(or_1113_cse, mux_tmp_869, fsm_output(3));
  mux_906_cse <= MUX_s_1_2_2(nand_110_nl, mux_905_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  or_1274_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_365_cse;
  or_1272_nl <= (COMP_LOOP_acc_psp_sva(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (NOT (COMP_LOOP_acc_psp_sva(1))) OR (fsm_output(7));
  mux_942_cse <= MUX_s_1_2_2(or_1274_nl, or_1272_nl, fsm_output(4));
  nand_336_cse <= NOT((fsm_output(4)) AND CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("101")) AND COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_967_nl <= MUX_s_1_2_2(nand_336_cse, mux_tmp_931, fsm_output(3));
  nand_121_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_931));
  mux_968_cse <= MUX_s_1_2_2(mux_967_nl, nand_121_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nor_662_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_365_cse);
  nor_663_nl <= NOT((COMP_LOOP_acc_psp_sva(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (NOT (COMP_LOOP_acc_psp_sva(1))) OR (fsm_output(7)));
  mux_973_cse <= MUX_s_1_2_2(nor_662_nl, nor_663_nl, fsm_output(4));
  nand_132_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_993));
  mux_1029_nl <= MUX_s_1_2_2(nand_336_cse, mux_tmp_993, fsm_output(3));
  mux_1030_cse <= MUX_s_1_2_2(nand_132_nl, mux_1029_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  or_1481_nl <= (COMP_LOOP_acc_13_psp_sva(0)) OR nand_303_cse;
  or_1480_nl <= (NOT (COMP_LOOP_acc_psp_sva(0))) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR (NOT (COMP_LOOP_acc_psp_sva(1))) OR (fsm_output(7));
  mux_1066_cse <= MUX_s_1_2_2(or_1481_nl, or_1480_nl, fsm_output(4));
  nand_300_cse <= NOT((fsm_output(4)) AND CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("110")) AND COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_1091_nl <= MUX_s_1_2_2(nand_300_cse, mux_tmp_1055, fsm_output(3));
  nand_143_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_1055));
  mux_1092_cse <= MUX_s_1_2_2(mux_1091_nl, nand_143_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nor_595_nl <= NOT((COMP_LOOP_acc_13_psp_sva(0)) OR nand_303_cse);
  nor_596_nl <= NOT((NOT (COMP_LOOP_acc_psp_sva(0))) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR (NOT (COMP_LOOP_acc_psp_sva(1))) OR (fsm_output(7)));
  mux_1097_cse <= MUX_s_1_2_2(nor_595_nl, nor_596_nl, fsm_output(4));
  nand_293_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_sva(4))
      AND (COMP_LOOP_acc_10_cse_10_1_sva(0)) AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("11")));
  nand_154_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_1117));
  mux_1153_nl <= MUX_s_1_2_2(nand_300_cse, mux_tmp_1117, fsm_output(3));
  mux_1154_cse <= MUX_s_1_2_2(nand_154_nl, mux_1153_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_264_cse <= NOT((fsm_output(4)) AND CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_1215_nl <= MUX_s_1_2_2(nand_264_cse, mux_tmp_1179, fsm_output(3));
  nand_165_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_1179));
  mux_1216_cse <= MUX_s_1_2_2(mux_1215_nl, nand_165_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_176_nl <= NOT((fsm_output(3)) AND (NOT mux_tmp_1241));
  mux_1277_nl <= MUX_s_1_2_2(nand_264_cse, mux_tmp_1241, fsm_output(3));
  mux_1278_cse <= MUX_s_1_2_2(nand_176_nl, mux_1277_nl, VEC_LOOP_j_10_0_sva_9_0(1));
  nand_204_cse <= NOT((COMP_LOOP_3_tmp_lshift_ncse_sva(3)) AND (fsm_output(3)));
  nand_205_cse <= NOT((COMP_LOOP_2_tmp_lshift_ncse_sva(4)) AND (fsm_output(3)));
  mux_1460_nl <= MUX_s_1_2_2(mux_tmp_1424, mux_tmp_1423, fsm_output(4));
  mux_1461_nl <= MUX_s_1_2_2(or_tmp_2025, mux_1460_nl, fsm_output(2));
  mux_1455_nl <= MUX_s_1_2_2((fsm_output(6)), mux_189_cse, fsm_output(3));
  mux_1456_nl <= MUX_s_1_2_2(and_456_cse, mux_1455_nl, fsm_output(4));
  mux_1457_nl <= MUX_s_1_2_2(mux_1456_nl, and_464_cse, fsm_output(2));
  mux_1462_rmff <= MUX_s_1_2_2(mux_1461_nl, (NOT mux_1457_nl), fsm_output(5));
  or_220_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"));
  or_212_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  and_316_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  nor_1023_cse <= NOT((fsm_output(2)) OR (fsm_output(4)));
  and_496_cse <= (fsm_output(1)) AND (fsm_output(3));
  or_32_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse <= NOT(CONV_SL_1_1(z_out_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  and_491_cse <= ((fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(3))) AND (fsm_output(7));
  mux_189_cse <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(6));
  and_33_cse <= (fsm_output(6)) AND or_212_cse AND (fsm_output(7));
  and_464_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  COMP_LOOP_tmp_or_cse <= and_dcpl_46 OR and_dcpl_49 OR and_dcpl_171 OR and_dcpl_172
      OR and_dcpl_173 OR and_dcpl_176;
  COMP_LOOP_or_59_cse <= and_dcpl_172 OR and_dcpl_176;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
  COMP_LOOP_tmp_nor_27_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse <= CONV_SL_1_1(z_out_7(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_nor_27_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
  COMP_LOOP_tmp_nor_29_cse <= NOT((z_out_7(3)) OR (z_out_7(1)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_cse <= (z_out_7(2)) AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_29_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
  COMP_LOOP_tmp_nor_78_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse <= (z_out_7(4)) AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_78_cse;
  COMP_LOOP_tmp_nor_30_cse <= NOT((z_out_7(3)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse <= CONV_SL_1_1(z_out_7(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_nor_30_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01100"));
  COMP_LOOP_tmp_nor_79_cse <= NOT((z_out_7(3)) OR (z_out_7(2)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse <= (z_out_7(4)) AND (z_out_7(1)) AND COMP_LOOP_tmp_nor_79_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
  COMP_LOOP_tmp_nor_32_cse <= NOT(CONV_SL_1_1(z_out_7(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse <= (z_out_7(4)) AND (z_out_7(1)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_27_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse <= (z_out_7(3)) AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_32_cse;
  COMP_LOOP_tmp_nor_81_cse <= NOT((z_out_7(3)) OR (z_out_7(1)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse <= (z_out_7(4)) AND (z_out_7(2)) AND COMP_LOOP_tmp_nor_81_cse;
  COMP_LOOP_tmp_nor_33_cse <= NOT((z_out_7(2)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse <= (z_out_7(3)) AND (z_out_7(1)) AND COMP_LOOP_tmp_nor_33_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse <= (z_out_7(4)) AND (z_out_7(2)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_29_cse;
  COMP_LOOP_tmp_nor_34_cse <= NOT(CONV_SL_1_1(z_out_7(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse <= (z_out_7(4)) AND (z_out_7(2)) AND (z_out_7(1))
      AND COMP_LOOP_tmp_nor_30_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_nor_34_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse <= (z_out_7(4)) AND (z_out_7(3)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_32_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse <= (z_out_7(4)) AND (z_out_7(3)) AND (z_out_7(1))
      AND COMP_LOOP_tmp_nor_33_cse;
  COMP_LOOP_tmp_or_12_cse <= and_dcpl_46 OR and_dcpl_49 OR and_dcpl_172 OR and_dcpl_173
      OR and_dcpl_176;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_tmp_nor_34_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
  COMP_LOOP_tmp_or_17_cse <= and_dcpl_46 OR and_dcpl_49 OR and_dcpl_172 OR and_dcpl_174;
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
  COMP_LOOP_or_42_cse <= and_dcpl_49 OR and_dcpl_172;
  COMP_LOOP_tmp_nor_1_cse <= NOT((z_out_7(4)) OR (z_out_7(3)) OR (z_out_7(2)) OR
      (z_out_7(0)));
  COMP_LOOP_or_41_cse <= and_dcpl_172 OR and_dcpl_173;
  COMP_LOOP_tmp_nor_101_cse <= NOT((z_out_7(4)) OR (z_out_7(3)) OR (z_out_7(1)) OR
      (z_out_7(0)));
  COMP_LOOP_tmp_nor_35_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
  COMP_LOOP_tmp_nor_105_cse <= NOT((z_out_7(4)) OR (z_out_7(2)) OR (z_out_7(1)) OR
      (z_out_7(0)));
  COMP_LOOP_or_39_cse <= and_dcpl_49 OR and_dcpl_172 OR and_dcpl_173;
  COMP_LOOP_or_36_itm <= and_dcpl_171 OR and_dcpl_222 OR and_dcpl_226 OR and_dcpl_229
      OR and_dcpl_232 OR and_dcpl_234 OR and_dcpl_236 OR and_dcpl_238;
  COMP_LOOP_tmp_or_35_cse <= and_dcpl_171 OR and_dcpl_174;
  COMP_LOOP_tmp_or_40_cse <= and_dcpl_173 OR and_dcpl_176;
  and_298_m1c <= and_dcpl_45 AND and_dcpl_175;
  and_1_cse <= (COMP_LOOP_2_tmp_mul_idiv_sva(0)) AND COMP_LOOP_tmp_nor_1_itm;
  nor_1025_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  and_456_cse <= ((fsm_output(3)) OR (fsm_output(6))) AND (fsm_output(7));
  mux_1588_nl <= MUX_s_1_2_2(mux_189_cse, and_464_cse, or_32_cse);
  mux_1589_nl <= MUX_s_1_2_2(mux_189_cse, mux_1588_nl, fsm_output(3));
  mux_1590_nl <= MUX_s_1_2_2(mux_1589_nl, and_464_cse, fsm_output(4));
  mux_1586_nl <= MUX_s_1_2_2(mux_189_cse, and_464_cse, fsm_output(3));
  mux_1587_nl <= MUX_s_1_2_2(mux_1586_nl, and_456_cse, fsm_output(4));
  mux_1591_nl <= MUX_s_1_2_2(mux_1590_nl, mux_1587_nl, fsm_output(2));
  mux_1592_tmp <= MUX_s_1_2_2(mux_1591_nl, (fsm_output(7)), fsm_output(5));
  and_490_cse <= (fsm_output(4)) AND (fsm_output(7));
  or_167_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  COMP_LOOP_1_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "000")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_1_acc_10_itm_10_1_1 <= COMP_LOOP_1_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_acc_psp_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
      DOWNTO 3)) + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0), 7));
  COMP_LOOP_acc_1_cse_6_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
      + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "101")), 10));
  COMP_LOOP_acc_1_cse_4_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
      + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "011")), 10));
  COMP_LOOP_acc_1_cse_2_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
      + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "001")), 10));
  COMP_LOOP_2_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "001")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_2_acc_10_itm_10_1_1 <= COMP_LOOP_2_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_3_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "010")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_3_acc_10_itm_10_1_1 <= COMP_LOOP_3_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_4_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "011")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_4_acc_10_itm_10_1_1 <= COMP_LOOP_4_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_5_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "100")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_5_acc_10_itm_10_1_1 <= COMP_LOOP_5_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_6_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "101")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_6_acc_10_itm_10_1_1 <= COMP_LOOP_6_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_7_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "110")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_7_acc_10_itm_10_1_1 <= COMP_LOOP_7_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_8_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "111")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_8_acc_10_itm_10_1_1 <= COMP_LOOP_8_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(1))
      AND COMP_LOOP_tmp_nor_49_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(2))
      AND COMP_LOOP_tmp_nor_1_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(3))
      AND COMP_LOOP_tmp_nor_14_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(4))
      AND COMP_LOOP_tmp_nor_3_itm;
  and_4_cse <= (COMP_LOOP_2_tmp_mul_idiv_sva(1)) AND COMP_LOOP_tmp_nor_14_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_119_rgt <= (COMP_LOOP_3_tmp_lshift_ncse_sva(1))
      AND COMP_LOOP_tmp_nor_26_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_121_rgt <= (COMP_LOOP_3_tmp_lshift_ncse_sva(2))
      AND COMP_LOOP_tmp_nor_28_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_125_rgt <= (COMP_LOOP_3_tmp_lshift_ncse_sva(3))
      AND COMP_LOOP_tmp_nor_31_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_165 <= (COMP_LOOP_2_tmp_mul_idiv_sva(4)) AND COMP_LOOP_tmp_nor_49_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 <= (COMP_LOOP_2_tmp_mul_idiv_sva(3)) AND COMP_LOOP_tmp_nor_42_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 <= (COMP_LOOP_2_tmp_mul_idiv_sva(2)) AND COMP_LOOP_tmp_nor_3_itm;
  nor_tmp_53 <= ((fsm_output(6)) OR (fsm_output(4))) AND (fsm_output(7));
  or_145_cse <= (fsm_output(4)) OR (fsm_output(7));
  and_485_cse <= (fsm_output(6)) AND (fsm_output(4));
  and_479_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"));
  or_tmp_142 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_28 <= NOT((fsm_output(2)) OR (fsm_output(5)));
  and_dcpl_29 <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_30 <= and_dcpl_29 AND and_dcpl_28;
  and_dcpl_31 <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_33 <= nor_1025_cse AND and_dcpl_31;
  and_dcpl_35 <= (fsm_output(2)) AND (fsm_output(5));
  and_dcpl_36 <= and_dcpl_29 AND and_dcpl_35;
  and_dcpl_38 <= and_464_cse AND and_dcpl_31;
  nor_tmp_95 <= ((fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1)))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_40 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_44 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_45 <= nor_1025_cse AND and_dcpl_44;
  and_dcpl_46 <= and_dcpl_45 AND and_dcpl_30;
  and_dcpl_48 <= nor_1025_cse AND and_316_cse;
  and_dcpl_49 <= and_dcpl_48 AND and_dcpl_30;
  and_dcpl_50 <= (fsm_output(2)) AND (NOT (fsm_output(5)));
  and_dcpl_52 <= and_479_cse AND and_dcpl_50;
  and_dcpl_54 <= and_dcpl_48 AND and_dcpl_52;
  and_dcpl_55 <= (NOT (fsm_output(2))) AND (fsm_output(5));
  and_dcpl_56 <= and_479_cse AND and_dcpl_55;
  and_dcpl_58 <= and_dcpl_48 AND and_dcpl_56;
  and_dcpl_59 <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_60 <= and_dcpl_59 AND and_dcpl_50;
  and_dcpl_61 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_62 <= and_dcpl_61 AND and_dcpl_44;
  and_dcpl_64 <= and_dcpl_61 AND and_316_cse;
  and_dcpl_65 <= and_dcpl_64 AND and_dcpl_60;
  and_dcpl_66 <= and_dcpl_59 AND and_dcpl_55;
  and_dcpl_68 <= and_dcpl_64 AND and_dcpl_66;
  and_dcpl_69 <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_70 <= and_dcpl_69 AND and_dcpl_50;
  and_dcpl_71 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_72 <= and_dcpl_71 AND and_dcpl_44;
  and_dcpl_74 <= and_dcpl_71 AND and_316_cse;
  and_dcpl_75 <= and_dcpl_74 AND and_dcpl_70;
  and_dcpl_76 <= and_dcpl_69 AND and_dcpl_55;
  and_dcpl_78 <= and_dcpl_74 AND and_dcpl_76;
  and_dcpl_79 <= and_dcpl_29 AND and_dcpl_50;
  and_dcpl_82 <= and_464_cse AND and_316_cse;
  and_dcpl_83 <= and_dcpl_82 AND and_dcpl_79;
  and_dcpl_85 <= nor_1025_cse AND and_dcpl_40;
  and_dcpl_89 <= and_dcpl_61 AND and_dcpl_31;
  and_dcpl_91 <= and_dcpl_61 AND and_dcpl_40;
  and_dcpl_95 <= and_dcpl_71 AND and_dcpl_31;
  and_dcpl_97 <= and_dcpl_71 AND and_dcpl_40;
  and_dcpl_102 <= and_464_cse AND and_dcpl_40;
  and_dcpl_104 <= and_dcpl_29 AND and_dcpl_55;
  or_238_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7)));
  or_236_nl <= (COMP_LOOP_acc_psp_sva(0)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR (COMP_LOOP_acc_psp_sva(1))
      OR (fsm_output(7));
  mux_322_cse <= MUX_s_1_2_2(or_238_nl, or_236_nl, fsm_output(4));
  or_284_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_282_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_311 <= MUX_s_1_2_2(or_284_nl, or_282_nl, fsm_output(4));
  nand_445_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(0)) AND (fsm_output(7)));
  nand_447_cse <= NOT((COMP_LOOP_acc_1_cse_6_sva(0)) AND (fsm_output(7)));
  nor_1001_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7))));
  nor_1002_nl <= NOT((COMP_LOOP_acc_psp_sva(0)) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR
      (COMP_LOOP_acc_psp_sva(1)) OR (fsm_output(7)));
  mux_353_cse <= MUX_s_1_2_2(nor_1001_nl, nor_1002_nl, fsm_output(4));
  nand_446_cse <= NOT((COMP_LOOP_acc_1_cse_sva(0)) AND (fsm_output(7)));
  nand_448_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_7_sva(0)) AND (fsm_output(7)));
  nor_98_cse <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")));
  nand_441_cse <= NOT((COMP_LOOP_acc_14_psp_sva(0)) AND (fsm_output(7)));
  nand_442_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(1)) AND (fsm_output(7)));
  or_388_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_386_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_373 <= MUX_s_1_2_2(or_388_nl, or_386_nl, fsm_output(4));
  nand_435_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7)));
  nand_437_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7)));
  or_446_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(7)));
  or_444_nl <= (COMP_LOOP_acc_psp_sva(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2))) OR
      (COMP_LOOP_acc_psp_sva(1)) OR (fsm_output(7));
  mux_446_cse <= MUX_s_1_2_2(or_446_nl, or_444_nl, fsm_output(4));
  or_492_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_490_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_435 <= MUX_s_1_2_2(or_492_nl, or_490_nl, fsm_output(4));
  nor_933_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(7))));
  nor_934_nl <= NOT((COMP_LOOP_acc_psp_sva(0)) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (COMP_LOOP_acc_psp_sva(1)) OR (fsm_output(7)));
  mux_477_cse <= MUX_s_1_2_2(nor_933_nl, nor_934_nl, fsm_output(4));
  nand_423_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7)));
  or_596_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_594_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_497 <= MUX_s_1_2_2(or_596_nl, or_594_nl, fsm_output(4));
  nand_417_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7)));
  nand_419_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7)));
  or_654_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(7)));
  or_652_nl <= (NOT (COMP_LOOP_acc_psp_sva(0))) OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR
      (COMP_LOOP_acc_psp_sva(1)) OR (fsm_output(7));
  mux_570_cse <= MUX_s_1_2_2(or_654_nl, or_652_nl, fsm_output(4));
  or_700_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_698_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_559 <= MUX_s_1_2_2(or_700_nl, or_698_nl, fsm_output(4));
  nand_411_cse <= NOT((COMP_LOOP_acc_1_cse_6_sva(3)) AND (COMP_LOOP_acc_1_cse_6_sva(0))
      AND (fsm_output(7)));
  nor_865_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(7))));
  nor_866_nl <= NOT((NOT (COMP_LOOP_acc_psp_sva(0))) OR (VEC_LOOP_j_10_0_sva_9_0(2))
      OR (COMP_LOOP_acc_psp_sva(1)) OR (fsm_output(7)));
  mux_601_cse <= MUX_s_1_2_2(nor_865_nl, nor_866_nl, fsm_output(4));
  or_804_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_802_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_621 <= MUX_s_1_2_2(or_804_nl, or_802_nl, fsm_output(4));
  nand_518_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(7)));
  or_860_nl <= (NOT (COMP_LOOP_acc_psp_sva(0))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (COMP_LOOP_acc_psp_sva(1)) OR (fsm_output(7));
  mux_694_cse <= MUX_s_1_2_2(nand_518_nl, or_860_nl, fsm_output(4));
  or_908_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_906_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_683 <= MUX_s_1_2_2(or_908_nl, or_906_nl, fsm_output(4));
  and_532_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(7));
  nor_798_nl <= NOT((NOT (COMP_LOOP_acc_psp_sva(0))) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(2)))
      OR (COMP_LOOP_acc_psp_sva(1)) OR (fsm_output(7)));
  mux_725_cse <= MUX_s_1_2_2(and_532_nl, nor_798_nl, fsm_output(4));
  nand_385_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7)));
  nand_472_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1009_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_745 <= MUX_s_1_2_2(nand_472_nl, or_1009_nl, fsm_output(4));
  nand_364_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_6_sva(4)) AND (fsm_output(7)));
  nand_365_cse <= NOT((COMP_LOOP_acc_13_psp_sva(2)) AND (fsm_output(7)));
  or_1112_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1110_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_807 <= MUX_s_1_2_2(or_1112_nl, or_1110_nl, fsm_output(4));
  nand_357_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_sva(0))
      AND (fsm_output(7)));
  nand_353_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(1))
      AND (fsm_output(7)));
  or_1216_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1214_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_869 <= MUX_s_1_2_2(or_1216_nl, or_1214_nl, fsm_output(4));
  or_1320_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1318_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_931 <= MUX_s_1_2_2(or_1320_nl, or_1318_nl, fsm_output(4));
  nand_469_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1422_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_993 <= MUX_s_1_2_2(nand_469_nl, or_1422_nl, fsm_output(4));
  nand_302_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7)));
  nand_303_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(7)));
  or_1527_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1525_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_1055 <= MUX_s_1_2_2(or_1527_nl, or_1525_nl, fsm_output(4));
  nand_294_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_sva(4))
      AND (COMP_LOOP_acc_10_cse_10_1_sva(0)) AND (fsm_output(7)));
  nand_297_cse <= NOT((COMP_LOOP_acc_1_cse_6_sva(4)) AND (COMP_LOOP_acc_1_cse_6_sva(3))
      AND (COMP_LOOP_acc_1_cse_6_sva(0)) AND (fsm_output(7)));
  nand_289_cse <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      AND (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) AND (fsm_output(7)));
  nand_466_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1627_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_1117 <= MUX_s_1_2_2(nand_466_nl, or_1627_nl, fsm_output(4));
  nand_266_cse <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7)));
  nand_268_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7)));
  nand_269_nl <= NOT((COMP_LOOP_acc_psp_sva(0)) AND (VEC_LOOP_j_10_0_sva_9_0(2))
      AND (COMP_LOOP_acc_psp_sva(1)) AND (NOT (fsm_output(7))));
  mux_1190_cse <= MUX_s_1_2_2(nand_268_nl, nand_269_nl, fsm_output(4));
  nand_463_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1727_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_1179 <= MUX_s_1_2_2(nand_463_nl, or_1727_nl, fsm_output(4));
  and_353_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7));
  and_354_nl <= (COMP_LOOP_acc_psp_sva(0)) AND (VEC_LOOP_j_10_0_sva_9_0(2)) AND (COMP_LOOP_acc_psp_sva(1))
      AND (NOT (fsm_output(7)));
  mux_1221_cse <= MUX_s_1_2_2(and_353_nl, and_354_nl, fsm_output(4));
  nand_459_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  nand_236_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("00")));
  mux_tmp_1241 <= MUX_s_1_2_2(nand_459_nl, nand_236_nl, fsm_output(4));
  and_dcpl_171 <= and_dcpl_33 AND and_dcpl_79;
  and_dcpl_172 <= and_dcpl_85 AND and_dcpl_79;
  and_dcpl_173 <= and_dcpl_45 AND and_dcpl_79;
  and_dcpl_174 <= and_dcpl_48 AND and_dcpl_79;
  and_dcpl_175 <= and_dcpl_69 AND and_dcpl_28;
  and_dcpl_176 <= and_dcpl_33 AND and_dcpl_175;
  and_dcpl_177 <= and_dcpl_85 AND and_dcpl_175;
  and_dcpl_178 <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_179 <= nor_1025_cse AND and_dcpl_178;
  not_tmp_617 <= NOT(CONV_SL_1_1(z_out_7(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      (fsm_output(1)));
  not_tmp_618 <= NOT((z_out_7(1)) AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")));
  not_tmp_625 <= NOT(CONV_SL_1_1(z_out_7(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND
      CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")));
  not_tmp_632 <= NOT((z_out_7(3)) AND (z_out_7(0)) AND (z_out_7(1)) AND (fsm_output(1)));
  mux_tmp_1423 <= MUX_s_1_2_2(or_167_cse, or_tmp_142, fsm_output(3));
  or_tmp_2024 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_1424 <= MUX_s_1_2_2((NOT and_464_cse), or_tmp_2024, fsm_output(3));
  or_tmp_2025 <= (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7));
  mux_tmp_1430 <= MUX_s_1_2_2(or_tmp_2024, or_167_cse, fsm_output(3));
  and_dcpl_220 <= and_dcpl_59 AND and_dcpl_28;
  and_dcpl_222 <= and_dcpl_33 AND and_dcpl_104;
  and_dcpl_223 <= and_dcpl_69 AND and_dcpl_35;
  and_dcpl_226 <= and_dcpl_33 AND and_479_cse AND and_dcpl_35;
  and_dcpl_229 <= and_dcpl_89 AND and_479_cse AND and_dcpl_28;
  and_dcpl_232 <= and_dcpl_89 AND and_dcpl_59 AND and_dcpl_35;
  and_dcpl_234 <= and_dcpl_95 AND and_dcpl_220;
  and_dcpl_236 <= and_dcpl_95 AND and_dcpl_223;
  and_dcpl_238 <= and_dcpl_38 AND and_dcpl_175;
  mux_240_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(4));
  mux_1470_nl <= MUX_s_1_2_2(and_490_cse, mux_240_nl, fsm_output(0));
  nand_tmp_184 <= NOT((fsm_output(3)) AND (NOT mux_1470_nl));
  or_2109_nl <= (fsm_output(0)) OR (NOT and_490_cse);
  mux_tmp_1437 <= MUX_s_1_2_2(or_145_cse, or_2109_nl, fsm_output(3));
  and_dcpl_244 <= (fsm_output(0)) AND (NOT (fsm_output(3)));
  or_dcpl_84 <= or_tmp_142 OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR or_212_cse OR (fsm_output(2)) OR (fsm_output(5));
  or_tmp_2048 <= and_316_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_1452 <= MUX_s_1_2_2((NOT or_tmp_2048), and_464_cse, or_212_cse);
  mux_1486_nl <= MUX_s_1_2_2(and_dcpl_82, and_464_cse, or_212_cse);
  mux_1488_nl <= MUX_s_1_2_2(mux_tmp_1452, mux_1486_nl, fsm_output(2));
  mux_1489_itm <= MUX_s_1_2_2(mux_1488_nl, and_464_cse, fsm_output(5));
  and_448_nl <= ((fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(6))) AND (fsm_output(7));
  mux_1490_nl <= MUX_s_1_2_2(and_464_cse, and_448_nl, fsm_output(3));
  mux_tmp_1456 <= MUX_s_1_2_2(mux_1490_nl, (fsm_output(7)), fsm_output(4));
  mux_1606_nl <= MUX_s_1_2_2(mux_189_cse, and_464_cse, and_316_cse);
  mux_tmp_1459 <= MUX_s_1_2_2(mux_1606_nl, and_464_cse, or_220_cse);
  and_tmp_11 <= (fsm_output(4)) AND ((fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(1)))
      AND (fsm_output(6));
  or_tmp_2054 <= and_316_cse OR (fsm_output(6));
  not_tmp_692 <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"))
      OR or_tmp_2054);
  or_tmp_2057 <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000")) OR
      and_316_cse;
  and_dcpl_252 <= or_tmp_2057 AND nor_1025_cse AND (NOT (fsm_output(5)));
  nor_340_nl <= NOT((fsm_output(3)) OR or_tmp_2054);
  and_511_nl <= (fsm_output(3)) AND (fsm_output(6));
  mux_tmp_1468 <= MUX_s_1_2_2(nor_340_nl, and_511_nl, fsm_output(4));
  and_tmp_13 <= (fsm_output(4)) AND ((fsm_output(3)) OR (fsm_output(1))) AND (fsm_output(6));
  nand_188_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")));
  mux_1510_nl <= MUX_s_1_2_2(or_tmp_2057, nand_188_nl, fsm_output(5));
  and_dcpl_256 <= mux_1510_nl AND nor_1025_cse;
  nor_tmp_324 <= (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(6));
  mux_1514_nl <= MUX_s_1_2_2(mux_tmp_1468, nor_tmp_324, fsm_output(2));
  mux_1515_nl <= MUX_s_1_2_2(mux_1514_nl, (fsm_output(6)), fsm_output(5));
  and_dcpl_259 <= NOT(mux_1515_nl OR (fsm_output(7)));
  mux_1599_nl <= MUX_s_1_2_2(mux_189_cse, and_464_cse, and_316_cse);
  mux_1516_nl <= MUX_s_1_2_2(mux_1599_nl, and_464_cse, fsm_output(3));
  mux_tmp_1482 <= MUX_s_1_2_2(mux_1516_nl, (fsm_output(7)), fsm_output(4));
  and_446_nl <= (and_496_cse OR (fsm_output(6))) AND (fsm_output(7));
  mux_tmp_1487 <= MUX_s_1_2_2(and_446_nl, (fsm_output(7)), fsm_output(4));
  mux_1525_nl <= MUX_s_1_2_2(nor_tmp_324, and_485_cse, fsm_output(2));
  mux_1526_nl <= MUX_s_1_2_2(not_tmp_692, mux_1525_nl, fsm_output(5));
  and_dcpl_260 <= NOT(mux_1526_nl OR (fsm_output(7)));
  mux_1530_nl <= MUX_s_1_2_2(mux_tmp_1482, nor_tmp_53, fsm_output(2));
  mux_1531_itm <= MUX_s_1_2_2(mux_1530_nl, (fsm_output(7)), fsm_output(5));
  and_306_nl <= ((fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(1))) AND CONV_SL_1_1(fsm_output(7
      DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  mux_1535_nl <= MUX_s_1_2_2(mux_tmp_1452, and_306_nl, fsm_output(2));
  mux_1536_itm <= MUX_s_1_2_2(mux_1535_nl, and_464_cse, fsm_output(5));
  mux_1537_nl <= MUX_s_1_2_2(nor_tmp_53, and_491_cse, fsm_output(2));
  mux_1538_itm <= MUX_s_1_2_2(mux_tmp_1459, mux_1537_nl, fsm_output(5));
  not_tmp_717 <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"))
      OR or_tmp_2048);
  mux_1542_nl <= MUX_s_1_2_2(mux_tmp_1452, and_33_cse, fsm_output(2));
  mux_1543_itm <= MUX_s_1_2_2(mux_1542_nl, and_464_cse, fsm_output(5));
  and_dcpl_262 <= nor_1023_cse AND (NOT (fsm_output(5)));
  and_dcpl_264 <= (NOT((NOT (fsm_output(1))) OR (fsm_output(6)) OR (fsm_output(7))))
      AND and_dcpl_244;
  nor_1128_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(1)));
  nor_1129_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(1))));
  mux_1551_nl <= MUX_s_1_2_2(nor_1128_nl, nor_1129_nl, fsm_output(2));
  and_dcpl_278 <= mux_1551_nl AND (NOT (fsm_output(7))) AND (NOT (fsm_output(6)))
      AND (fsm_output(0)) AND and_dcpl_178;
  or_tmp_2075 <= (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7));
  or_dcpl_109 <= or_tmp_142 OR (NOT and_316_cse) OR or_212_cse OR (NOT (fsm_output(2)))
      OR (fsm_output(5));
  STAGE_LOOP_i_3_0_sva_mx0c1 <= and_dcpl_38 AND and_dcpl_36;
  VEC_LOOP_j_10_0_sva_9_0_mx0c0 <= and_dcpl_85 AND and_dcpl_30;
  COMP_LOOP_tmp_mux1h_itm_mx0c0 <= and_dcpl_264 AND and_dcpl_262 AND CONV_SL_1_1(COMP_LOOP_1_tmp_mul_idiv_sva_1_0=STD_LOGIC_VECTOR'("00"));
  COMP_LOOP_tmp_mux1h_itm_mx0c1 <= and_dcpl_264 AND and_dcpl_262 AND CONV_SL_1_1(COMP_LOOP_1_tmp_mul_idiv_sva_1_0=STD_LOGIC_VECTOR'("01"));
  COMP_LOOP_tmp_mux1h_itm_mx0c2 <= and_dcpl_264 AND and_dcpl_262 AND CONV_SL_1_1(COMP_LOOP_1_tmp_mul_idiv_sva_1_0=STD_LOGIC_VECTOR'("10"));
  COMP_LOOP_tmp_mux1h_itm_mx0c3 <= and_dcpl_264 AND and_dcpl_262 AND CONV_SL_1_1(COMP_LOOP_1_tmp_mul_idiv_sva_1_0=STD_LOGIC_VECTOR'("11"));
  mux_1553_nl <= MUX_s_1_2_2(mux_tmp_1430, or_tmp_2075, fsm_output(4));
  nand_185_nl <= NOT((fsm_output(4)) AND (NOT mux_tmp_1424));
  mux_1554_nl <= MUX_s_1_2_2(mux_1553_nl, nand_185_nl, fsm_output(2));
  nand_473_nl <= NOT((fsm_output(4)) AND (fsm_output(3)) AND (NOT (fsm_output(6)))
      AND (fsm_output(7)));
  or_2171_nl <= (fsm_output(4)) OR mux_tmp_1423;
  mux_1552_nl <= MUX_s_1_2_2(nand_473_nl, or_2171_nl, fsm_output(2));
  mux_1555_nl <= MUX_s_1_2_2(mux_1554_nl, mux_1552_nl, fsm_output(5));
  COMP_LOOP_1_acc_8_itm_mx0c4 <= (NOT mux_1555_nl) AND and_dcpl_40;
  or_229_nl <= or_32_cse OR or_212_cse;
  mux_1574_nl <= MUX_s_1_2_2(or_212_cse, or_229_nl, fsm_output(2));
  mux_1573_nl <= MUX_s_1_2_2((fsm_output(4)), or_212_cse, fsm_output(2));
  mux_1575_nl <= MUX_s_1_2_2(mux_1574_nl, (NOT mux_1573_nl), fsm_output(5));
  and_294_tmp <= mux_1575_nl AND nor_1025_cse;
  mux_1577_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), or_212_cse);
  nor_1059_nl <= NOT((fsm_output(1)) OR (fsm_output(6)));
  mux_1576_nl <= MUX_s_1_2_2(nor_1059_nl, (fsm_output(6)), or_212_cse);
  mux_1578_nl <= MUX_s_1_2_2(mux_1577_nl, mux_1576_nl, fsm_output(2));
  mux_1579_nl <= MUX_s_1_2_2(mux_1578_nl, (fsm_output(6)), fsm_output(5));
  nor_1119_tmp <= NOT(mux_1579_nl OR (fsm_output(7)));
  nor_1062_nl <= NOT((fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(6)));
  nor_1063_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR or_tmp_2054);
  mux_1580_nl <= MUX_s_1_2_2(nor_1062_nl, nor_1063_nl, fsm_output(2));
  and_520_nl <= or_220_cse AND (fsm_output(6));
  mux_1581_nl <= MUX_s_1_2_2(mux_1580_nl, and_520_nl, fsm_output(5));
  nor_tmp <= NOT(mux_1581_nl OR (fsm_output(7)));
  nor_1117_tmp <= NOT((NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 3)/=STD_LOGIC_VECTOR'("0000"))))
      OR (fsm_output(7)));
  and_54_nl <= ((fsm_output(6)) XOR (fsm_output(3))) AND ((fsm_output(7)) XOR (fsm_output(4)))
      AND and_dcpl_40 AND ((fsm_output(2)) XOR (fsm_output(5)));
  vec_rsc_0_0_i_d_d_pff <= MUX_v_64_2_2(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z,
      COMP_LOOP_1_acc_8_itm, and_54_nl);
  and_64_nl <= and_dcpl_45 AND and_dcpl_52;
  and_68_nl <= and_dcpl_45 AND and_dcpl_56;
  and_74_nl <= and_dcpl_62 AND and_dcpl_60;
  and_78_nl <= and_dcpl_62 AND and_dcpl_66;
  and_84_nl <= and_dcpl_72 AND and_dcpl_70;
  and_88_nl <= and_dcpl_72 AND and_dcpl_76;
  and_92_nl <= and_464_cse AND and_dcpl_44 AND and_dcpl_79;
  vec_rsc_0_0_i_radr_d_pff <= MUX1HOT_v_5_16_2((COMP_LOOP_1_acc_10_itm_10_1_1(9 DOWNTO
      5)), (COMP_LOOP_acc_psp_sva(6 DOWNTO 2)), (COMP_LOOP_acc_1_cse_2_sva(9 DOWNTO
      5)), (COMP_LOOP_acc_10_cse_10_1_2_sva(9 DOWNTO 5)), (COMP_LOOP_acc_11_psp_sva(8
      DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_3_sva(9 DOWNTO 5)), (COMP_LOOP_acc_1_cse_4_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_4_sva(9 DOWNTO 5)), (COMP_LOOP_acc_13_psp_sva(7
      DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_5_sva(9 DOWNTO 5)), (COMP_LOOP_acc_1_cse_6_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_6_sva(9 DOWNTO 5)), (COMP_LOOP_acc_14_psp_sva(8
      DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_7_sva(9 DOWNTO 5)), (COMP_LOOP_acc_1_cse_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_sva(9 DOWNTO 5)), STD_LOGIC_VECTOR'(
      and_dcpl_46 & and_dcpl_49 & and_64_nl & and_dcpl_54 & and_68_nl & and_dcpl_58
      & and_74_nl & and_dcpl_65 & and_78_nl & and_dcpl_68 & and_84_nl & and_dcpl_75
      & and_88_nl & and_dcpl_78 & and_92_nl & and_dcpl_83));
  and_95_nl <= and_dcpl_33 AND and_dcpl_52;
  and_97_nl <= and_dcpl_85 AND and_dcpl_52;
  and_98_nl <= and_dcpl_33 AND and_dcpl_56;
  and_99_nl <= and_dcpl_85 AND and_dcpl_56;
  and_101_nl <= and_dcpl_89 AND and_dcpl_60;
  and_103_nl <= and_dcpl_91 AND and_dcpl_60;
  and_104_nl <= and_dcpl_89 AND and_dcpl_66;
  and_105_nl <= and_dcpl_91 AND and_dcpl_66;
  and_107_nl <= and_dcpl_95 AND and_dcpl_70;
  and_109_nl <= and_dcpl_97 AND and_dcpl_70;
  and_110_nl <= and_dcpl_95 AND and_dcpl_76;
  and_111_nl <= and_dcpl_97 AND and_dcpl_76;
  and_112_nl <= and_dcpl_38 AND and_dcpl_79;
  and_114_nl <= and_dcpl_102 AND and_dcpl_79;
  and_116_nl <= and_dcpl_38 AND and_dcpl_104;
  and_117_nl <= and_dcpl_102 AND and_dcpl_104;
  vec_rsc_0_0_i_wadr_d_pff <= MUX1HOT_v_5_16_2((COMP_LOOP_acc_10_cse_10_1_1_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_psp_sva(6 DOWNTO 2)), (COMP_LOOP_acc_10_cse_10_1_2_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_1_cse_2_sva(9 DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_3_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_11_psp_sva(8 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_4_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_1_cse_4_sva(9 DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_5_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_13_psp_sva(7 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_6_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_1_cse_6_sva(9 DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_7_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_14_psp_sva(8 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_sva(9
      DOWNTO 5)), (COMP_LOOP_acc_1_cse_sva(9 DOWNTO 5)), STD_LOGIC_VECTOR'( and_95_nl
      & and_97_nl & and_98_nl & and_99_nl & and_101_nl & and_103_nl & and_104_nl
      & and_105_nl & and_107_nl & and_109_nl & and_110_nl & and_111_nl & and_112_nl
      & and_114_nl & and_116_nl & and_117_nl));
  nor_1010_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(7))));
  nor_1011_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(7)));
  mux_333_nl <= MUX_s_1_2_2(nor_1010_nl, nor_1011_nl, fsm_output(4));
  nor_1012_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(7))));
  nor_1013_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(7)));
  mux_332_nl <= MUX_s_1_2_2(nor_1012_nl, nor_1013_nl, fsm_output(4));
  mux_334_nl <= MUX_s_1_2_2(mux_333_nl, mux_332_nl, fsm_output(0));
  and_443_nl <= (fsm_output(6)) AND mux_334_nl;
  or_257_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(7)));
  or_255_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(7));
  mux_330_nl <= MUX_s_1_2_2(or_257_nl, or_255_nl, fsm_output(4));
  or_254_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(7)));
  or_252_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(7));
  mux_329_nl <= MUX_s_1_2_2(or_254_nl, or_252_nl, fsm_output(4));
  mux_331_nl <= MUX_s_1_2_2(mux_330_nl, mux_329_nl, fsm_output(0));
  nor_1014_nl <= NOT((fsm_output(6)) OR mux_331_nl);
  mux_335_nl <= MUX_s_1_2_2(and_443_nl, nor_1014_nl, fsm_output(3));
  nand_506_nl <= NOT((fsm_output(5)) AND mux_335_nl);
  nor_1016_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(7))));
  nor_1017_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(7)));
  mux_326_nl <= MUX_s_1_2_2(nor_1016_nl, nor_1017_nl, fsm_output(4));
  or_246_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7)));
  or_244_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7));
  mux_325_nl <= MUX_s_1_2_2(or_246_nl, or_244_nl, fsm_output(4));
  nor_1018_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_325_nl);
  mux_327_nl <= MUX_s_1_2_2(mux_326_nl, nor_1018_nl, fsm_output(0));
  nand_8_nl <= NOT((fsm_output(6)) AND mux_327_nl);
  or_242_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(7)));
  or_240_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(7));
  mux_323_nl <= MUX_s_1_2_2(or_242_nl, or_240_nl, fsm_output(4));
  or_239_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR mux_322_cse;
  mux_324_nl <= MUX_s_1_2_2(mux_323_nl, or_239_nl, fsm_output(0));
  or_243_nl <= (fsm_output(6)) OR mux_324_nl;
  mux_328_nl <= MUX_s_1_2_2(nand_8_nl, or_243_nl, fsm_output(3));
  or_2280_nl <= (fsm_output(5)) OR mux_328_nl;
  mux_336_nl <= MUX_s_1_2_2(nand_506_nl, or_2280_nl, fsm_output(2));
  vec_rsc_0_0_i_we_d_pff <= NOT(mux_336_nl OR (fsm_output(1)));
  nor_1003_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_1004_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_350_nl <= MUX_s_1_2_2(nor_1003_nl, nor_1004_nl, fsm_output(0));
  nor_1005_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_348_cse);
  nor_1006_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_1007_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_1008_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_344_nl <= MUX_s_1_2_2(nor_1007_nl, nor_1008_nl, fsm_output(4));
  mux_345_nl <= MUX_s_1_2_2(nor_1006_nl, mux_344_nl, fsm_output(3));
  mux_349_nl <= MUX_s_1_2_2(nor_1005_nl, mux_345_nl, fsm_output(0));
  mux_351_nl <= MUX_s_1_2_2(mux_350_nl, mux_349_nl, fsm_output(5));
  or_276_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_274_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_341_nl <= MUX_s_1_2_2(or_276_nl, or_274_nl, fsm_output(4));
  or_273_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_271_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_340_nl <= MUX_s_1_2_2(or_273_nl, or_271_nl, fsm_output(4));
  mux_342_nl <= MUX_s_1_2_2(mux_341_nl, mux_340_nl, fsm_output(3));
  or_270_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR nand_443_cse;
  or_268_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_338_nl <= MUX_s_1_2_2(or_270_nl, or_268_nl, fsm_output(4));
  or_267_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_265_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_337_nl <= MUX_s_1_2_2(or_267_nl, or_265_nl, fsm_output(4));
  mux_339_nl <= MUX_s_1_2_2(mux_338_nl, mux_337_nl, fsm_output(3));
  mux_343_nl <= MUX_s_1_2_2(mux_342_nl, mux_339_nl, fsm_output(0));
  nor_1009_nl <= NOT((fsm_output(5)) OR mux_343_nl);
  mux_352_nl <= MUX_s_1_2_2(mux_351_nl, nor_1009_nl, fsm_output(2));
  vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_352_nl AND (fsm_output(1));
  nor_991_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_445_cse);
  nor_992_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (fsm_output(7)));
  mux_364_nl <= MUX_s_1_2_2(nor_991_nl, nor_992_nl, fsm_output(4));
  nor_993_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_446_cse);
  nor_994_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (fsm_output(7)));
  mux_363_nl <= MUX_s_1_2_2(nor_993_nl, nor_994_nl, fsm_output(4));
  mux_365_nl <= MUX_s_1_2_2(mux_364_nl, mux_363_nl, fsm_output(0));
  and_440_nl <= (fsm_output(6)) AND mux_365_nl;
  or_308_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT (fsm_output(7)));
  or_306_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (fsm_output(7));
  mux_361_nl <= MUX_s_1_2_2(or_308_nl, or_306_nl, fsm_output(4));
  or_305_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_447_cse;
  or_303_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (fsm_output(7));
  mux_360_nl <= MUX_s_1_2_2(or_305_nl, or_303_nl, fsm_output(4));
  mux_362_nl <= MUX_s_1_2_2(mux_361_nl, mux_360_nl, fsm_output(0));
  nor_995_nl <= NOT((fsm_output(6)) OR mux_362_nl);
  mux_366_nl <= MUX_s_1_2_2(and_440_nl, nor_995_nl, fsm_output(3));
  nand_505_nl <= NOT((fsm_output(5)) AND mux_366_nl);
  nor_997_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_448_cse);
  nor_998_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (fsm_output(7)));
  mux_357_nl <= MUX_s_1_2_2(nor_997_nl, nor_998_nl, fsm_output(4));
  nor_999_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(7))));
  nor_1000_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(7)));
  mux_356_nl <= MUX_s_1_2_2(nor_999_nl, nor_1000_nl, fsm_output(4));
  and_441_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_356_nl;
  mux_358_nl <= MUX_s_1_2_2(mux_357_nl, and_441_nl, fsm_output(0));
  nand_14_nl <= NOT((fsm_output(6)) AND mux_358_nl);
  or_294_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT (fsm_output(7)));
  or_292_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (fsm_output(7));
  mux_354_nl <= MUX_s_1_2_2(or_294_nl, or_292_nl, fsm_output(4));
  nand_12_nl <= NOT(nor_98_cse AND mux_353_cse);
  mux_355_nl <= MUX_s_1_2_2(mux_354_nl, nand_12_nl, fsm_output(0));
  or_295_nl <= (fsm_output(6)) OR mux_355_nl;
  mux_359_nl <= MUX_s_1_2_2(nand_14_nl, or_295_nl, fsm_output(3));
  or_2279_nl <= (fsm_output(5)) OR mux_359_nl;
  mux_367_nl <= MUX_s_1_2_2(nand_505_nl, or_2279_nl, fsm_output(2));
  vec_rsc_0_1_i_we_d_pff <= NOT(mux_367_nl OR (fsm_output(1)));
  nor_985_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_986_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_381_nl <= MUX_s_1_2_2(nor_985_nl, nor_986_nl, fsm_output(0));
  and_438_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_348_cse);
  nor_987_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_988_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_989_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_375_nl <= MUX_s_1_2_2(nor_988_nl, nor_989_nl, fsm_output(4));
  mux_376_nl <= MUX_s_1_2_2(nor_987_nl, mux_375_nl, fsm_output(3));
  mux_380_nl <= MUX_s_1_2_2(and_438_nl, mux_376_nl, fsm_output(0));
  mux_382_nl <= MUX_s_1_2_2(mux_381_nl, mux_380_nl, fsm_output(5));
  or_327_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_325_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_372_nl <= MUX_s_1_2_2(or_327_nl, or_325_nl, fsm_output(4));
  or_324_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_322_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_371_nl <= MUX_s_1_2_2(or_324_nl, or_322_nl, fsm_output(4));
  mux_373_nl <= MUX_s_1_2_2(mux_372_nl, mux_371_nl, fsm_output(3));
  or_321_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_444_cse;
  or_319_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_369_nl <= MUX_s_1_2_2(or_321_nl, or_319_nl, fsm_output(4));
  or_318_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_316_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_368_nl <= MUX_s_1_2_2(or_318_nl, or_316_nl, fsm_output(4));
  mux_370_nl <= MUX_s_1_2_2(mux_369_nl, mux_368_nl, fsm_output(3));
  mux_374_nl <= MUX_s_1_2_2(mux_373_nl, mux_370_nl, fsm_output(0));
  nor_990_nl <= NOT((fsm_output(5)) OR mux_374_nl);
  mux_383_nl <= MUX_s_1_2_2(mux_382_nl, nor_990_nl, fsm_output(2));
  vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_383_nl AND (fsm_output(1));
  nor_976_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(7))));
  nor_977_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(7)));
  mux_395_nl <= MUX_s_1_2_2(nor_976_nl, nor_977_nl, fsm_output(4));
  nor_978_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(7))));
  nor_979_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(7)));
  mux_394_nl <= MUX_s_1_2_2(nor_978_nl, nor_979_nl, fsm_output(4));
  mux_396_nl <= MUX_s_1_2_2(mux_395_nl, mux_394_nl, fsm_output(0));
  and_437_nl <= (fsm_output(6)) AND mux_396_nl;
  or_361_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(7)));
  or_359_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(7));
  mux_392_nl <= MUX_s_1_2_2(or_361_nl, or_359_nl, fsm_output(4));
  or_358_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(7)));
  or_356_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(7));
  mux_391_nl <= MUX_s_1_2_2(or_358_nl, or_356_nl, fsm_output(4));
  mux_393_nl <= MUX_s_1_2_2(mux_392_nl, mux_391_nl, fsm_output(0));
  nor_980_nl <= NOT((fsm_output(6)) OR mux_393_nl);
  mux_397_nl <= MUX_s_1_2_2(and_437_nl, nor_980_nl, fsm_output(3));
  nand_504_nl <= NOT((fsm_output(5)) AND mux_397_nl);
  nor_982_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(7))));
  nor_983_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(7)));
  mux_388_nl <= MUX_s_1_2_2(nor_982_nl, nor_983_nl, fsm_output(4));
  or_350_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))
      OR nand_441_cse;
  or_348_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7));
  mux_387_nl <= MUX_s_1_2_2(or_350_nl, or_348_nl, fsm_output(4));
  nor_984_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_387_nl);
  mux_389_nl <= MUX_s_1_2_2(mux_388_nl, nor_984_nl, fsm_output(0));
  nand_19_nl <= NOT((fsm_output(6)) AND mux_389_nl);
  or_346_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      OR nand_442_cse;
  or_344_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(7));
  mux_385_nl <= MUX_s_1_2_2(or_346_nl, or_344_nl, fsm_output(4));
  or_343_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR mux_322_cse;
  mux_386_nl <= MUX_s_1_2_2(mux_385_nl, or_343_nl, fsm_output(0));
  or_347_nl <= (fsm_output(6)) OR mux_386_nl;
  mux_390_nl <= MUX_s_1_2_2(nand_19_nl, or_347_nl, fsm_output(3));
  or_2278_nl <= (fsm_output(5)) OR mux_390_nl;
  mux_398_nl <= MUX_s_1_2_2(nand_504_nl, or_2278_nl, fsm_output(2));
  vec_rsc_0_2_i_we_d_pff <= NOT(mux_398_nl OR (fsm_output(1)));
  nor_969_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_970_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_412_nl <= MUX_s_1_2_2(nor_969_nl, nor_970_nl, fsm_output(0));
  nor_971_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_410_cse);
  nor_972_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_973_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_974_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_406_nl <= MUX_s_1_2_2(nor_973_nl, nor_974_nl, fsm_output(4));
  mux_407_nl <= MUX_s_1_2_2(nor_972_nl, mux_406_nl, fsm_output(3));
  mux_411_nl <= MUX_s_1_2_2(nor_971_nl, mux_407_nl, fsm_output(0));
  mux_413_nl <= MUX_s_1_2_2(mux_412_nl, mux_411_nl, fsm_output(5));
  or_380_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_378_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_403_nl <= MUX_s_1_2_2(or_380_nl, or_378_nl, fsm_output(4));
  or_377_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_375_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_402_nl <= MUX_s_1_2_2(or_377_nl, or_375_nl, fsm_output(4));
  mux_404_nl <= MUX_s_1_2_2(mux_403_nl, mux_402_nl, fsm_output(3));
  or_374_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR nand_443_cse;
  or_372_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_400_nl <= MUX_s_1_2_2(or_374_nl, or_372_nl, fsm_output(4));
  or_371_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_369_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_399_nl <= MUX_s_1_2_2(or_371_nl, or_369_nl, fsm_output(4));
  mux_401_nl <= MUX_s_1_2_2(mux_400_nl, mux_399_nl, fsm_output(3));
  mux_405_nl <= MUX_s_1_2_2(mux_404_nl, mux_401_nl, fsm_output(0));
  nor_975_nl <= NOT((fsm_output(5)) OR mux_405_nl);
  mux_414_nl <= MUX_s_1_2_2(mux_413_nl, nor_975_nl, fsm_output(2));
  vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_414_nl AND (fsm_output(1));
  nor_957_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR nand_445_cse);
  nor_958_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (fsm_output(7)));
  mux_426_nl <= MUX_s_1_2_2(nor_957_nl, nor_958_nl, fsm_output(4));
  nor_959_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"))
      OR nand_435_cse);
  nor_960_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (fsm_output(7)));
  mux_425_nl <= MUX_s_1_2_2(nor_959_nl, nor_960_nl, fsm_output(4));
  mux_427_nl <= MUX_s_1_2_2(mux_426_nl, mux_425_nl, fsm_output(0));
  and_434_nl <= (fsm_output(6)) AND mux_427_nl;
  or_412_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT (fsm_output(7)));
  or_410_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (fsm_output(7));
  mux_423_nl <= MUX_s_1_2_2(or_412_nl, or_410_nl, fsm_output(4));
  or_409_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR nand_447_cse;
  or_407_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (fsm_output(7));
  mux_422_nl <= MUX_s_1_2_2(or_409_nl, or_407_nl, fsm_output(4));
  mux_424_nl <= MUX_s_1_2_2(mux_423_nl, mux_422_nl, fsm_output(0));
  nor_961_nl <= NOT((fsm_output(6)) OR mux_424_nl);
  mux_428_nl <= MUX_s_1_2_2(and_434_nl, nor_961_nl, fsm_output(3));
  nand_503_nl <= NOT((fsm_output(5)) AND mux_428_nl);
  nor_963_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"))
      OR nand_437_cse);
  nor_964_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (fsm_output(7)));
  mux_419_nl <= MUX_s_1_2_2(nor_963_nl, nor_964_nl, fsm_output(4));
  nor_965_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))
      OR nand_441_cse);
  nor_966_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(7)));
  mux_418_nl <= MUX_s_1_2_2(nor_965_nl, nor_966_nl, fsm_output(4));
  and_435_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_418_nl;
  mux_420_nl <= MUX_s_1_2_2(mux_419_nl, and_435_nl, fsm_output(0));
  nand_25_nl <= NOT((fsm_output(6)) AND mux_420_nl);
  or_398_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      OR nand_442_cse;
  or_396_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (fsm_output(7));
  mux_416_nl <= MUX_s_1_2_2(or_398_nl, or_396_nl, fsm_output(4));
  nand_23_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_353_cse);
  mux_417_nl <= MUX_s_1_2_2(mux_416_nl, nand_23_nl, fsm_output(0));
  or_399_nl <= (fsm_output(6)) OR mux_417_nl;
  mux_421_nl <= MUX_s_1_2_2(nand_25_nl, or_399_nl, fsm_output(3));
  or_2277_nl <= (fsm_output(5)) OR mux_421_nl;
  mux_429_nl <= MUX_s_1_2_2(nand_503_nl, or_2277_nl, fsm_output(2));
  vec_rsc_0_3_i_we_d_pff <= NOT(mux_429_nl OR (fsm_output(1)));
  nor_951_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_952_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_443_nl <= MUX_s_1_2_2(nor_951_nl, nor_952_nl, fsm_output(0));
  and_432_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_410_cse);
  nor_953_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_954_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_955_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_437_nl <= MUX_s_1_2_2(nor_954_nl, nor_955_nl, fsm_output(4));
  mux_438_nl <= MUX_s_1_2_2(nor_953_nl, mux_437_nl, fsm_output(3));
  mux_442_nl <= MUX_s_1_2_2(and_432_nl, mux_438_nl, fsm_output(0));
  mux_444_nl <= MUX_s_1_2_2(mux_443_nl, mux_442_nl, fsm_output(5));
  or_431_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_429_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_434_nl <= MUX_s_1_2_2(or_431_nl, or_429_nl, fsm_output(4));
  or_428_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_426_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_433_nl <= MUX_s_1_2_2(or_428_nl, or_426_nl, fsm_output(4));
  mux_435_nl <= MUX_s_1_2_2(mux_434_nl, mux_433_nl, fsm_output(3));
  or_425_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR nand_444_cse;
  or_423_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_431_nl <= MUX_s_1_2_2(or_425_nl, or_423_nl, fsm_output(4));
  or_422_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_420_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_430_nl <= MUX_s_1_2_2(or_422_nl, or_420_nl, fsm_output(4));
  mux_432_nl <= MUX_s_1_2_2(mux_431_nl, mux_430_nl, fsm_output(3));
  mux_436_nl <= MUX_s_1_2_2(mux_435_nl, mux_432_nl, fsm_output(0));
  nor_956_nl <= NOT((fsm_output(5)) OR mux_436_nl);
  mux_445_nl <= MUX_s_1_2_2(mux_444_nl, nor_956_nl, fsm_output(2));
  vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_445_nl AND (fsm_output(1));
  nor_942_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(7))));
  nor_943_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(7)));
  mux_457_nl <= MUX_s_1_2_2(nor_942_nl, nor_943_nl, fsm_output(4));
  nor_944_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(7))));
  nor_945_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(7)));
  mux_456_nl <= MUX_s_1_2_2(nor_944_nl, nor_945_nl, fsm_output(4));
  mux_458_nl <= MUX_s_1_2_2(mux_457_nl, mux_456_nl, fsm_output(0));
  and_431_nl <= (fsm_output(6)) AND mux_458_nl;
  or_465_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(7)));
  or_463_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(7));
  mux_454_nl <= MUX_s_1_2_2(or_465_nl, or_463_nl, fsm_output(4));
  or_462_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(7)));
  or_460_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(7));
  mux_453_nl <= MUX_s_1_2_2(or_462_nl, or_460_nl, fsm_output(4));
  mux_455_nl <= MUX_s_1_2_2(mux_454_nl, mux_453_nl, fsm_output(0));
  nor_946_nl <= NOT((fsm_output(6)) OR mux_455_nl);
  mux_459_nl <= MUX_s_1_2_2(and_431_nl, nor_946_nl, fsm_output(3));
  nand_502_nl <= NOT((fsm_output(5)) AND mux_459_nl);
  nor_948_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(7))));
  nor_949_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(7)));
  mux_450_nl <= MUX_s_1_2_2(nor_948_nl, nor_949_nl, fsm_output(4));
  or_454_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7)));
  or_452_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7));
  mux_449_nl <= MUX_s_1_2_2(or_454_nl, or_452_nl, fsm_output(4));
  nor_950_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_449_nl);
  mux_451_nl <= MUX_s_1_2_2(mux_450_nl, nor_950_nl, fsm_output(0));
  nand_30_nl <= NOT((fsm_output(6)) AND mux_451_nl);
  or_450_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(7)));
  or_448_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(7));
  mux_447_nl <= MUX_s_1_2_2(or_450_nl, or_448_nl, fsm_output(4));
  or_447_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR mux_446_cse;
  mux_448_nl <= MUX_s_1_2_2(mux_447_nl, or_447_nl, fsm_output(0));
  or_451_nl <= (fsm_output(6)) OR mux_448_nl;
  mux_452_nl <= MUX_s_1_2_2(nand_30_nl, or_451_nl, fsm_output(3));
  or_2276_nl <= (fsm_output(5)) OR mux_452_nl;
  mux_460_nl <= MUX_s_1_2_2(nand_502_nl, or_2276_nl, fsm_output(2));
  vec_rsc_0_4_i_we_d_pff <= NOT(mux_460_nl OR (fsm_output(1)));
  nor_935_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_936_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_474_nl <= MUX_s_1_2_2(nor_935_nl, nor_936_nl, fsm_output(0));
  nor_937_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_472_cse);
  nor_938_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_939_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_940_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_468_nl <= MUX_s_1_2_2(nor_939_nl, nor_940_nl, fsm_output(4));
  mux_469_nl <= MUX_s_1_2_2(nor_938_nl, mux_468_nl, fsm_output(3));
  mux_473_nl <= MUX_s_1_2_2(nor_937_nl, mux_469_nl, fsm_output(0));
  mux_475_nl <= MUX_s_1_2_2(mux_474_nl, mux_473_nl, fsm_output(5));
  or_484_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_482_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_465_nl <= MUX_s_1_2_2(or_484_nl, or_482_nl, fsm_output(4));
  or_481_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_479_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_464_nl <= MUX_s_1_2_2(or_481_nl, or_479_nl, fsm_output(4));
  mux_466_nl <= MUX_s_1_2_2(mux_465_nl, mux_464_nl, fsm_output(3));
  or_478_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR nand_443_cse;
  or_476_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_462_nl <= MUX_s_1_2_2(or_478_nl, or_476_nl, fsm_output(4));
  or_475_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_473_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_461_nl <= MUX_s_1_2_2(or_475_nl, or_473_nl, fsm_output(4));
  mux_463_nl <= MUX_s_1_2_2(mux_462_nl, mux_461_nl, fsm_output(3));
  mux_467_nl <= MUX_s_1_2_2(mux_466_nl, mux_463_nl, fsm_output(0));
  nor_941_nl <= NOT((fsm_output(5)) OR mux_467_nl);
  mux_476_nl <= MUX_s_1_2_2(mux_475_nl, nor_941_nl, fsm_output(2));
  vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_476_nl AND (fsm_output(1));
  nor_923_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_445_cse);
  nor_924_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (fsm_output(7)));
  mux_488_nl <= MUX_s_1_2_2(nor_923_nl, nor_924_nl, fsm_output(4));
  nor_925_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_446_cse);
  nor_926_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (fsm_output(7)));
  mux_487_nl <= MUX_s_1_2_2(nor_925_nl, nor_926_nl, fsm_output(4));
  mux_489_nl <= MUX_s_1_2_2(mux_488_nl, mux_487_nl, fsm_output(0));
  and_428_nl <= (fsm_output(6)) AND mux_489_nl;
  or_516_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT (fsm_output(7)));
  or_514_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (fsm_output(7));
  mux_485_nl <= MUX_s_1_2_2(or_516_nl, or_514_nl, fsm_output(4));
  or_513_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_447_cse;
  or_511_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (fsm_output(7));
  mux_484_nl <= MUX_s_1_2_2(or_513_nl, or_511_nl, fsm_output(4));
  mux_486_nl <= MUX_s_1_2_2(mux_485_nl, mux_484_nl, fsm_output(0));
  nor_927_nl <= NOT((fsm_output(6)) OR mux_486_nl);
  mux_490_nl <= MUX_s_1_2_2(and_428_nl, nor_927_nl, fsm_output(3));
  nand_501_nl <= NOT((fsm_output(5)) AND mux_490_nl);
  nor_929_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_448_cse);
  nor_930_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (fsm_output(7)));
  mux_481_nl <= MUX_s_1_2_2(nor_929_nl, nor_930_nl, fsm_output(4));
  nor_931_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(7))));
  nor_932_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(7)));
  mux_480_nl <= MUX_s_1_2_2(nor_931_nl, nor_932_nl, fsm_output(4));
  and_429_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_480_nl;
  mux_482_nl <= MUX_s_1_2_2(mux_481_nl, and_429_nl, fsm_output(0));
  nand_36_nl <= NOT((fsm_output(6)) AND mux_482_nl);
  or_502_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT (fsm_output(7)));
  or_500_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (fsm_output(7));
  mux_478_nl <= MUX_s_1_2_2(or_502_nl, or_500_nl, fsm_output(4));
  nand_34_nl <= NOT(nor_98_cse AND mux_477_cse);
  mux_479_nl <= MUX_s_1_2_2(mux_478_nl, nand_34_nl, fsm_output(0));
  or_503_nl <= (fsm_output(6)) OR mux_479_nl;
  mux_483_nl <= MUX_s_1_2_2(nand_36_nl, or_503_nl, fsm_output(3));
  or_2275_nl <= (fsm_output(5)) OR mux_483_nl;
  mux_491_nl <= MUX_s_1_2_2(nand_501_nl, or_2275_nl, fsm_output(2));
  vec_rsc_0_5_i_we_d_pff <= NOT(mux_491_nl OR (fsm_output(1)));
  nor_917_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_918_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_505_nl <= MUX_s_1_2_2(nor_917_nl, nor_918_nl, fsm_output(0));
  and_426_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_472_cse);
  nor_919_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_920_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_921_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_499_nl <= MUX_s_1_2_2(nor_920_nl, nor_921_nl, fsm_output(4));
  mux_500_nl <= MUX_s_1_2_2(nor_919_nl, mux_499_nl, fsm_output(3));
  mux_504_nl <= MUX_s_1_2_2(and_426_nl, mux_500_nl, fsm_output(0));
  mux_506_nl <= MUX_s_1_2_2(mux_505_nl, mux_504_nl, fsm_output(5));
  or_535_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_533_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_496_nl <= MUX_s_1_2_2(or_535_nl, or_533_nl, fsm_output(4));
  or_532_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_530_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_495_nl <= MUX_s_1_2_2(or_532_nl, or_530_nl, fsm_output(4));
  mux_497_nl <= MUX_s_1_2_2(mux_496_nl, mux_495_nl, fsm_output(3));
  or_529_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_444_cse;
  or_527_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_493_nl <= MUX_s_1_2_2(or_529_nl, or_527_nl, fsm_output(4));
  or_526_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_524_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_492_nl <= MUX_s_1_2_2(or_526_nl, or_524_nl, fsm_output(4));
  mux_494_nl <= MUX_s_1_2_2(mux_493_nl, mux_492_nl, fsm_output(3));
  mux_498_nl <= MUX_s_1_2_2(mux_497_nl, mux_494_nl, fsm_output(0));
  nor_922_nl <= NOT((fsm_output(5)) OR mux_498_nl);
  mux_507_nl <= MUX_s_1_2_2(mux_506_nl, nor_922_nl, fsm_output(2));
  vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_507_nl AND (fsm_output(1));
  nor_908_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(7))));
  nor_909_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(7)));
  mux_519_nl <= MUX_s_1_2_2(nor_908_nl, nor_909_nl, fsm_output(4));
  nor_910_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(7))));
  nor_911_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(7)));
  mux_518_nl <= MUX_s_1_2_2(nor_910_nl, nor_911_nl, fsm_output(4));
  mux_520_nl <= MUX_s_1_2_2(mux_519_nl, mux_518_nl, fsm_output(0));
  and_425_nl <= (fsm_output(6)) AND mux_520_nl;
  or_569_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(7)));
  or_567_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(7));
  mux_516_nl <= MUX_s_1_2_2(or_569_nl, or_567_nl, fsm_output(4));
  or_566_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(7)));
  or_564_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(7));
  mux_515_nl <= MUX_s_1_2_2(or_566_nl, or_564_nl, fsm_output(4));
  mux_517_nl <= MUX_s_1_2_2(mux_516_nl, mux_515_nl, fsm_output(0));
  nor_912_nl <= NOT((fsm_output(6)) OR mux_517_nl);
  mux_521_nl <= MUX_s_1_2_2(and_425_nl, nor_912_nl, fsm_output(3));
  nand_500_nl <= NOT((fsm_output(5)) AND mux_521_nl);
  nor_914_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(7))));
  nor_915_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(7)));
  mux_512_nl <= MUX_s_1_2_2(nor_914_nl, nor_915_nl, fsm_output(4));
  or_558_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR nand_423_cse;
  or_556_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7));
  mux_511_nl <= MUX_s_1_2_2(or_558_nl, or_556_nl, fsm_output(4));
  nor_916_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_511_nl);
  mux_513_nl <= MUX_s_1_2_2(mux_512_nl, nor_916_nl, fsm_output(0));
  nand_41_nl <= NOT((fsm_output(6)) AND mux_513_nl);
  or_554_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      OR nand_442_cse;
  or_552_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(7));
  mux_509_nl <= MUX_s_1_2_2(or_554_nl, or_552_nl, fsm_output(4));
  or_551_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR mux_446_cse;
  mux_510_nl <= MUX_s_1_2_2(mux_509_nl, or_551_nl, fsm_output(0));
  or_555_nl <= (fsm_output(6)) OR mux_510_nl;
  mux_514_nl <= MUX_s_1_2_2(nand_41_nl, or_555_nl, fsm_output(3));
  or_2274_nl <= (fsm_output(5)) OR mux_514_nl;
  mux_522_nl <= MUX_s_1_2_2(nand_500_nl, or_2274_nl, fsm_output(2));
  vec_rsc_0_6_i_we_d_pff <= NOT(mux_522_nl OR (fsm_output(1)));
  nor_901_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_902_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_536_nl <= MUX_s_1_2_2(nor_901_nl, nor_902_nl, fsm_output(0));
  nor_903_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_534_cse);
  nor_904_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_905_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_906_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_530_nl <= MUX_s_1_2_2(nor_905_nl, nor_906_nl, fsm_output(4));
  mux_531_nl <= MUX_s_1_2_2(nor_904_nl, mux_530_nl, fsm_output(3));
  mux_535_nl <= MUX_s_1_2_2(nor_903_nl, mux_531_nl, fsm_output(0));
  mux_537_nl <= MUX_s_1_2_2(mux_536_nl, mux_535_nl, fsm_output(5));
  or_588_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_586_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_527_nl <= MUX_s_1_2_2(or_588_nl, or_586_nl, fsm_output(4));
  or_585_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_583_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_526_nl <= MUX_s_1_2_2(or_585_nl, or_583_nl, fsm_output(4));
  mux_528_nl <= MUX_s_1_2_2(mux_527_nl, mux_526_nl, fsm_output(3));
  or_582_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR nand_443_cse;
  or_580_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_524_nl <= MUX_s_1_2_2(or_582_nl, or_580_nl, fsm_output(4));
  or_579_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_577_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_523_nl <= MUX_s_1_2_2(or_579_nl, or_577_nl, fsm_output(4));
  mux_525_nl <= MUX_s_1_2_2(mux_524_nl, mux_523_nl, fsm_output(3));
  mux_529_nl <= MUX_s_1_2_2(mux_528_nl, mux_525_nl, fsm_output(0));
  nor_907_nl <= NOT((fsm_output(5)) OR mux_529_nl);
  mux_538_nl <= MUX_s_1_2_2(mux_537_nl, nor_907_nl, fsm_output(2));
  vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_538_nl AND (fsm_output(1));
  nor_889_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011"))
      OR nand_445_cse);
  nor_890_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (fsm_output(7)));
  mux_550_nl <= MUX_s_1_2_2(nor_889_nl, nor_890_nl, fsm_output(4));
  nor_891_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR nand_417_cse);
  nor_892_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (fsm_output(7)));
  mux_549_nl <= MUX_s_1_2_2(nor_891_nl, nor_892_nl, fsm_output(4));
  mux_551_nl <= MUX_s_1_2_2(mux_550_nl, mux_549_nl, fsm_output(0));
  and_422_nl <= (fsm_output(6)) AND mux_551_nl;
  or_620_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT (fsm_output(7)));
  or_618_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (fsm_output(7));
  mux_547_nl <= MUX_s_1_2_2(or_620_nl, or_618_nl, fsm_output(4));
  or_617_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011"))
      OR nand_447_cse;
  or_615_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (fsm_output(7));
  mux_546_nl <= MUX_s_1_2_2(or_617_nl, or_615_nl, fsm_output(4));
  mux_548_nl <= MUX_s_1_2_2(mux_547_nl, mux_546_nl, fsm_output(0));
  nor_893_nl <= NOT((fsm_output(6)) OR mux_548_nl);
  mux_552_nl <= MUX_s_1_2_2(and_422_nl, nor_893_nl, fsm_output(3));
  nand_499_nl <= NOT((fsm_output(5)) AND mux_552_nl);
  nor_895_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR nand_419_cse);
  nor_896_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (fsm_output(7)));
  mux_543_nl <= MUX_s_1_2_2(nor_895_nl, nor_896_nl, fsm_output(4));
  nor_897_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR nand_423_cse);
  nor_898_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(7)));
  mux_542_nl <= MUX_s_1_2_2(nor_897_nl, nor_898_nl, fsm_output(4));
  and_423_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_542_nl;
  mux_544_nl <= MUX_s_1_2_2(mux_543_nl, and_423_nl, fsm_output(0));
  nand_47_nl <= NOT((fsm_output(6)) AND mux_544_nl);
  or_606_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      OR nand_442_cse;
  or_604_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (fsm_output(7));
  mux_540_nl <= MUX_s_1_2_2(or_606_nl, or_604_nl, fsm_output(4));
  nand_45_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_477_cse);
  mux_541_nl <= MUX_s_1_2_2(mux_540_nl, nand_45_nl, fsm_output(0));
  or_607_nl <= (fsm_output(6)) OR mux_541_nl;
  mux_545_nl <= MUX_s_1_2_2(nand_47_nl, or_607_nl, fsm_output(3));
  or_2273_nl <= (fsm_output(5)) OR mux_545_nl;
  mux_553_nl <= MUX_s_1_2_2(nand_499_nl, or_2273_nl, fsm_output(2));
  vec_rsc_0_7_i_we_d_pff <= NOT(mux_553_nl OR (fsm_output(1)));
  nor_883_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_884_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_567_nl <= MUX_s_1_2_2(nor_883_nl, nor_884_nl, fsm_output(0));
  and_420_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_534_cse);
  nor_885_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_886_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_887_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_561_nl <= MUX_s_1_2_2(nor_886_nl, nor_887_nl, fsm_output(4));
  mux_562_nl <= MUX_s_1_2_2(nor_885_nl, mux_561_nl, fsm_output(3));
  mux_566_nl <= MUX_s_1_2_2(and_420_nl, mux_562_nl, fsm_output(0));
  mux_568_nl <= MUX_s_1_2_2(mux_567_nl, mux_566_nl, fsm_output(5));
  or_639_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_637_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_558_nl <= MUX_s_1_2_2(or_639_nl, or_637_nl, fsm_output(4));
  or_636_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_634_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_557_nl <= MUX_s_1_2_2(or_636_nl, or_634_nl, fsm_output(4));
  mux_559_nl <= MUX_s_1_2_2(mux_558_nl, mux_557_nl, fsm_output(3));
  or_633_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0011"))
      OR nand_444_cse;
  or_631_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_555_nl <= MUX_s_1_2_2(or_633_nl, or_631_nl, fsm_output(4));
  or_630_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_628_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_554_nl <= MUX_s_1_2_2(or_630_nl, or_628_nl, fsm_output(4));
  mux_556_nl <= MUX_s_1_2_2(mux_555_nl, mux_554_nl, fsm_output(3));
  mux_560_nl <= MUX_s_1_2_2(mux_559_nl, mux_556_nl, fsm_output(0));
  nor_888_nl <= NOT((fsm_output(5)) OR mux_560_nl);
  mux_569_nl <= MUX_s_1_2_2(mux_568_nl, nor_888_nl, fsm_output(2));
  vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_569_nl AND (fsm_output(1));
  nor_874_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(7))));
  nor_875_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(7)));
  mux_581_nl <= MUX_s_1_2_2(nor_874_nl, nor_875_nl, fsm_output(4));
  nor_876_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(7))));
  nor_877_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(7)));
  mux_580_nl <= MUX_s_1_2_2(nor_876_nl, nor_877_nl, fsm_output(4));
  mux_582_nl <= MUX_s_1_2_2(mux_581_nl, mux_580_nl, fsm_output(0));
  and_419_nl <= (fsm_output(6)) AND mux_582_nl;
  or_673_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(7)));
  or_671_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(7));
  mux_578_nl <= MUX_s_1_2_2(or_673_nl, or_671_nl, fsm_output(4));
  or_670_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(7)));
  or_668_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(7));
  mux_577_nl <= MUX_s_1_2_2(or_670_nl, or_668_nl, fsm_output(4));
  mux_579_nl <= MUX_s_1_2_2(mux_578_nl, mux_577_nl, fsm_output(0));
  nor_878_nl <= NOT((fsm_output(6)) OR mux_579_nl);
  mux_583_nl <= MUX_s_1_2_2(and_419_nl, nor_878_nl, fsm_output(3));
  nand_498_nl <= NOT((fsm_output(5)) AND mux_583_nl);
  nor_880_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(7))));
  nor_881_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(7)));
  mux_574_nl <= MUX_s_1_2_2(nor_880_nl, nor_881_nl, fsm_output(4));
  or_662_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7)));
  or_660_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7));
  mux_573_nl <= MUX_s_1_2_2(or_662_nl, or_660_nl, fsm_output(4));
  nor_882_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_573_nl);
  mux_575_nl <= MUX_s_1_2_2(mux_574_nl, nor_882_nl, fsm_output(0));
  nand_52_nl <= NOT((fsm_output(6)) AND mux_575_nl);
  or_658_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(7)));
  or_656_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(7));
  mux_571_nl <= MUX_s_1_2_2(or_658_nl, or_656_nl, fsm_output(4));
  or_655_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR mux_570_cse;
  mux_572_nl <= MUX_s_1_2_2(mux_571_nl, or_655_nl, fsm_output(0));
  or_659_nl <= (fsm_output(6)) OR mux_572_nl;
  mux_576_nl <= MUX_s_1_2_2(nand_52_nl, or_659_nl, fsm_output(3));
  or_2272_nl <= (fsm_output(5)) OR mux_576_nl;
  mux_584_nl <= MUX_s_1_2_2(nand_498_nl, or_2272_nl, fsm_output(2));
  vec_rsc_0_8_i_we_d_pff <= NOT(mux_584_nl OR (fsm_output(1)));
  nor_867_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_868_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_598_nl <= MUX_s_1_2_2(nor_867_nl, nor_868_nl, fsm_output(0));
  nor_869_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_596_cse);
  nor_870_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_871_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_872_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_592_nl <= MUX_s_1_2_2(nor_871_nl, nor_872_nl, fsm_output(4));
  mux_593_nl <= MUX_s_1_2_2(nor_870_nl, mux_592_nl, fsm_output(3));
  mux_597_nl <= MUX_s_1_2_2(nor_869_nl, mux_593_nl, fsm_output(0));
  mux_599_nl <= MUX_s_1_2_2(mux_598_nl, mux_597_nl, fsm_output(5));
  or_692_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_690_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_589_nl <= MUX_s_1_2_2(or_692_nl, or_690_nl, fsm_output(4));
  or_689_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_687_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_588_nl <= MUX_s_1_2_2(or_689_nl, or_687_nl, fsm_output(4));
  mux_590_nl <= MUX_s_1_2_2(mux_589_nl, mux_588_nl, fsm_output(3));
  or_686_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR nand_443_cse;
  or_684_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_586_nl <= MUX_s_1_2_2(or_686_nl, or_684_nl, fsm_output(4));
  or_683_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_681_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_585_nl <= MUX_s_1_2_2(or_683_nl, or_681_nl, fsm_output(4));
  mux_587_nl <= MUX_s_1_2_2(mux_586_nl, mux_585_nl, fsm_output(3));
  mux_591_nl <= MUX_s_1_2_2(mux_590_nl, mux_587_nl, fsm_output(0));
  nor_873_nl <= NOT((fsm_output(5)) OR mux_591_nl);
  mux_600_nl <= MUX_s_1_2_2(mux_599_nl, nor_873_nl, fsm_output(2));
  vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_600_nl AND (fsm_output(1));
  nor_855_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_445_cse);
  nor_856_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (fsm_output(7)));
  mux_612_nl <= MUX_s_1_2_2(nor_855_nl, nor_856_nl, fsm_output(4));
  nor_857_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_446_cse);
  nor_858_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (fsm_output(7)));
  mux_611_nl <= MUX_s_1_2_2(nor_857_nl, nor_858_nl, fsm_output(4));
  mux_613_nl <= MUX_s_1_2_2(mux_612_nl, mux_611_nl, fsm_output(0));
  and_416_nl <= (fsm_output(6)) AND mux_613_nl;
  or_724_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT (fsm_output(7)));
  or_722_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (fsm_output(7));
  mux_609_nl <= MUX_s_1_2_2(or_724_nl, or_722_nl, fsm_output(4));
  or_721_nl <= (COMP_LOOP_acc_1_cse_6_sva(2)) OR (COMP_LOOP_acc_1_cse_6_sva(1)) OR
      (COMP_LOOP_acc_1_cse_6_sva(4)) OR nand_411_cse;
  or_719_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (fsm_output(7));
  mux_608_nl <= MUX_s_1_2_2(or_721_nl, or_719_nl, fsm_output(4));
  mux_610_nl <= MUX_s_1_2_2(mux_609_nl, mux_608_nl, fsm_output(0));
  nor_859_nl <= NOT((fsm_output(6)) OR mux_610_nl);
  mux_614_nl <= MUX_s_1_2_2(and_416_nl, nor_859_nl, fsm_output(3));
  nand_497_nl <= NOT((fsm_output(5)) AND mux_614_nl);
  nor_861_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_448_cse);
  nor_862_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (fsm_output(7)));
  mux_605_nl <= MUX_s_1_2_2(nor_861_nl, nor_862_nl, fsm_output(4));
  nor_863_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(7))));
  nor_864_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(7)));
  mux_604_nl <= MUX_s_1_2_2(nor_863_nl, nor_864_nl, fsm_output(4));
  and_417_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_604_nl;
  mux_606_nl <= MUX_s_1_2_2(mux_605_nl, and_417_nl, fsm_output(0));
  nand_58_nl <= NOT((fsm_output(6)) AND mux_606_nl);
  or_710_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT (fsm_output(7)));
  or_708_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (fsm_output(7));
  mux_602_nl <= MUX_s_1_2_2(or_710_nl, or_708_nl, fsm_output(4));
  nand_56_nl <= NOT(nor_98_cse AND mux_601_cse);
  mux_603_nl <= MUX_s_1_2_2(mux_602_nl, nand_56_nl, fsm_output(0));
  or_711_nl <= (fsm_output(6)) OR mux_603_nl;
  mux_607_nl <= MUX_s_1_2_2(nand_58_nl, or_711_nl, fsm_output(3));
  or_2271_nl <= (fsm_output(5)) OR mux_607_nl;
  mux_615_nl <= MUX_s_1_2_2(nand_497_nl, or_2271_nl, fsm_output(2));
  vec_rsc_0_9_i_we_d_pff <= NOT(mux_615_nl OR (fsm_output(1)));
  nor_849_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_850_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_629_nl <= MUX_s_1_2_2(nor_849_nl, nor_850_nl, fsm_output(0));
  and_414_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_596_cse);
  nor_851_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_852_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_853_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_623_nl <= MUX_s_1_2_2(nor_852_nl, nor_853_nl, fsm_output(4));
  mux_624_nl <= MUX_s_1_2_2(nor_851_nl, mux_623_nl, fsm_output(3));
  mux_628_nl <= MUX_s_1_2_2(and_414_nl, mux_624_nl, fsm_output(0));
  mux_630_nl <= MUX_s_1_2_2(mux_629_nl, mux_628_nl, fsm_output(5));
  or_743_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_741_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_620_nl <= MUX_s_1_2_2(or_743_nl, or_741_nl, fsm_output(4));
  or_740_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_738_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_619_nl <= MUX_s_1_2_2(or_740_nl, or_738_nl, fsm_output(4));
  mux_621_nl <= MUX_s_1_2_2(mux_620_nl, mux_619_nl, fsm_output(3));
  or_737_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_444_cse;
  or_735_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_617_nl <= MUX_s_1_2_2(or_737_nl, or_735_nl, fsm_output(4));
  or_734_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_732_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_616_nl <= MUX_s_1_2_2(or_734_nl, or_732_nl, fsm_output(4));
  mux_618_nl <= MUX_s_1_2_2(mux_617_nl, mux_616_nl, fsm_output(3));
  mux_622_nl <= MUX_s_1_2_2(mux_621_nl, mux_618_nl, fsm_output(0));
  nor_854_nl <= NOT((fsm_output(5)) OR mux_622_nl);
  mux_631_nl <= MUX_s_1_2_2(mux_630_nl, nor_854_nl, fsm_output(2));
  vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_631_nl AND (fsm_output(1));
  nor_840_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(7))));
  nor_841_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(7)));
  mux_643_nl <= MUX_s_1_2_2(nor_840_nl, nor_841_nl, fsm_output(4));
  nor_842_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(7))));
  nor_843_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(7)));
  mux_642_nl <= MUX_s_1_2_2(nor_842_nl, nor_843_nl, fsm_output(4));
  mux_644_nl <= MUX_s_1_2_2(mux_643_nl, mux_642_nl, fsm_output(0));
  and_413_nl <= (fsm_output(6)) AND mux_644_nl;
  or_777_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(7)));
  or_775_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(7));
  mux_640_nl <= MUX_s_1_2_2(or_777_nl, or_775_nl, fsm_output(4));
  or_774_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(7)));
  or_772_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(7));
  mux_639_nl <= MUX_s_1_2_2(or_774_nl, or_772_nl, fsm_output(4));
  mux_641_nl <= MUX_s_1_2_2(mux_640_nl, mux_639_nl, fsm_output(0));
  nor_844_nl <= NOT((fsm_output(6)) OR mux_641_nl);
  mux_645_nl <= MUX_s_1_2_2(and_413_nl, nor_844_nl, fsm_output(3));
  nand_496_nl <= NOT((fsm_output(5)) AND mux_645_nl);
  nor_846_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(7))));
  nor_847_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(7)));
  mux_636_nl <= MUX_s_1_2_2(nor_846_nl, nor_847_nl, fsm_output(4));
  or_766_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"))
      OR nand_441_cse;
  or_764_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7));
  mux_635_nl <= MUX_s_1_2_2(or_766_nl, or_764_nl, fsm_output(4));
  nor_848_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_635_nl);
  mux_637_nl <= MUX_s_1_2_2(mux_636_nl, nor_848_nl, fsm_output(0));
  nand_63_nl <= NOT((fsm_output(6)) AND mux_637_nl);
  or_762_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      OR nand_442_cse;
  or_760_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(7));
  mux_633_nl <= MUX_s_1_2_2(or_762_nl, or_760_nl, fsm_output(4));
  or_759_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR mux_570_cse;
  mux_634_nl <= MUX_s_1_2_2(mux_633_nl, or_759_nl, fsm_output(0));
  or_763_nl <= (fsm_output(6)) OR mux_634_nl;
  mux_638_nl <= MUX_s_1_2_2(nand_63_nl, or_763_nl, fsm_output(3));
  or_2270_nl <= (fsm_output(5)) OR mux_638_nl;
  mux_646_nl <= MUX_s_1_2_2(nand_496_nl, or_2270_nl, fsm_output(2));
  vec_rsc_0_10_i_we_d_pff <= NOT(mux_646_nl OR (fsm_output(1)));
  nor_833_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_834_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_660_nl <= MUX_s_1_2_2(nor_833_nl, nor_834_nl, fsm_output(0));
  nor_835_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_658_cse);
  nor_836_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_837_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_838_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_654_nl <= MUX_s_1_2_2(nor_837_nl, nor_838_nl, fsm_output(4));
  mux_655_nl <= MUX_s_1_2_2(nor_836_nl, mux_654_nl, fsm_output(3));
  mux_659_nl <= MUX_s_1_2_2(nor_835_nl, mux_655_nl, fsm_output(0));
  mux_661_nl <= MUX_s_1_2_2(mux_660_nl, mux_659_nl, fsm_output(5));
  or_796_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_794_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_651_nl <= MUX_s_1_2_2(or_796_nl, or_794_nl, fsm_output(4));
  or_793_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_791_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_650_nl <= MUX_s_1_2_2(or_793_nl, or_791_nl, fsm_output(4));
  mux_652_nl <= MUX_s_1_2_2(mux_651_nl, mux_650_nl, fsm_output(3));
  or_790_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR nand_443_cse;
  or_788_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_648_nl <= MUX_s_1_2_2(or_790_nl, or_788_nl, fsm_output(4));
  or_787_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_785_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_647_nl <= MUX_s_1_2_2(or_787_nl, or_785_nl, fsm_output(4));
  mux_649_nl <= MUX_s_1_2_2(mux_648_nl, mux_647_nl, fsm_output(3));
  mux_653_nl <= MUX_s_1_2_2(mux_652_nl, mux_649_nl, fsm_output(0));
  nor_839_nl <= NOT((fsm_output(5)) OR mux_653_nl);
  mux_662_nl <= MUX_s_1_2_2(mux_661_nl, nor_839_nl, fsm_output(2));
  vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_662_nl AND (fsm_output(1));
  nor_821_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101"))
      OR nand_445_cse);
  nor_822_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (fsm_output(7)));
  mux_674_nl <= MUX_s_1_2_2(nor_821_nl, nor_822_nl, fsm_output(4));
  nor_823_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("010"))
      OR nand_435_cse);
  nor_824_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (fsm_output(7)));
  mux_673_nl <= MUX_s_1_2_2(nor_823_nl, nor_824_nl, fsm_output(4));
  mux_675_nl <= MUX_s_1_2_2(mux_674_nl, mux_673_nl, fsm_output(0));
  and_410_nl <= (fsm_output(6)) AND mux_675_nl;
  or_828_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT (fsm_output(7)));
  or_826_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (fsm_output(7));
  mux_671_nl <= MUX_s_1_2_2(or_828_nl, or_826_nl, fsm_output(4));
  or_825_nl <= (COMP_LOOP_acc_1_cse_6_sva(2)) OR (NOT (COMP_LOOP_acc_1_cse_6_sva(1)))
      OR (COMP_LOOP_acc_1_cse_6_sva(4)) OR nand_411_cse;
  or_823_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (fsm_output(7));
  mux_670_nl <= MUX_s_1_2_2(or_825_nl, or_823_nl, fsm_output(4));
  mux_672_nl <= MUX_s_1_2_2(mux_671_nl, mux_670_nl, fsm_output(0));
  nor_825_nl <= NOT((fsm_output(6)) OR mux_672_nl);
  mux_676_nl <= MUX_s_1_2_2(and_410_nl, nor_825_nl, fsm_output(3));
  nand_495_nl <= NOT((fsm_output(5)) AND mux_676_nl);
  nor_827_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("010"))
      OR nand_437_cse);
  nor_828_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (fsm_output(7)));
  mux_667_nl <= MUX_s_1_2_2(nor_827_nl, nor_828_nl, fsm_output(4));
  nor_829_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"))
      OR nand_441_cse);
  nor_830_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(7)));
  mux_666_nl <= MUX_s_1_2_2(nor_829_nl, nor_830_nl, fsm_output(4));
  and_411_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_666_nl;
  mux_668_nl <= MUX_s_1_2_2(mux_667_nl, and_411_nl, fsm_output(0));
  nand_69_nl <= NOT((fsm_output(6)) AND mux_668_nl);
  or_814_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      OR nand_442_cse;
  or_812_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (fsm_output(7));
  mux_664_nl <= MUX_s_1_2_2(or_814_nl, or_812_nl, fsm_output(4));
  nand_67_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_601_cse);
  mux_665_nl <= MUX_s_1_2_2(mux_664_nl, nand_67_nl, fsm_output(0));
  or_815_nl <= (fsm_output(6)) OR mux_665_nl;
  mux_669_nl <= MUX_s_1_2_2(nand_69_nl, or_815_nl, fsm_output(3));
  or_2269_nl <= (fsm_output(5)) OR mux_669_nl;
  mux_677_nl <= MUX_s_1_2_2(nand_495_nl, or_2269_nl, fsm_output(2));
  vec_rsc_0_11_i_we_d_pff <= NOT(mux_677_nl OR (fsm_output(1)));
  nor_815_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_816_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_691_nl <= MUX_s_1_2_2(nor_815_nl, nor_816_nl, fsm_output(0));
  and_408_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_658_cse);
  nor_817_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_818_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_819_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_685_nl <= MUX_s_1_2_2(nor_818_nl, nor_819_nl, fsm_output(4));
  mux_686_nl <= MUX_s_1_2_2(nor_817_nl, mux_685_nl, fsm_output(3));
  mux_690_nl <= MUX_s_1_2_2(and_408_nl, mux_686_nl, fsm_output(0));
  mux_692_nl <= MUX_s_1_2_2(mux_691_nl, mux_690_nl, fsm_output(5));
  or_847_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_845_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_682_nl <= MUX_s_1_2_2(or_847_nl, or_845_nl, fsm_output(4));
  or_844_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_842_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_681_nl <= MUX_s_1_2_2(or_844_nl, or_842_nl, fsm_output(4));
  mux_683_nl <= MUX_s_1_2_2(mux_682_nl, mux_681_nl, fsm_output(3));
  or_841_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0101"))
      OR nand_444_cse;
  or_839_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_679_nl <= MUX_s_1_2_2(or_841_nl, or_839_nl, fsm_output(4));
  or_838_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_836_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_678_nl <= MUX_s_1_2_2(or_838_nl, or_836_nl, fsm_output(4));
  mux_680_nl <= MUX_s_1_2_2(mux_679_nl, mux_678_nl, fsm_output(3));
  mux_684_nl <= MUX_s_1_2_2(mux_683_nl, mux_680_nl, fsm_output(0));
  nor_820_nl <= NOT((fsm_output(5)) OR mux_684_nl);
  mux_693_nl <= MUX_s_1_2_2(mux_692_nl, nor_820_nl, fsm_output(2));
  vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_693_nl AND (fsm_output(1));
  nor_806_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(7))));
  nor_807_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(7)));
  mux_705_nl <= MUX_s_1_2_2(nor_806_nl, nor_807_nl, fsm_output(4));
  nor_808_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(7))));
  nor_809_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(7)));
  mux_704_nl <= MUX_s_1_2_2(nor_808_nl, nor_809_nl, fsm_output(4));
  mux_706_nl <= MUX_s_1_2_2(mux_705_nl, mux_704_nl, fsm_output(0));
  and_407_nl <= (fsm_output(6)) AND mux_706_nl;
  or_881_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(7)));
  or_879_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(7));
  mux_702_nl <= MUX_s_1_2_2(or_881_nl, or_879_nl, fsm_output(4));
  or_878_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(7)));
  or_876_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(7));
  mux_701_nl <= MUX_s_1_2_2(or_878_nl, or_876_nl, fsm_output(4));
  mux_703_nl <= MUX_s_1_2_2(mux_702_nl, mux_701_nl, fsm_output(0));
  nor_810_nl <= NOT((fsm_output(6)) OR mux_703_nl);
  mux_707_nl <= MUX_s_1_2_2(and_407_nl, nor_810_nl, fsm_output(3));
  nand_494_nl <= NOT((fsm_output(5)) AND mux_707_nl);
  nor_812_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(7))));
  nor_813_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(7)));
  mux_698_nl <= MUX_s_1_2_2(nor_812_nl, nor_813_nl, fsm_output(4));
  or_870_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7)));
  or_868_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7));
  mux_697_nl <= MUX_s_1_2_2(or_870_nl, or_868_nl, fsm_output(4));
  nor_814_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_697_nl);
  mux_699_nl <= MUX_s_1_2_2(mux_698_nl, nor_814_nl, fsm_output(0));
  nand_74_nl <= NOT((fsm_output(6)) AND mux_699_nl);
  or_866_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(7)));
  or_864_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(7));
  mux_695_nl <= MUX_s_1_2_2(or_866_nl, or_864_nl, fsm_output(4));
  or_863_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR mux_694_cse;
  mux_696_nl <= MUX_s_1_2_2(mux_695_nl, or_863_nl, fsm_output(0));
  or_867_nl <= (fsm_output(6)) OR mux_696_nl;
  mux_700_nl <= MUX_s_1_2_2(nand_74_nl, or_867_nl, fsm_output(3));
  or_2268_nl <= (fsm_output(5)) OR mux_700_nl;
  mux_708_nl <= MUX_s_1_2_2(nand_494_nl, or_2268_nl, fsm_output(2));
  vec_rsc_0_12_i_we_d_pff <= NOT(mux_708_nl OR (fsm_output(1)));
  nor_799_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_800_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_722_nl <= MUX_s_1_2_2(nor_799_nl, nor_800_nl, fsm_output(0));
  nor_801_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_720_cse);
  nor_802_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_803_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_804_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_716_nl <= MUX_s_1_2_2(nor_803_nl, nor_804_nl, fsm_output(4));
  mux_717_nl <= MUX_s_1_2_2(nor_802_nl, mux_716_nl, fsm_output(3));
  mux_721_nl <= MUX_s_1_2_2(nor_801_nl, mux_717_nl, fsm_output(0));
  mux_723_nl <= MUX_s_1_2_2(mux_722_nl, mux_721_nl, fsm_output(5));
  or_900_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_898_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_713_nl <= MUX_s_1_2_2(or_900_nl, or_898_nl, fsm_output(4));
  or_897_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_895_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_712_nl <= MUX_s_1_2_2(or_897_nl, or_895_nl, fsm_output(4));
  mux_714_nl <= MUX_s_1_2_2(mux_713_nl, mux_712_nl, fsm_output(3));
  or_894_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR nand_443_cse;
  or_892_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_710_nl <= MUX_s_1_2_2(or_894_nl, or_892_nl, fsm_output(4));
  or_891_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_889_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_709_nl <= MUX_s_1_2_2(or_891_nl, or_889_nl, fsm_output(4));
  mux_711_nl <= MUX_s_1_2_2(mux_710_nl, mux_709_nl, fsm_output(3));
  mux_715_nl <= MUX_s_1_2_2(mux_714_nl, mux_711_nl, fsm_output(0));
  nor_805_nl <= NOT((fsm_output(5)) OR mux_715_nl);
  mux_724_nl <= MUX_s_1_2_2(mux_723_nl, nor_805_nl, fsm_output(2));
  vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_724_nl AND (fsm_output(1));
  nor_787_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_445_cse);
  nor_788_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (fsm_output(7)));
  mux_736_nl <= MUX_s_1_2_2(nor_787_nl, nor_788_nl, fsm_output(4));
  nor_789_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_446_cse);
  nor_790_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (fsm_output(7)));
  mux_735_nl <= MUX_s_1_2_2(nor_789_nl, nor_790_nl, fsm_output(4));
  mux_737_nl <= MUX_s_1_2_2(mux_736_nl, mux_735_nl, fsm_output(0));
  and_404_nl <= (fsm_output(6)) AND mux_737_nl;
  or_932_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT (fsm_output(7)));
  or_930_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (fsm_output(7));
  mux_733_nl <= MUX_s_1_2_2(or_932_nl, or_930_nl, fsm_output(4));
  or_929_nl <= (NOT (COMP_LOOP_acc_1_cse_6_sva(2))) OR (COMP_LOOP_acc_1_cse_6_sva(1))
      OR (COMP_LOOP_acc_1_cse_6_sva(4)) OR nand_411_cse;
  or_927_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (fsm_output(7));
  mux_732_nl <= MUX_s_1_2_2(or_929_nl, or_927_nl, fsm_output(4));
  mux_734_nl <= MUX_s_1_2_2(mux_733_nl, mux_732_nl, fsm_output(0));
  nor_791_nl <= NOT((fsm_output(6)) OR mux_734_nl);
  mux_738_nl <= MUX_s_1_2_2(and_404_nl, nor_791_nl, fsm_output(3));
  nand_493_nl <= NOT((fsm_output(5)) AND mux_738_nl);
  nor_793_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_448_cse);
  nor_794_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (fsm_output(7)));
  mux_729_nl <= MUX_s_1_2_2(nor_793_nl, nor_794_nl, fsm_output(4));
  nor_795_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(7))));
  nor_796_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(7)));
  mux_728_nl <= MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output(4));
  and_405_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_728_nl;
  mux_730_nl <= MUX_s_1_2_2(mux_729_nl, and_405_nl, fsm_output(0));
  nand_80_nl <= NOT((fsm_output(6)) AND mux_730_nl);
  or_918_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT (fsm_output(7)));
  or_916_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (fsm_output(7));
  mux_726_nl <= MUX_s_1_2_2(or_918_nl, or_916_nl, fsm_output(4));
  nand_78_nl <= NOT(nor_98_cse AND mux_725_cse);
  mux_727_nl <= MUX_s_1_2_2(mux_726_nl, nand_78_nl, fsm_output(0));
  or_919_nl <= (fsm_output(6)) OR mux_727_nl;
  mux_731_nl <= MUX_s_1_2_2(nand_80_nl, or_919_nl, fsm_output(3));
  or_2267_nl <= (fsm_output(5)) OR mux_731_nl;
  mux_739_nl <= MUX_s_1_2_2(nand_493_nl, or_2267_nl, fsm_output(2));
  vec_rsc_0_13_i_we_d_pff <= NOT(mux_739_nl OR (fsm_output(1)));
  nor_781_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_782_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_753_nl <= MUX_s_1_2_2(nor_781_nl, nor_782_nl, fsm_output(0));
  and_402_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_720_cse);
  nor_783_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_784_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_785_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_747_nl <= MUX_s_1_2_2(nor_784_nl, nor_785_nl, fsm_output(4));
  mux_748_nl <= MUX_s_1_2_2(nor_783_nl, mux_747_nl, fsm_output(3));
  mux_752_nl <= MUX_s_1_2_2(and_402_nl, mux_748_nl, fsm_output(0));
  mux_754_nl <= MUX_s_1_2_2(mux_753_nl, mux_752_nl, fsm_output(5));
  or_951_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_949_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_744_nl <= MUX_s_1_2_2(or_951_nl, or_949_nl, fsm_output(4));
  or_948_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_946_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_743_nl <= MUX_s_1_2_2(or_948_nl, or_946_nl, fsm_output(4));
  mux_745_nl <= MUX_s_1_2_2(mux_744_nl, mux_743_nl, fsm_output(3));
  or_945_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_444_cse;
  or_943_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_741_nl <= MUX_s_1_2_2(or_945_nl, or_943_nl, fsm_output(4));
  or_942_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_940_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_740_nl <= MUX_s_1_2_2(or_942_nl, or_940_nl, fsm_output(4));
  mux_742_nl <= MUX_s_1_2_2(mux_741_nl, mux_740_nl, fsm_output(3));
  mux_746_nl <= MUX_s_1_2_2(mux_745_nl, mux_742_nl, fsm_output(0));
  nor_786_nl <= NOT((fsm_output(5)) OR mux_746_nl);
  mux_755_nl <= MUX_s_1_2_2(mux_754_nl, nor_786_nl, fsm_output(2));
  vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_755_nl AND (fsm_output(1));
  nor_772_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(7))));
  nor_773_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(7)));
  mux_767_nl <= MUX_s_1_2_2(nor_772_nl, nor_773_nl, fsm_output(4));
  nor_774_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(7))));
  nor_775_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(7)));
  mux_766_nl <= MUX_s_1_2_2(nor_774_nl, nor_775_nl, fsm_output(4));
  mux_768_nl <= MUX_s_1_2_2(mux_767_nl, mux_766_nl, fsm_output(0));
  and_401_nl <= (fsm_output(6)) AND mux_768_nl;
  or_984_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(7)));
  or_982_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(7));
  mux_764_nl <= MUX_s_1_2_2(or_984_nl, or_982_nl, fsm_output(4));
  or_981_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(7)));
  or_979_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(7));
  mux_763_nl <= MUX_s_1_2_2(or_981_nl, or_979_nl, fsm_output(4));
  mux_765_nl <= MUX_s_1_2_2(mux_764_nl, mux_763_nl, fsm_output(0));
  nor_776_nl <= NOT((fsm_output(6)) OR mux_765_nl);
  mux_769_nl <= MUX_s_1_2_2(and_401_nl, nor_776_nl, fsm_output(3));
  nand_492_nl <= NOT((fsm_output(5)) AND mux_769_nl);
  nor_778_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(7))));
  nor_779_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(7)));
  mux_760_nl <= MUX_s_1_2_2(nor_778_nl, nor_779_nl, fsm_output(4));
  or_973_nl <= (COMP_LOOP_acc_14_psp_sva(3)) OR nand_385_cse;
  or_972_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7));
  mux_759_nl <= MUX_s_1_2_2(or_973_nl, or_972_nl, fsm_output(4));
  nor_780_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_759_nl);
  mux_761_nl <= MUX_s_1_2_2(mux_760_nl, nor_780_nl, fsm_output(0));
  nand_85_nl <= NOT((fsm_output(6)) AND mux_761_nl);
  or_970_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      OR nand_442_cse;
  or_968_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(7));
  mux_757_nl <= MUX_s_1_2_2(or_970_nl, or_968_nl, fsm_output(4));
  or_967_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR mux_694_cse;
  mux_758_nl <= MUX_s_1_2_2(mux_757_nl, or_967_nl, fsm_output(0));
  or_971_nl <= (fsm_output(6)) OR mux_758_nl;
  mux_762_nl <= MUX_s_1_2_2(nand_85_nl, or_971_nl, fsm_output(3));
  or_2266_nl <= (fsm_output(5)) OR mux_762_nl;
  mux_770_nl <= MUX_s_1_2_2(nand_492_nl, or_2266_nl, fsm_output(2));
  vec_rsc_0_14_i_we_d_pff <= NOT(mux_770_nl OR (fsm_output(1)));
  nor_765_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_766_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_784_nl <= MUX_s_1_2_2(nor_765_nl, nor_766_nl, fsm_output(0));
  nor_767_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_782_cse);
  nor_768_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_769_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_770_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_778_nl <= MUX_s_1_2_2(nor_769_nl, nor_770_nl, fsm_output(4));
  mux_779_nl <= MUX_s_1_2_2(nor_768_nl, mux_778_nl, fsm_output(3));
  mux_783_nl <= MUX_s_1_2_2(nor_767_nl, mux_779_nl, fsm_output(0));
  mux_785_nl <= MUX_s_1_2_2(mux_784_nl, mux_783_nl, fsm_output(5));
  or_1003_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1001_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_775_nl <= MUX_s_1_2_2(or_1003_nl, or_1001_nl, fsm_output(4));
  or_1000_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_998_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_774_nl <= MUX_s_1_2_2(or_1000_nl, or_998_nl, fsm_output(4));
  mux_776_nl <= MUX_s_1_2_2(mux_775_nl, mux_774_nl, fsm_output(3));
  or_997_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR nand_443_cse;
  or_995_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_772_nl <= MUX_s_1_2_2(or_997_nl, or_995_nl, fsm_output(4));
  or_994_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_992_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_771_nl <= MUX_s_1_2_2(or_994_nl, or_992_nl, fsm_output(4));
  mux_773_nl <= MUX_s_1_2_2(mux_772_nl, mux_771_nl, fsm_output(3));
  mux_777_nl <= MUX_s_1_2_2(mux_776_nl, mux_773_nl, fsm_output(0));
  nor_771_nl <= NOT((fsm_output(5)) OR mux_777_nl);
  mux_786_nl <= MUX_s_1_2_2(mux_785_nl, nor_771_nl, fsm_output(2));
  vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_786_nl AND (fsm_output(1));
  nor_753_nl <= NOT(nand_371_cse OR nand_445_cse);
  nor_754_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (fsm_output(7)));
  mux_798_nl <= MUX_s_1_2_2(nor_753_nl, nor_754_nl, fsm_output(4));
  nor_755_nl <= NOT((COMP_LOOP_acc_1_cse_sva(4)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(7)))));
  nor_756_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (fsm_output(7)));
  mux_797_nl <= MUX_s_1_2_2(nor_755_nl, nor_756_nl, fsm_output(4));
  mux_799_nl <= MUX_s_1_2_2(mux_798_nl, mux_797_nl, fsm_output(0));
  and_398_nl <= (fsm_output(6)) AND mux_799_nl;
  nand_516_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND (fsm_output(7)));
  or_1031_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (fsm_output(7));
  mux_795_nl <= MUX_s_1_2_2(nand_516_nl, or_1031_nl, fsm_output(4));
  or_1030_nl <= (NOT (COMP_LOOP_acc_1_cse_6_sva(2))) OR (NOT (COMP_LOOP_acc_1_cse_6_sva(1)))
      OR (COMP_LOOP_acc_1_cse_6_sva(4)) OR nand_411_cse;
  or_1028_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (fsm_output(7));
  mux_794_nl <= MUX_s_1_2_2(or_1030_nl, or_1028_nl, fsm_output(4));
  mux_796_nl <= MUX_s_1_2_2(mux_795_nl, mux_794_nl, fsm_output(0));
  nor_757_nl <= NOT((fsm_output(6)) OR mux_796_nl);
  mux_800_nl <= MUX_s_1_2_2(and_398_nl, nor_757_nl, fsm_output(3));
  nand_491_nl <= NOT((fsm_output(5)) AND mux_800_nl);
  nor_759_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_7_sva(4)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(7)))));
  nor_760_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (fsm_output(7)));
  mux_791_nl <= MUX_s_1_2_2(nor_759_nl, nor_760_nl, fsm_output(4));
  nor_761_nl <= NOT((COMP_LOOP_acc_14_psp_sva(3)) OR nand_385_cse);
  nor_762_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(7)));
  mux_790_nl <= MUX_s_1_2_2(nor_761_nl, nor_762_nl, fsm_output(4));
  and_399_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_790_nl;
  mux_792_nl <= MUX_s_1_2_2(mux_791_nl, and_399_nl, fsm_output(0));
  nand_91_nl <= NOT((fsm_output(6)) AND mux_792_nl);
  or_1021_nl <= (NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      AND (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) AND (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(4)))))
      OR nand_442_cse;
  or_1019_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (fsm_output(7));
  mux_788_nl <= MUX_s_1_2_2(or_1021_nl, or_1019_nl, fsm_output(4));
  nand_89_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_725_cse);
  mux_789_nl <= MUX_s_1_2_2(mux_788_nl, nand_89_nl, fsm_output(0));
  or_1022_nl <= (fsm_output(6)) OR mux_789_nl;
  mux_793_nl <= MUX_s_1_2_2(nand_91_nl, or_1022_nl, fsm_output(3));
  or_2265_nl <= (fsm_output(5)) OR mux_793_nl;
  mux_801_nl <= MUX_s_1_2_2(nand_491_nl, or_2265_nl, fsm_output(2));
  vec_rsc_0_15_i_we_d_pff <= NOT(mux_801_nl OR (fsm_output(1)));
  nor_748_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_749_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_815_nl <= MUX_s_1_2_2(nor_748_nl, nor_749_nl, fsm_output(0));
  and_395_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_782_cse);
  and_396_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND (fsm_output(4)) AND (fsm_output(6)) AND (NOT (fsm_output(7)));
  and_527_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  nor_751_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_809_nl <= MUX_s_1_2_2(and_527_nl, nor_751_nl, fsm_output(4));
  mux_810_nl <= MUX_s_1_2_2(and_396_nl, mux_809_nl, fsm_output(3));
  mux_814_nl <= MUX_s_1_2_2(and_395_nl, mux_810_nl, fsm_output(0));
  mux_816_nl <= MUX_s_1_2_2(mux_815_nl, mux_814_nl, fsm_output(5));
  or_1051_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)) OR nand_443_cse;
  nand_369_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("01")));
  mux_806_nl <= MUX_s_1_2_2(or_1051_nl, nand_369_nl, fsm_output(4));
  nand_515_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1046_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_805_nl <= MUX_s_1_2_2(nand_515_nl, or_1046_nl, fsm_output(4));
  mux_807_nl <= MUX_s_1_2_2(mux_806_nl, mux_805_nl, fsm_output(3));
  or_1045_nl <= nand_371_cse OR nand_444_cse;
  nand_373_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_803_nl <= MUX_s_1_2_2(or_1045_nl, nand_373_nl, fsm_output(4));
  nand_471_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  or_1040_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_802_nl <= MUX_s_1_2_2(nand_471_nl, or_1040_nl, fsm_output(4));
  mux_804_nl <= MUX_s_1_2_2(mux_803_nl, mux_802_nl, fsm_output(3));
  mux_808_nl <= MUX_s_1_2_2(mux_807_nl, mux_804_nl, fsm_output(0));
  nor_752_nl <= NOT((fsm_output(5)) OR mux_808_nl);
  mux_817_nl <= MUX_s_1_2_2(mux_816_nl, nor_752_nl, fsm_output(2));
  vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_817_nl AND (fsm_output(1));
  nor_739_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (fsm_output(7))));
  nor_740_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(7)));
  mux_829_nl <= MUX_s_1_2_2(nor_739_nl, nor_740_nl, fsm_output(4));
  nor_741_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (fsm_output(7))));
  nor_742_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(7)));
  mux_828_nl <= MUX_s_1_2_2(nor_741_nl, nor_742_nl, fsm_output(4));
  mux_830_nl <= MUX_s_1_2_2(mux_829_nl, mux_828_nl, fsm_output(0));
  and_394_nl <= (fsm_output(6)) AND mux_830_nl;
  or_1085_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_364_cse;
  or_1083_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(7));
  mux_826_nl <= MUX_s_1_2_2(or_1085_nl, or_1083_nl, fsm_output(4));
  or_1082_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (fsm_output(7)));
  or_1080_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(7));
  mux_825_nl <= MUX_s_1_2_2(or_1082_nl, or_1080_nl, fsm_output(4));
  mux_827_nl <= MUX_s_1_2_2(mux_826_nl, mux_825_nl, fsm_output(0));
  nor_743_nl <= NOT((fsm_output(6)) OR mux_827_nl);
  mux_831_nl <= MUX_s_1_2_2(and_394_nl, nor_743_nl, fsm_output(3));
  nand_490_nl <= NOT((fsm_output(5)) AND mux_831_nl);
  nor_745_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (fsm_output(7))));
  nor_746_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(7)));
  mux_822_nl <= MUX_s_1_2_2(nor_745_nl, nor_746_nl, fsm_output(4));
  or_1074_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7)));
  or_1072_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7));
  mux_821_nl <= MUX_s_1_2_2(or_1074_nl, or_1072_nl, fsm_output(4));
  nor_747_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_821_nl);
  mux_823_nl <= MUX_s_1_2_2(mux_822_nl, nor_747_nl, fsm_output(0));
  nand_96_nl <= NOT((fsm_output(6)) AND mux_823_nl);
  or_1070_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (fsm_output(7)));
  or_1068_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(7));
  mux_819_nl <= MUX_s_1_2_2(or_1070_nl, or_1068_nl, fsm_output(4));
  or_1067_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR mux_818_cse;
  mux_820_nl <= MUX_s_1_2_2(mux_819_nl, or_1067_nl, fsm_output(0));
  or_1071_nl <= (fsm_output(6)) OR mux_820_nl;
  mux_824_nl <= MUX_s_1_2_2(nand_96_nl, or_1071_nl, fsm_output(3));
  or_2264_nl <= (fsm_output(5)) OR mux_824_nl;
  mux_832_nl <= MUX_s_1_2_2(nand_490_nl, or_2264_nl, fsm_output(2));
  vec_rsc_0_16_i_we_d_pff <= NOT(mux_832_nl OR (fsm_output(1)));
  nor_732_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_733_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_846_nl <= MUX_s_1_2_2(nor_732_nl, nor_733_nl, fsm_output(0));
  nor_734_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_844_cse);
  nor_735_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_736_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_737_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_840_nl <= MUX_s_1_2_2(nor_736_nl, nor_737_nl, fsm_output(4));
  mux_841_nl <= MUX_s_1_2_2(nor_735_nl, mux_840_nl, fsm_output(3));
  mux_845_nl <= MUX_s_1_2_2(nor_734_nl, mux_841_nl, fsm_output(0));
  mux_847_nl <= MUX_s_1_2_2(mux_846_nl, mux_845_nl, fsm_output(5));
  or_1104_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1102_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_837_nl <= MUX_s_1_2_2(or_1104_nl, or_1102_nl, fsm_output(4));
  or_1101_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1099_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_836_nl <= MUX_s_1_2_2(or_1101_nl, or_1099_nl, fsm_output(4));
  mux_838_nl <= MUX_s_1_2_2(mux_837_nl, mux_836_nl, fsm_output(3));
  or_1098_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR nand_443_cse;
  or_1096_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_834_nl <= MUX_s_1_2_2(or_1098_nl, or_1096_nl, fsm_output(4));
  or_1095_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1093_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_833_nl <= MUX_s_1_2_2(or_1095_nl, or_1093_nl, fsm_output(4));
  mux_835_nl <= MUX_s_1_2_2(mux_834_nl, mux_833_nl, fsm_output(3));
  mux_839_nl <= MUX_s_1_2_2(mux_838_nl, mux_835_nl, fsm_output(0));
  nor_738_nl <= NOT((fsm_output(5)) OR mux_839_nl);
  mux_848_nl <= MUX_s_1_2_2(mux_847_nl, nor_738_nl, fsm_output(2));
  vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_848_nl AND (fsm_output(1));
  nor_720_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))
      OR nand_357_cse);
  nor_721_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (fsm_output(7)));
  mux_860_nl <= MUX_s_1_2_2(nor_720_nl, nor_721_nl, fsm_output(4));
  nor_722_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"))
      OR nand_446_cse);
  nor_723_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (fsm_output(7)));
  mux_859_nl <= MUX_s_1_2_2(nor_722_nl, nor_723_nl, fsm_output(4));
  mux_861_nl <= MUX_s_1_2_2(mux_860_nl, mux_859_nl, fsm_output(0));
  and_391_nl <= (fsm_output(6)) AND mux_861_nl;
  or_1136_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR nand_364_cse;
  or_1134_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (fsm_output(7));
  mux_857_nl <= MUX_s_1_2_2(or_1136_nl, or_1134_nl, fsm_output(4));
  or_1133_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"))
      OR nand_447_cse;
  or_1131_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (fsm_output(7));
  mux_856_nl <= MUX_s_1_2_2(or_1133_nl, or_1131_nl, fsm_output(4));
  mux_858_nl <= MUX_s_1_2_2(mux_857_nl, mux_856_nl, fsm_output(0));
  nor_724_nl <= NOT((fsm_output(6)) OR mux_858_nl);
  mux_862_nl <= MUX_s_1_2_2(and_391_nl, nor_724_nl, fsm_output(3));
  nand_489_nl <= NOT((fsm_output(5)) AND mux_862_nl);
  nor_726_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"))
      OR nand_448_cse);
  nor_727_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (fsm_output(7)));
  mux_853_nl <= MUX_s_1_2_2(nor_726_nl, nor_727_nl, fsm_output(4));
  nor_728_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(7))));
  nor_729_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(7)));
  mux_852_nl <= MUX_s_1_2_2(nor_728_nl, nor_729_nl, fsm_output(4));
  and_392_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_852_nl;
  mux_854_nl <= MUX_s_1_2_2(mux_853_nl, and_392_nl, fsm_output(0));
  nand_102_nl <= NOT((fsm_output(6)) AND mux_854_nl);
  or_1122_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT (fsm_output(7)));
  or_1120_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (fsm_output(7));
  mux_850_nl <= MUX_s_1_2_2(or_1122_nl, or_1120_nl, fsm_output(4));
  nand_100_nl <= NOT(nor_98_cse AND mux_849_cse);
  mux_851_nl <= MUX_s_1_2_2(mux_850_nl, nand_100_nl, fsm_output(0));
  or_1123_nl <= (fsm_output(6)) OR mux_851_nl;
  mux_855_nl <= MUX_s_1_2_2(nand_102_nl, or_1123_nl, fsm_output(3));
  or_2263_nl <= (fsm_output(5)) OR mux_855_nl;
  mux_863_nl <= MUX_s_1_2_2(nand_489_nl, or_2263_nl, fsm_output(2));
  vec_rsc_0_17_i_we_d_pff <= NOT(mux_863_nl OR (fsm_output(1)));
  nor_714_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_715_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_877_nl <= MUX_s_1_2_2(nor_714_nl, nor_715_nl, fsm_output(0));
  and_389_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_844_cse);
  nor_716_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_717_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_718_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_871_nl <= MUX_s_1_2_2(nor_717_nl, nor_718_nl, fsm_output(4));
  mux_872_nl <= MUX_s_1_2_2(nor_716_nl, mux_871_nl, fsm_output(3));
  mux_876_nl <= MUX_s_1_2_2(and_389_nl, mux_872_nl, fsm_output(0));
  mux_878_nl <= MUX_s_1_2_2(mux_877_nl, mux_876_nl, fsm_output(5));
  or_1155_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1153_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_868_nl <= MUX_s_1_2_2(or_1155_nl, or_1153_nl, fsm_output(4));
  or_1152_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1150_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_867_nl <= MUX_s_1_2_2(or_1152_nl, or_1150_nl, fsm_output(4));
  mux_869_nl <= MUX_s_1_2_2(mux_868_nl, mux_867_nl, fsm_output(3));
  or_1149_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))
      OR nand_356_cse;
  or_1147_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_865_nl <= MUX_s_1_2_2(or_1149_nl, or_1147_nl, fsm_output(4));
  or_1146_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1144_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_864_nl <= MUX_s_1_2_2(or_1146_nl, or_1144_nl, fsm_output(4));
  mux_866_nl <= MUX_s_1_2_2(mux_865_nl, mux_864_nl, fsm_output(3));
  mux_870_nl <= MUX_s_1_2_2(mux_869_nl, mux_866_nl, fsm_output(0));
  nor_719_nl <= NOT((fsm_output(5)) OR mux_870_nl);
  mux_879_nl <= MUX_s_1_2_2(mux_878_nl, nor_719_nl, fsm_output(2));
  vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_879_nl AND (fsm_output(1));
  nor_705_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(7))));
  nor_706_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(7)));
  mux_891_nl <= MUX_s_1_2_2(nor_705_nl, nor_706_nl, fsm_output(4));
  nor_707_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(7))));
  nor_708_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(7)));
  mux_890_nl <= MUX_s_1_2_2(nor_707_nl, nor_708_nl, fsm_output(4));
  mux_892_nl <= MUX_s_1_2_2(mux_891_nl, mux_890_nl, fsm_output(0));
  and_388_nl <= (fsm_output(6)) AND mux_892_nl;
  or_1189_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_364_cse;
  or_1187_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(7));
  mux_888_nl <= MUX_s_1_2_2(or_1189_nl, or_1187_nl, fsm_output(4));
  or_1186_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(7)));
  or_1184_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(7));
  mux_887_nl <= MUX_s_1_2_2(or_1186_nl, or_1184_nl, fsm_output(4));
  mux_889_nl <= MUX_s_1_2_2(mux_888_nl, mux_887_nl, fsm_output(0));
  nor_709_nl <= NOT((fsm_output(6)) OR mux_889_nl);
  mux_893_nl <= MUX_s_1_2_2(and_388_nl, nor_709_nl, fsm_output(3));
  nand_488_nl <= NOT((fsm_output(5)) AND mux_893_nl);
  nor_711_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(7))));
  nor_712_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(7)));
  mux_884_nl <= MUX_s_1_2_2(nor_711_nl, nor_712_nl, fsm_output(4));
  or_1178_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100"))
      OR nand_441_cse;
  or_1176_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7));
  mux_883_nl <= MUX_s_1_2_2(or_1178_nl, or_1176_nl, fsm_output(4));
  nor_713_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_883_nl);
  mux_885_nl <= MUX_s_1_2_2(mux_884_nl, nor_713_nl, fsm_output(0));
  nand_107_nl <= NOT((fsm_output(6)) AND mux_885_nl);
  or_1174_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) OR nand_353_cse;
  or_1172_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(7));
  mux_881_nl <= MUX_s_1_2_2(or_1174_nl, or_1172_nl, fsm_output(4));
  or_1171_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR mux_818_cse;
  mux_882_nl <= MUX_s_1_2_2(mux_881_nl, or_1171_nl, fsm_output(0));
  or_1175_nl <= (fsm_output(6)) OR mux_882_nl;
  mux_886_nl <= MUX_s_1_2_2(nand_107_nl, or_1175_nl, fsm_output(3));
  or_2262_nl <= (fsm_output(5)) OR mux_886_nl;
  mux_894_nl <= MUX_s_1_2_2(nand_488_nl, or_2262_nl, fsm_output(2));
  vec_rsc_0_18_i_we_d_pff <= NOT(mux_894_nl OR (fsm_output(1)));
  nor_698_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_699_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_908_nl <= MUX_s_1_2_2(nor_698_nl, nor_699_nl, fsm_output(0));
  nor_700_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_906_cse);
  nor_701_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_702_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_703_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_902_nl <= MUX_s_1_2_2(nor_702_nl, nor_703_nl, fsm_output(4));
  mux_903_nl <= MUX_s_1_2_2(nor_701_nl, mux_902_nl, fsm_output(3));
  mux_907_nl <= MUX_s_1_2_2(nor_700_nl, mux_903_nl, fsm_output(0));
  mux_909_nl <= MUX_s_1_2_2(mux_908_nl, mux_907_nl, fsm_output(5));
  or_1208_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1206_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_899_nl <= MUX_s_1_2_2(or_1208_nl, or_1206_nl, fsm_output(4));
  or_1205_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1203_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_898_nl <= MUX_s_1_2_2(or_1205_nl, or_1203_nl, fsm_output(4));
  mux_900_nl <= MUX_s_1_2_2(mux_899_nl, mux_898_nl, fsm_output(3));
  or_1202_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR nand_443_cse;
  or_1200_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_896_nl <= MUX_s_1_2_2(or_1202_nl, or_1200_nl, fsm_output(4));
  or_1199_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1197_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_895_nl <= MUX_s_1_2_2(or_1199_nl, or_1197_nl, fsm_output(4));
  mux_897_nl <= MUX_s_1_2_2(mux_896_nl, mux_895_nl, fsm_output(3));
  mux_901_nl <= MUX_s_1_2_2(mux_900_nl, mux_897_nl, fsm_output(0));
  nor_704_nl <= NOT((fsm_output(5)) OR mux_901_nl);
  mux_910_nl <= MUX_s_1_2_2(mux_909_nl, nor_704_nl, fsm_output(2));
  vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_910_nl AND (fsm_output(1));
  nor_686_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001"))
      OR nand_357_cse);
  nor_687_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (fsm_output(7)));
  mux_922_nl <= MUX_s_1_2_2(nor_686_nl, nor_687_nl, fsm_output(4));
  nor_688_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("100"))
      OR nand_435_cse);
  nor_689_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (fsm_output(7)));
  mux_921_nl <= MUX_s_1_2_2(nor_688_nl, nor_689_nl, fsm_output(4));
  mux_923_nl <= MUX_s_1_2_2(mux_922_nl, mux_921_nl, fsm_output(0));
  and_385_nl <= (fsm_output(6)) AND mux_923_nl;
  or_1240_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR nand_364_cse;
  or_1238_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (fsm_output(7));
  mux_919_nl <= MUX_s_1_2_2(or_1240_nl, or_1238_nl, fsm_output(4));
  or_1237_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1001"))
      OR nand_447_cse;
  or_1235_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (fsm_output(7));
  mux_918_nl <= MUX_s_1_2_2(or_1237_nl, or_1235_nl, fsm_output(4));
  mux_920_nl <= MUX_s_1_2_2(mux_919_nl, mux_918_nl, fsm_output(0));
  nor_690_nl <= NOT((fsm_output(6)) OR mux_920_nl);
  mux_924_nl <= MUX_s_1_2_2(and_385_nl, nor_690_nl, fsm_output(3));
  nand_487_nl <= NOT((fsm_output(5)) AND mux_924_nl);
  nor_692_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("100"))
      OR nand_437_cse);
  nor_693_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (fsm_output(7)));
  mux_915_nl <= MUX_s_1_2_2(nor_692_nl, nor_693_nl, fsm_output(4));
  nor_694_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100"))
      OR nand_441_cse);
  nor_695_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(7)));
  mux_914_nl <= MUX_s_1_2_2(nor_694_nl, nor_695_nl, fsm_output(4));
  and_386_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_914_nl;
  mux_916_nl <= MUX_s_1_2_2(mux_915_nl, and_386_nl, fsm_output(0));
  nand_113_nl <= NOT((fsm_output(6)) AND mux_916_nl);
  or_1226_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) OR nand_353_cse;
  or_1224_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (fsm_output(7));
  mux_912_nl <= MUX_s_1_2_2(or_1226_nl, or_1224_nl, fsm_output(4));
  nand_111_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_849_cse);
  mux_913_nl <= MUX_s_1_2_2(mux_912_nl, nand_111_nl, fsm_output(0));
  or_1227_nl <= (fsm_output(6)) OR mux_913_nl;
  mux_917_nl <= MUX_s_1_2_2(nand_113_nl, or_1227_nl, fsm_output(3));
  or_2261_nl <= (fsm_output(5)) OR mux_917_nl;
  mux_925_nl <= MUX_s_1_2_2(nand_487_nl, or_2261_nl, fsm_output(2));
  vec_rsc_0_19_i_we_d_pff <= NOT(mux_925_nl OR (fsm_output(1)));
  nor_680_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_681_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_939_nl <= MUX_s_1_2_2(nor_680_nl, nor_681_nl, fsm_output(0));
  and_383_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_906_cse);
  nor_682_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_683_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_684_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_933_nl <= MUX_s_1_2_2(nor_683_nl, nor_684_nl, fsm_output(4));
  mux_934_nl <= MUX_s_1_2_2(nor_682_nl, mux_933_nl, fsm_output(3));
  mux_938_nl <= MUX_s_1_2_2(and_383_nl, mux_934_nl, fsm_output(0));
  mux_940_nl <= MUX_s_1_2_2(mux_939_nl, mux_938_nl, fsm_output(5));
  or_1259_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1257_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_930_nl <= MUX_s_1_2_2(or_1259_nl, or_1257_nl, fsm_output(4));
  or_1256_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1254_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_929_nl <= MUX_s_1_2_2(or_1256_nl, or_1254_nl, fsm_output(4));
  mux_931_nl <= MUX_s_1_2_2(mux_930_nl, mux_929_nl, fsm_output(3));
  or_1253_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001"))
      OR nand_356_cse;
  or_1251_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_927_nl <= MUX_s_1_2_2(or_1253_nl, or_1251_nl, fsm_output(4));
  or_1250_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1248_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_926_nl <= MUX_s_1_2_2(or_1250_nl, or_1248_nl, fsm_output(4));
  mux_928_nl <= MUX_s_1_2_2(mux_927_nl, mux_926_nl, fsm_output(3));
  mux_932_nl <= MUX_s_1_2_2(mux_931_nl, mux_928_nl, fsm_output(0));
  nor_685_nl <= NOT((fsm_output(5)) OR mux_932_nl);
  mux_941_nl <= MUX_s_1_2_2(mux_940_nl, nor_685_nl, fsm_output(2));
  vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_941_nl AND (fsm_output(1));
  nor_671_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (fsm_output(7))));
  nor_672_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(7)));
  mux_953_nl <= MUX_s_1_2_2(nor_671_nl, nor_672_nl, fsm_output(4));
  nor_673_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (fsm_output(7))));
  nor_674_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(7)));
  mux_952_nl <= MUX_s_1_2_2(nor_673_nl, nor_674_nl, fsm_output(4));
  mux_954_nl <= MUX_s_1_2_2(mux_953_nl, mux_952_nl, fsm_output(0));
  and_382_nl <= (fsm_output(6)) AND mux_954_nl;
  or_1293_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_364_cse;
  or_1291_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(7));
  mux_950_nl <= MUX_s_1_2_2(or_1293_nl, or_1291_nl, fsm_output(4));
  or_1290_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (fsm_output(7)));
  or_1288_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(7));
  mux_949_nl <= MUX_s_1_2_2(or_1290_nl, or_1288_nl, fsm_output(4));
  mux_951_nl <= MUX_s_1_2_2(mux_950_nl, mux_949_nl, fsm_output(0));
  nor_675_nl <= NOT((fsm_output(6)) OR mux_951_nl);
  mux_955_nl <= MUX_s_1_2_2(and_382_nl, nor_675_nl, fsm_output(3));
  nand_486_nl <= NOT((fsm_output(5)) AND mux_955_nl);
  nor_677_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (fsm_output(7))));
  nor_678_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(7)));
  mux_946_nl <= MUX_s_1_2_2(nor_677_nl, nor_678_nl, fsm_output(4));
  or_1282_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7)));
  or_1280_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7));
  mux_945_nl <= MUX_s_1_2_2(or_1282_nl, or_1280_nl, fsm_output(4));
  nor_679_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_945_nl);
  mux_947_nl <= MUX_s_1_2_2(mux_946_nl, nor_679_nl, fsm_output(0));
  nand_118_nl <= NOT((fsm_output(6)) AND mux_947_nl);
  or_1278_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (fsm_output(7)));
  or_1276_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(7));
  mux_943_nl <= MUX_s_1_2_2(or_1278_nl, or_1276_nl, fsm_output(4));
  or_1275_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR mux_942_cse;
  mux_944_nl <= MUX_s_1_2_2(mux_943_nl, or_1275_nl, fsm_output(0));
  or_1279_nl <= (fsm_output(6)) OR mux_944_nl;
  mux_948_nl <= MUX_s_1_2_2(nand_118_nl, or_1279_nl, fsm_output(3));
  or_2260_nl <= (fsm_output(5)) OR mux_948_nl;
  mux_956_nl <= MUX_s_1_2_2(nand_486_nl, or_2260_nl, fsm_output(2));
  vec_rsc_0_20_i_we_d_pff <= NOT(mux_956_nl OR (fsm_output(1)));
  nor_664_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_665_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_970_nl <= MUX_s_1_2_2(nor_664_nl, nor_665_nl, fsm_output(0));
  nor_666_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_968_cse);
  nor_667_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_668_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_669_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_964_nl <= MUX_s_1_2_2(nor_668_nl, nor_669_nl, fsm_output(4));
  mux_965_nl <= MUX_s_1_2_2(nor_667_nl, mux_964_nl, fsm_output(3));
  mux_969_nl <= MUX_s_1_2_2(nor_666_nl, mux_965_nl, fsm_output(0));
  mux_971_nl <= MUX_s_1_2_2(mux_970_nl, mux_969_nl, fsm_output(5));
  or_1312_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1310_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_961_nl <= MUX_s_1_2_2(or_1312_nl, or_1310_nl, fsm_output(4));
  or_1309_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1307_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_960_nl <= MUX_s_1_2_2(or_1309_nl, or_1307_nl, fsm_output(4));
  mux_962_nl <= MUX_s_1_2_2(mux_961_nl, mux_960_nl, fsm_output(3));
  or_1306_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR nand_443_cse;
  or_1304_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_958_nl <= MUX_s_1_2_2(or_1306_nl, or_1304_nl, fsm_output(4));
  or_1303_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1301_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_957_nl <= MUX_s_1_2_2(or_1303_nl, or_1301_nl, fsm_output(4));
  mux_959_nl <= MUX_s_1_2_2(mux_958_nl, mux_957_nl, fsm_output(3));
  mux_963_nl <= MUX_s_1_2_2(mux_962_nl, mux_959_nl, fsm_output(0));
  nor_670_nl <= NOT((fsm_output(5)) OR mux_963_nl);
  mux_972_nl <= MUX_s_1_2_2(mux_971_nl, nor_670_nl, fsm_output(2));
  vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_972_nl AND (fsm_output(1));
  nor_652_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"))
      OR nand_357_cse);
  nor_653_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (fsm_output(7)));
  mux_984_nl <= MUX_s_1_2_2(nor_652_nl, nor_653_nl, fsm_output(4));
  nor_654_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"))
      OR nand_446_cse);
  nor_655_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (fsm_output(7)));
  mux_983_nl <= MUX_s_1_2_2(nor_654_nl, nor_655_nl, fsm_output(4));
  mux_985_nl <= MUX_s_1_2_2(mux_984_nl, mux_983_nl, fsm_output(0));
  and_379_nl <= (fsm_output(6)) AND mux_985_nl;
  or_1344_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR nand_364_cse;
  or_1342_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (fsm_output(7));
  mux_981_nl <= MUX_s_1_2_2(or_1344_nl, or_1342_nl, fsm_output(4));
  or_1341_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"))
      OR nand_447_cse;
  or_1339_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (fsm_output(7));
  mux_980_nl <= MUX_s_1_2_2(or_1341_nl, or_1339_nl, fsm_output(4));
  mux_982_nl <= MUX_s_1_2_2(mux_981_nl, mux_980_nl, fsm_output(0));
  nor_656_nl <= NOT((fsm_output(6)) OR mux_982_nl);
  mux_986_nl <= MUX_s_1_2_2(and_379_nl, nor_656_nl, fsm_output(3));
  nand_485_nl <= NOT((fsm_output(5)) AND mux_986_nl);
  nor_658_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"))
      OR nand_448_cse);
  nor_659_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (fsm_output(7)));
  mux_977_nl <= MUX_s_1_2_2(nor_658_nl, nor_659_nl, fsm_output(4));
  nor_660_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(7))));
  nor_661_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(7)));
  mux_976_nl <= MUX_s_1_2_2(nor_660_nl, nor_661_nl, fsm_output(4));
  and_380_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_976_nl;
  mux_978_nl <= MUX_s_1_2_2(mux_977_nl, and_380_nl, fsm_output(0));
  nand_124_nl <= NOT((fsm_output(6)) AND mux_978_nl);
  or_1330_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT (fsm_output(7)));
  or_1328_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (fsm_output(7));
  mux_974_nl <= MUX_s_1_2_2(or_1330_nl, or_1328_nl, fsm_output(4));
  nand_122_nl <= NOT(nor_98_cse AND mux_973_cse);
  mux_975_nl <= MUX_s_1_2_2(mux_974_nl, nand_122_nl, fsm_output(0));
  or_1331_nl <= (fsm_output(6)) OR mux_975_nl;
  mux_979_nl <= MUX_s_1_2_2(nand_124_nl, or_1331_nl, fsm_output(3));
  or_2259_nl <= (fsm_output(5)) OR mux_979_nl;
  mux_987_nl <= MUX_s_1_2_2(nand_485_nl, or_2259_nl, fsm_output(2));
  vec_rsc_0_21_i_we_d_pff <= NOT(mux_987_nl OR (fsm_output(1)));
  nor_646_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_647_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1001_nl <= MUX_s_1_2_2(nor_646_nl, nor_647_nl, fsm_output(0));
  and_377_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_968_cse);
  nor_648_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_649_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_650_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_995_nl <= MUX_s_1_2_2(nor_649_nl, nor_650_nl, fsm_output(4));
  mux_996_nl <= MUX_s_1_2_2(nor_648_nl, mux_995_nl, fsm_output(3));
  mux_1000_nl <= MUX_s_1_2_2(and_377_nl, mux_996_nl, fsm_output(0));
  mux_1002_nl <= MUX_s_1_2_2(mux_1001_nl, mux_1000_nl, fsm_output(5));
  or_1363_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1361_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_992_nl <= MUX_s_1_2_2(or_1363_nl, or_1361_nl, fsm_output(4));
  or_1360_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1358_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_991_nl <= MUX_s_1_2_2(or_1360_nl, or_1358_nl, fsm_output(4));
  mux_993_nl <= MUX_s_1_2_2(mux_992_nl, mux_991_nl, fsm_output(3));
  or_1357_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"))
      OR nand_356_cse;
  or_1355_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_989_nl <= MUX_s_1_2_2(or_1357_nl, or_1355_nl, fsm_output(4));
  or_1354_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1352_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_988_nl <= MUX_s_1_2_2(or_1354_nl, or_1352_nl, fsm_output(4));
  mux_990_nl <= MUX_s_1_2_2(mux_989_nl, mux_988_nl, fsm_output(3));
  mux_994_nl <= MUX_s_1_2_2(mux_993_nl, mux_990_nl, fsm_output(0));
  nor_651_nl <= NOT((fsm_output(5)) OR mux_994_nl);
  mux_1003_nl <= MUX_s_1_2_2(mux_1002_nl, nor_651_nl, fsm_output(2));
  vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1003_nl AND (fsm_output(1));
  nor_637_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(7))));
  nor_638_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(7)));
  mux_1015_nl <= MUX_s_1_2_2(nor_637_nl, nor_638_nl, fsm_output(4));
  nor_639_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(7))));
  nor_640_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(7)));
  mux_1014_nl <= MUX_s_1_2_2(nor_639_nl, nor_640_nl, fsm_output(4));
  mux_1016_nl <= MUX_s_1_2_2(mux_1015_nl, mux_1014_nl, fsm_output(0));
  and_376_nl <= (fsm_output(6)) AND mux_1016_nl;
  or_1397_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_364_cse;
  or_1395_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(7));
  mux_1012_nl <= MUX_s_1_2_2(or_1397_nl, or_1395_nl, fsm_output(4));
  or_1394_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(7)));
  or_1392_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(7));
  mux_1011_nl <= MUX_s_1_2_2(or_1394_nl, or_1392_nl, fsm_output(4));
  mux_1013_nl <= MUX_s_1_2_2(mux_1012_nl, mux_1011_nl, fsm_output(0));
  nor_641_nl <= NOT((fsm_output(6)) OR mux_1013_nl);
  mux_1017_nl <= MUX_s_1_2_2(and_376_nl, nor_641_nl, fsm_output(3));
  nand_484_nl <= NOT((fsm_output(5)) AND mux_1017_nl);
  nor_643_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(7))));
  nor_644_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(7)));
  mux_1008_nl <= MUX_s_1_2_2(nor_643_nl, nor_644_nl, fsm_output(4));
  or_1386_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10"))
      OR nand_423_cse;
  or_1384_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7));
  mux_1007_nl <= MUX_s_1_2_2(or_1386_nl, or_1384_nl, fsm_output(4));
  nor_645_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1007_nl);
  mux_1009_nl <= MUX_s_1_2_2(mux_1008_nl, nor_645_nl, fsm_output(0));
  nand_129_nl <= NOT((fsm_output(6)) AND mux_1009_nl);
  or_1382_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) OR nand_353_cse;
  or_1380_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(7));
  mux_1005_nl <= MUX_s_1_2_2(or_1382_nl, or_1380_nl, fsm_output(4));
  or_1379_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR mux_942_cse;
  mux_1006_nl <= MUX_s_1_2_2(mux_1005_nl, or_1379_nl, fsm_output(0));
  or_1383_nl <= (fsm_output(6)) OR mux_1006_nl;
  mux_1010_nl <= MUX_s_1_2_2(nand_129_nl, or_1383_nl, fsm_output(3));
  or_2258_nl <= (fsm_output(5)) OR mux_1010_nl;
  mux_1018_nl <= MUX_s_1_2_2(nand_484_nl, or_2258_nl, fsm_output(2));
  vec_rsc_0_22_i_we_d_pff <= NOT(mux_1018_nl OR (fsm_output(1)));
  nor_630_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_631_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1032_nl <= MUX_s_1_2_2(nor_630_nl, nor_631_nl, fsm_output(0));
  nor_632_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1030_cse);
  nor_633_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_634_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_635_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1026_nl <= MUX_s_1_2_2(nor_634_nl, nor_635_nl, fsm_output(4));
  mux_1027_nl <= MUX_s_1_2_2(nor_633_nl, mux_1026_nl, fsm_output(3));
  mux_1031_nl <= MUX_s_1_2_2(nor_632_nl, mux_1027_nl, fsm_output(0));
  mux_1033_nl <= MUX_s_1_2_2(mux_1032_nl, mux_1031_nl, fsm_output(5));
  or_1416_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1414_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_1023_nl <= MUX_s_1_2_2(or_1416_nl, or_1414_nl, fsm_output(4));
  or_1413_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1411_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1022_nl <= MUX_s_1_2_2(or_1413_nl, or_1411_nl, fsm_output(4));
  mux_1024_nl <= MUX_s_1_2_2(mux_1023_nl, mux_1022_nl, fsm_output(3));
  or_1410_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR nand_443_cse;
  or_1408_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_1020_nl <= MUX_s_1_2_2(or_1410_nl, or_1408_nl, fsm_output(4));
  or_1407_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1405_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1019_nl <= MUX_s_1_2_2(or_1407_nl, or_1405_nl, fsm_output(4));
  mux_1021_nl <= MUX_s_1_2_2(mux_1020_nl, mux_1019_nl, fsm_output(3));
  mux_1025_nl <= MUX_s_1_2_2(mux_1024_nl, mux_1021_nl, fsm_output(0));
  nor_636_nl <= NOT((fsm_output(5)) OR mux_1025_nl);
  mux_1034_nl <= MUX_s_1_2_2(mux_1033_nl, nor_636_nl, fsm_output(2));
  vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1034_nl AND (fsm_output(1));
  nor_618_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011"))
      OR nand_357_cse);
  nor_619_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (fsm_output(7)));
  mux_1046_nl <= MUX_s_1_2_2(nor_618_nl, nor_619_nl, fsm_output(4));
  nor_620_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10"))
      OR nand_417_cse);
  nor_621_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (fsm_output(7)));
  mux_1045_nl <= MUX_s_1_2_2(nor_620_nl, nor_621_nl, fsm_output(4));
  mux_1047_nl <= MUX_s_1_2_2(mux_1046_nl, mux_1045_nl, fsm_output(0));
  and_373_nl <= (fsm_output(6)) AND mux_1047_nl;
  or_1448_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))))
      OR nand_364_cse;
  or_1446_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (fsm_output(7));
  mux_1043_nl <= MUX_s_1_2_2(or_1448_nl, or_1446_nl, fsm_output(4));
  or_1445_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1011"))))
      OR nand_447_cse;
  or_1443_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (fsm_output(7));
  mux_1042_nl <= MUX_s_1_2_2(or_1445_nl, or_1443_nl, fsm_output(4));
  mux_1044_nl <= MUX_s_1_2_2(mux_1043_nl, mux_1042_nl, fsm_output(0));
  nor_622_nl <= NOT((fsm_output(6)) OR mux_1044_nl);
  mux_1048_nl <= MUX_s_1_2_2(and_373_nl, nor_622_nl, fsm_output(3));
  nand_483_nl <= NOT((fsm_output(5)) AND mux_1048_nl);
  nor_624_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10"))
      OR nand_419_cse);
  nor_625_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (fsm_output(7)));
  mux_1039_nl <= MUX_s_1_2_2(nor_624_nl, nor_625_nl, fsm_output(4));
  nor_626_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10"))
      OR nand_423_cse);
  nor_627_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(7)));
  mux_1038_nl <= MUX_s_1_2_2(nor_626_nl, nor_627_nl, fsm_output(4));
  and_374_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1038_nl;
  mux_1040_nl <= MUX_s_1_2_2(mux_1039_nl, and_374_nl, fsm_output(0));
  nand_135_nl <= NOT((fsm_output(6)) AND mux_1040_nl);
  or_1434_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) OR nand_353_cse;
  or_1432_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (fsm_output(7));
  mux_1036_nl <= MUX_s_1_2_2(or_1434_nl, or_1432_nl, fsm_output(4));
  nand_133_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_973_cse);
  mux_1037_nl <= MUX_s_1_2_2(mux_1036_nl, nand_133_nl, fsm_output(0));
  or_1435_nl <= (fsm_output(6)) OR mux_1037_nl;
  mux_1041_nl <= MUX_s_1_2_2(nand_135_nl, or_1435_nl, fsm_output(3));
  or_2257_nl <= (fsm_output(5)) OR mux_1041_nl;
  mux_1049_nl <= MUX_s_1_2_2(nand_483_nl, or_2257_nl, fsm_output(2));
  vec_rsc_0_23_i_we_d_pff <= NOT(mux_1049_nl OR (fsm_output(1)));
  nor_613_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_614_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1063_nl <= MUX_s_1_2_2(nor_613_nl, nor_614_nl, fsm_output(0));
  and_370_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_1030_cse);
  and_371_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND (fsm_output(4)) AND (fsm_output(6)) AND (NOT (fsm_output(7)));
  and_526_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  nor_616_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1057_nl <= MUX_s_1_2_2(and_526_nl, nor_616_nl, fsm_output(4));
  mux_1058_nl <= MUX_s_1_2_2(and_371_nl, mux_1057_nl, fsm_output(3));
  mux_1062_nl <= MUX_s_1_2_2(and_370_nl, mux_1058_nl, fsm_output(0));
  mux_1064_nl <= MUX_s_1_2_2(mux_1063_nl, mux_1062_nl, fsm_output(5));
  or_1467_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)) OR nand_443_cse;
  nand_307_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("01")));
  mux_1054_nl <= MUX_s_1_2_2(or_1467_nl, nand_307_nl, fsm_output(4));
  nand_514_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1462_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1053_nl <= MUX_s_1_2_2(nand_514_nl, or_1462_nl, fsm_output(4));
  mux_1055_nl <= MUX_s_1_2_2(mux_1054_nl, mux_1053_nl, fsm_output(3));
  or_1461_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011"))
      OR nand_356_cse;
  nand_310_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_1051_nl <= MUX_s_1_2_2(or_1461_nl, nand_310_nl, fsm_output(4));
  nand_468_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  or_1456_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1050_nl <= MUX_s_1_2_2(nand_468_nl, or_1456_nl, fsm_output(4));
  mux_1052_nl <= MUX_s_1_2_2(mux_1051_nl, mux_1050_nl, fsm_output(3));
  mux_1056_nl <= MUX_s_1_2_2(mux_1055_nl, mux_1052_nl, fsm_output(0));
  nor_617_nl <= NOT((fsm_output(5)) OR mux_1056_nl);
  mux_1065_nl <= MUX_s_1_2_2(mux_1064_nl, nor_617_nl, fsm_output(2));
  vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1065_nl AND (fsm_output(1));
  nor_604_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (fsm_output(7))));
  nor_605_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(7)));
  mux_1077_nl <= MUX_s_1_2_2(nor_604_nl, nor_605_nl, fsm_output(4));
  nor_606_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (fsm_output(7))));
  nor_607_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(7)));
  mux_1076_nl <= MUX_s_1_2_2(nor_606_nl, nor_607_nl, fsm_output(4));
  mux_1078_nl <= MUX_s_1_2_2(mux_1077_nl, mux_1076_nl, fsm_output(0));
  and_369_nl <= (fsm_output(6)) AND mux_1078_nl;
  or_1500_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_302_cse;
  or_1498_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(7));
  mux_1074_nl <= MUX_s_1_2_2(or_1500_nl, or_1498_nl, fsm_output(4));
  or_1497_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (fsm_output(7)));
  or_1495_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(7));
  mux_1073_nl <= MUX_s_1_2_2(or_1497_nl, or_1495_nl, fsm_output(4));
  mux_1075_nl <= MUX_s_1_2_2(mux_1074_nl, mux_1073_nl, fsm_output(0));
  nor_608_nl <= NOT((fsm_output(6)) OR mux_1075_nl);
  mux_1079_nl <= MUX_s_1_2_2(and_369_nl, nor_608_nl, fsm_output(3));
  nand_482_nl <= NOT((fsm_output(5)) AND mux_1079_nl);
  nor_610_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (fsm_output(7))));
  nor_611_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(7)));
  mux_1070_nl <= MUX_s_1_2_2(nor_610_nl, nor_611_nl, fsm_output(4));
  or_1489_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7)));
  or_1487_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7));
  mux_1069_nl <= MUX_s_1_2_2(or_1489_nl, or_1487_nl, fsm_output(4));
  nor_612_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1069_nl);
  mux_1071_nl <= MUX_s_1_2_2(mux_1070_nl, nor_612_nl, fsm_output(0));
  nand_140_nl <= NOT((fsm_output(6)) AND mux_1071_nl);
  or_1485_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (fsm_output(7)));
  or_1483_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(7));
  mux_1067_nl <= MUX_s_1_2_2(or_1485_nl, or_1483_nl, fsm_output(4));
  or_1482_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1066_cse;
  mux_1068_nl <= MUX_s_1_2_2(mux_1067_nl, or_1482_nl, fsm_output(0));
  or_1486_nl <= (fsm_output(6)) OR mux_1068_nl;
  mux_1072_nl <= MUX_s_1_2_2(nand_140_nl, or_1486_nl, fsm_output(3));
  or_2256_nl <= (fsm_output(5)) OR mux_1072_nl;
  mux_1080_nl <= MUX_s_1_2_2(nand_482_nl, or_2256_nl, fsm_output(2));
  vec_rsc_0_24_i_we_d_pff <= NOT(mux_1080_nl OR (fsm_output(1)));
  nor_597_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_598_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1094_nl <= MUX_s_1_2_2(nor_597_nl, nor_598_nl, fsm_output(0));
  nor_599_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1092_cse);
  nor_600_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_601_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_602_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1088_nl <= MUX_s_1_2_2(nor_601_nl, nor_602_nl, fsm_output(4));
  mux_1089_nl <= MUX_s_1_2_2(nor_600_nl, mux_1088_nl, fsm_output(3));
  mux_1093_nl <= MUX_s_1_2_2(nor_599_nl, mux_1089_nl, fsm_output(0));
  mux_1095_nl <= MUX_s_1_2_2(mux_1094_nl, mux_1093_nl, fsm_output(5));
  or_1519_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1517_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_1085_nl <= MUX_s_1_2_2(or_1519_nl, or_1517_nl, fsm_output(4));
  or_1516_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1514_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1084_nl <= MUX_s_1_2_2(or_1516_nl, or_1514_nl, fsm_output(4));
  mux_1086_nl <= MUX_s_1_2_2(mux_1085_nl, mux_1084_nl, fsm_output(3));
  or_1513_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR nand_443_cse;
  or_1511_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_1082_nl <= MUX_s_1_2_2(or_1513_nl, or_1511_nl, fsm_output(4));
  or_1510_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1508_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1081_nl <= MUX_s_1_2_2(or_1510_nl, or_1508_nl, fsm_output(4));
  mux_1083_nl <= MUX_s_1_2_2(mux_1082_nl, mux_1081_nl, fsm_output(3));
  mux_1087_nl <= MUX_s_1_2_2(mux_1086_nl, mux_1083_nl, fsm_output(0));
  nor_603_nl <= NOT((fsm_output(5)) OR mux_1087_nl);
  mux_1096_nl <= MUX_s_1_2_2(mux_1095_nl, nor_603_nl, fsm_output(2));
  vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1096_nl AND (fsm_output(1));
  nor_585_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR nand_294_cse);
  nor_586_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (fsm_output(7)));
  mux_1108_nl <= MUX_s_1_2_2(nor_585_nl, nor_586_nl, fsm_output(4));
  nor_587_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100"))
      OR nand_446_cse);
  nor_588_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (fsm_output(7)));
  mux_1107_nl <= MUX_s_1_2_2(nor_587_nl, nor_588_nl, fsm_output(4));
  mux_1109_nl <= MUX_s_1_2_2(mux_1108_nl, mux_1107_nl, fsm_output(0));
  and_366_nl <= (fsm_output(6)) AND mux_1109_nl;
  or_1550_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_302_cse;
  or_1548_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (fsm_output(7));
  mux_1105_nl <= MUX_s_1_2_2(or_1550_nl, or_1548_nl, fsm_output(4));
  or_1547_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR nand_297_cse;
  or_1545_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (fsm_output(7));
  mux_1104_nl <= MUX_s_1_2_2(or_1547_nl, or_1545_nl, fsm_output(4));
  mux_1106_nl <= MUX_s_1_2_2(mux_1105_nl, mux_1104_nl, fsm_output(0));
  nor_589_nl <= NOT((fsm_output(6)) OR mux_1106_nl);
  mux_1110_nl <= MUX_s_1_2_2(and_366_nl, nor_589_nl, fsm_output(3));
  nand_481_nl <= NOT((fsm_output(5)) AND mux_1110_nl);
  nor_591_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100"))
      OR nand_448_cse);
  nor_592_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (fsm_output(7)));
  mux_1101_nl <= MUX_s_1_2_2(nor_591_nl, nor_592_nl, fsm_output(4));
  nor_593_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(7))));
  nor_594_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(7)));
  mux_1100_nl <= MUX_s_1_2_2(nor_593_nl, nor_594_nl, fsm_output(4));
  and_367_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1100_nl;
  mux_1102_nl <= MUX_s_1_2_2(mux_1101_nl, and_367_nl, fsm_output(0));
  nand_146_nl <= NOT((fsm_output(6)) AND mux_1102_nl);
  or_1536_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT (fsm_output(7)));
  or_1534_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (fsm_output(7));
  mux_1098_nl <= MUX_s_1_2_2(or_1536_nl, or_1534_nl, fsm_output(4));
  nand_144_nl <= NOT(nor_98_cse AND mux_1097_cse);
  mux_1099_nl <= MUX_s_1_2_2(mux_1098_nl, nand_144_nl, fsm_output(0));
  or_1537_nl <= (fsm_output(6)) OR mux_1099_nl;
  mux_1103_nl <= MUX_s_1_2_2(nand_146_nl, or_1537_nl, fsm_output(3));
  or_2255_nl <= (fsm_output(5)) OR mux_1103_nl;
  mux_1111_nl <= MUX_s_1_2_2(nand_481_nl, or_2255_nl, fsm_output(2));
  vec_rsc_0_25_i_we_d_pff <= NOT(mux_1111_nl OR (fsm_output(1)));
  nor_579_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_580_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1125_nl <= MUX_s_1_2_2(nor_579_nl, nor_580_nl, fsm_output(0));
  and_364_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_1092_cse);
  nor_581_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_582_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_583_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1119_nl <= MUX_s_1_2_2(nor_582_nl, nor_583_nl, fsm_output(4));
  mux_1120_nl <= MUX_s_1_2_2(nor_581_nl, mux_1119_nl, fsm_output(3));
  mux_1124_nl <= MUX_s_1_2_2(and_364_nl, mux_1120_nl, fsm_output(0));
  mux_1126_nl <= MUX_s_1_2_2(mux_1125_nl, mux_1124_nl, fsm_output(5));
  or_1569_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1567_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_1116_nl <= MUX_s_1_2_2(or_1569_nl, or_1567_nl, fsm_output(4));
  or_1566_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1564_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1115_nl <= MUX_s_1_2_2(or_1566_nl, or_1564_nl, fsm_output(4));
  mux_1117_nl <= MUX_s_1_2_2(mux_1116_nl, mux_1115_nl, fsm_output(3));
  or_1563_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR nand_293_cse;
  or_1561_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_1113_nl <= MUX_s_1_2_2(or_1563_nl, or_1561_nl, fsm_output(4));
  or_1560_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1558_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1112_nl <= MUX_s_1_2_2(or_1560_nl, or_1558_nl, fsm_output(4));
  mux_1114_nl <= MUX_s_1_2_2(mux_1113_nl, mux_1112_nl, fsm_output(3));
  mux_1118_nl <= MUX_s_1_2_2(mux_1117_nl, mux_1114_nl, fsm_output(0));
  nor_584_nl <= NOT((fsm_output(5)) OR mux_1118_nl);
  mux_1127_nl <= MUX_s_1_2_2(mux_1126_nl, nor_584_nl, fsm_output(2));
  vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1127_nl AND (fsm_output(1));
  nor_570_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(7))));
  nor_571_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(7)));
  mux_1139_nl <= MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output(4));
  nor_572_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(7))));
  nor_573_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(7)));
  mux_1138_nl <= MUX_s_1_2_2(nor_572_nl, nor_573_nl, fsm_output(4));
  mux_1140_nl <= MUX_s_1_2_2(mux_1139_nl, mux_1138_nl, fsm_output(0));
  and_363_nl <= (fsm_output(6)) AND mux_1140_nl;
  or_1602_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_302_cse;
  or_1600_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(7));
  mux_1136_nl <= MUX_s_1_2_2(or_1602_nl, or_1600_nl, fsm_output(4));
  or_1599_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(7)));
  or_1597_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(7));
  mux_1135_nl <= MUX_s_1_2_2(or_1599_nl, or_1597_nl, fsm_output(4));
  mux_1137_nl <= MUX_s_1_2_2(mux_1136_nl, mux_1135_nl, fsm_output(0));
  nor_574_nl <= NOT((fsm_output(6)) OR mux_1137_nl);
  mux_1141_nl <= MUX_s_1_2_2(and_363_nl, nor_574_nl, fsm_output(3));
  nand_480_nl <= NOT((fsm_output(5)) AND mux_1141_nl);
  nor_576_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(7))));
  nor_577_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(7)));
  mux_1132_nl <= MUX_s_1_2_2(nor_576_nl, nor_577_nl, fsm_output(4));
  or_1591_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110"))
      OR nand_441_cse;
  or_1589_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7));
  mux_1131_nl <= MUX_s_1_2_2(or_1591_nl, or_1589_nl, fsm_output(4));
  nor_578_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1131_nl);
  mux_1133_nl <= MUX_s_1_2_2(mux_1132_nl, nor_578_nl, fsm_output(0));
  nand_151_nl <= NOT((fsm_output(6)) AND mux_1133_nl);
  or_1587_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR nand_289_cse;
  or_1585_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(7));
  mux_1129_nl <= MUX_s_1_2_2(or_1587_nl, or_1585_nl, fsm_output(4));
  or_1584_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1066_cse;
  mux_1130_nl <= MUX_s_1_2_2(mux_1129_nl, or_1584_nl, fsm_output(0));
  or_1588_nl <= (fsm_output(6)) OR mux_1130_nl;
  mux_1134_nl <= MUX_s_1_2_2(nand_151_nl, or_1588_nl, fsm_output(3));
  or_2254_nl <= (fsm_output(5)) OR mux_1134_nl;
  mux_1142_nl <= MUX_s_1_2_2(nand_480_nl, or_2254_nl, fsm_output(2));
  vec_rsc_0_26_i_we_d_pff <= NOT(mux_1142_nl OR (fsm_output(1)));
  nor_563_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_564_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1156_nl <= MUX_s_1_2_2(nor_563_nl, nor_564_nl, fsm_output(0));
  nor_565_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1154_cse);
  nor_566_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_567_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_568_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1150_nl <= MUX_s_1_2_2(nor_567_nl, nor_568_nl, fsm_output(4));
  mux_1151_nl <= MUX_s_1_2_2(nor_566_nl, mux_1150_nl, fsm_output(3));
  mux_1155_nl <= MUX_s_1_2_2(nor_565_nl, mux_1151_nl, fsm_output(0));
  mux_1157_nl <= MUX_s_1_2_2(mux_1156_nl, mux_1155_nl, fsm_output(5));
  or_1621_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1619_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_1147_nl <= MUX_s_1_2_2(or_1621_nl, or_1619_nl, fsm_output(4));
  or_1618_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1616_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1146_nl <= MUX_s_1_2_2(or_1618_nl, or_1616_nl, fsm_output(4));
  mux_1148_nl <= MUX_s_1_2_2(mux_1147_nl, mux_1146_nl, fsm_output(3));
  or_1615_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR nand_443_cse;
  or_1613_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_1144_nl <= MUX_s_1_2_2(or_1615_nl, or_1613_nl, fsm_output(4));
  or_1612_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1610_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1143_nl <= MUX_s_1_2_2(or_1612_nl, or_1610_nl, fsm_output(4));
  mux_1145_nl <= MUX_s_1_2_2(mux_1144_nl, mux_1143_nl, fsm_output(3));
  mux_1149_nl <= MUX_s_1_2_2(mux_1148_nl, mux_1145_nl, fsm_output(0));
  nor_569_nl <= NOT((fsm_output(5)) OR mux_1149_nl);
  mux_1158_nl <= MUX_s_1_2_2(mux_1157_nl, nor_569_nl, fsm_output(2));
  vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1158_nl AND (fsm_output(1));
  nor_551_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"))
      OR nand_294_cse);
  nor_552_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (fsm_output(7)));
  mux_1170_nl <= MUX_s_1_2_2(nor_551_nl, nor_552_nl, fsm_output(4));
  nor_553_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("110"))
      OR nand_435_cse);
  nor_554_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (fsm_output(7)));
  mux_1169_nl <= MUX_s_1_2_2(nor_553_nl, nor_554_nl, fsm_output(4));
  mux_1171_nl <= MUX_s_1_2_2(mux_1170_nl, mux_1169_nl, fsm_output(0));
  and_360_nl <= (fsm_output(6)) AND mux_1171_nl;
  or_1651_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR nand_302_cse;
  or_1649_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (fsm_output(7));
  mux_1167_nl <= MUX_s_1_2_2(or_1651_nl, or_1649_nl, fsm_output(4));
  or_1648_nl <= (COMP_LOOP_acc_1_cse_6_sva(2)) OR (NOT((COMP_LOOP_acc_1_cse_6_sva(1))
      AND (COMP_LOOP_acc_1_cse_6_sva(4)) AND (COMP_LOOP_acc_1_cse_6_sva(3)) AND (COMP_LOOP_acc_1_cse_6_sva(0))
      AND (fsm_output(7))));
  or_1647_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (fsm_output(7));
  mux_1166_nl <= MUX_s_1_2_2(or_1648_nl, or_1647_nl, fsm_output(4));
  mux_1168_nl <= MUX_s_1_2_2(mux_1167_nl, mux_1166_nl, fsm_output(0));
  nor_555_nl <= NOT((fsm_output(6)) OR mux_1168_nl);
  mux_1172_nl <= MUX_s_1_2_2(and_360_nl, nor_555_nl, fsm_output(3));
  nand_479_nl <= NOT((fsm_output(5)) AND mux_1172_nl);
  nor_557_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("110"))
      OR nand_437_cse);
  nor_558_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (fsm_output(7)));
  mux_1163_nl <= MUX_s_1_2_2(nor_557_nl, nor_558_nl, fsm_output(4));
  nor_559_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("110"))
      OR nand_441_cse);
  nor_560_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(7)));
  mux_1162_nl <= MUX_s_1_2_2(nor_559_nl, nor_560_nl, fsm_output(4));
  and_361_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1162_nl;
  mux_1164_nl <= MUX_s_1_2_2(mux_1163_nl, and_361_nl, fsm_output(0));
  nand_157_nl <= NOT((fsm_output(6)) AND mux_1164_nl);
  or_1638_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR nand_289_cse;
  or_1636_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (fsm_output(7));
  mux_1160_nl <= MUX_s_1_2_2(or_1638_nl, or_1636_nl, fsm_output(4));
  nand_155_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_1097_cse);
  mux_1161_nl <= MUX_s_1_2_2(mux_1160_nl, nand_155_nl, fsm_output(0));
  or_1639_nl <= (fsm_output(6)) OR mux_1161_nl;
  mux_1165_nl <= MUX_s_1_2_2(nand_157_nl, or_1639_nl, fsm_output(3));
  or_2253_nl <= (fsm_output(5)) OR mux_1165_nl;
  mux_1173_nl <= MUX_s_1_2_2(nand_479_nl, or_2253_nl, fsm_output(2));
  vec_rsc_0_27_i_we_d_pff <= NOT(mux_1173_nl OR (fsm_output(1)));
  nor_546_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_547_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1187_nl <= MUX_s_1_2_2(nor_546_nl, nor_547_nl, fsm_output(0));
  and_357_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_1154_cse);
  and_358_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND (fsm_output(4)) AND (fsm_output(6)) AND (NOT (fsm_output(7)));
  and_525_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  nor_549_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1181_nl <= MUX_s_1_2_2(and_525_nl, nor_549_nl, fsm_output(4));
  mux_1182_nl <= MUX_s_1_2_2(and_358_nl, mux_1181_nl, fsm_output(3));
  mux_1186_nl <= MUX_s_1_2_2(and_357_nl, mux_1182_nl, fsm_output(0));
  mux_1188_nl <= MUX_s_1_2_2(mux_1187_nl, mux_1186_nl, fsm_output(5));
  or_1670_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)) OR nand_443_cse;
  nand_273_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("01")));
  mux_1178_nl <= MUX_s_1_2_2(or_1670_nl, nand_273_nl, fsm_output(4));
  nand_513_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1665_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1177_nl <= MUX_s_1_2_2(nand_513_nl, or_1665_nl, fsm_output(4));
  mux_1179_nl <= MUX_s_1_2_2(mux_1178_nl, mux_1177_nl, fsm_output(3));
  or_1664_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"))
      OR nand_293_cse;
  nand_276_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_1175_nl <= MUX_s_1_2_2(or_1664_nl, nand_276_nl, fsm_output(4));
  nand_465_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  or_1659_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1174_nl <= MUX_s_1_2_2(nand_465_nl, or_1659_nl, fsm_output(4));
  mux_1176_nl <= MUX_s_1_2_2(mux_1175_nl, mux_1174_nl, fsm_output(3));
  mux_1180_nl <= MUX_s_1_2_2(mux_1179_nl, mux_1176_nl, fsm_output(0));
  nor_550_nl <= NOT((fsm_output(5)) OR mux_1180_nl);
  mux_1189_nl <= MUX_s_1_2_2(mux_1188_nl, nor_550_nl, fsm_output(2));
  vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1189_nl AND (fsm_output(1));
  nor_537_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (fsm_output(7))));
  nor_538_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(7)));
  mux_1201_nl <= MUX_s_1_2_2(nor_537_nl, nor_538_nl, fsm_output(4));
  nor_539_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (fsm_output(7))));
  nor_540_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(7)));
  mux_1200_nl <= MUX_s_1_2_2(nor_539_nl, nor_540_nl, fsm_output(4));
  mux_1202_nl <= MUX_s_1_2_2(mux_1201_nl, mux_1200_nl, fsm_output(0));
  and_356_nl <= (fsm_output(6)) AND mux_1202_nl;
  or_1702_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_266_cse;
  or_1700_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(7));
  mux_1198_nl <= MUX_s_1_2_2(or_1702_nl, or_1700_nl, fsm_output(4));
  or_1699_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (fsm_output(7)));
  or_1697_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(7));
  mux_1197_nl <= MUX_s_1_2_2(or_1699_nl, or_1697_nl, fsm_output(4));
  mux_1199_nl <= MUX_s_1_2_2(mux_1198_nl, mux_1197_nl, fsm_output(0));
  nor_541_nl <= NOT((fsm_output(6)) OR mux_1199_nl);
  mux_1203_nl <= MUX_s_1_2_2(and_356_nl, nor_541_nl, fsm_output(3));
  nand_478_nl <= NOT((fsm_output(5)) AND mux_1203_nl);
  nor_543_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (fsm_output(7))));
  nor_544_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(7)));
  mux_1194_nl <= MUX_s_1_2_2(nor_543_nl, nor_544_nl, fsm_output(4));
  nand_519_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(7)));
  or_1689_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7));
  mux_1193_nl <= MUX_s_1_2_2(nand_519_nl, or_1689_nl, fsm_output(4));
  nor_545_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1193_nl);
  mux_1195_nl <= MUX_s_1_2_2(mux_1194_nl, nor_545_nl, fsm_output(0));
  nand_162_nl <= NOT((fsm_output(6)) AND mux_1195_nl);
  or_1687_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (fsm_output(7)));
  or_1685_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(7));
  mux_1191_nl <= MUX_s_1_2_2(or_1687_nl, or_1685_nl, fsm_output(4));
  or_1684_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1190_cse;
  mux_1192_nl <= MUX_s_1_2_2(mux_1191_nl, or_1684_nl, fsm_output(0));
  or_1688_nl <= (fsm_output(6)) OR mux_1192_nl;
  mux_1196_nl <= MUX_s_1_2_2(nand_162_nl, or_1688_nl, fsm_output(3));
  or_2252_nl <= (fsm_output(5)) OR mux_1196_nl;
  mux_1204_nl <= MUX_s_1_2_2(nand_478_nl, or_2252_nl, fsm_output(2));
  vec_rsc_0_28_i_we_d_pff <= NOT(mux_1204_nl OR (fsm_output(1)));
  nor_530_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_531_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1218_nl <= MUX_s_1_2_2(nor_530_nl, nor_531_nl, fsm_output(0));
  nor_532_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1216_cse);
  nor_533_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(6))) OR (fsm_output(7)));
  nor_534_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  nor_535_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1212_nl <= MUX_s_1_2_2(nor_534_nl, nor_535_nl, fsm_output(4));
  mux_1213_nl <= MUX_s_1_2_2(nor_533_nl, mux_1212_nl, fsm_output(3));
  mux_1217_nl <= MUX_s_1_2_2(nor_532_nl, mux_1213_nl, fsm_output(0));
  mux_1219_nl <= MUX_s_1_2_2(mux_1218_nl, mux_1217_nl, fsm_output(5));
  or_1721_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR nand_443_cse;
  or_1719_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_1209_nl <= MUX_s_1_2_2(or_1721_nl, or_1719_nl, fsm_output(4));
  or_1718_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("10"));
  or_1716_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1208_nl <= MUX_s_1_2_2(or_1718_nl, or_1716_nl, fsm_output(4));
  mux_1210_nl <= MUX_s_1_2_2(mux_1209_nl, mux_1208_nl, fsm_output(3));
  or_1715_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR nand_443_cse;
  or_1713_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_1206_nl <= MUX_s_1_2_2(or_1715_nl, or_1713_nl, fsm_output(4));
  or_1712_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1710_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1205_nl <= MUX_s_1_2_2(or_1712_nl, or_1710_nl, fsm_output(4));
  mux_1207_nl <= MUX_s_1_2_2(mux_1206_nl, mux_1205_nl, fsm_output(3));
  mux_1211_nl <= MUX_s_1_2_2(mux_1210_nl, mux_1207_nl, fsm_output(0));
  nor_536_nl <= NOT((fsm_output(5)) OR mux_1211_nl);
  mux_1220_nl <= MUX_s_1_2_2(mux_1219_nl, nor_536_nl, fsm_output(2));
  vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1220_nl AND (fsm_output(1));
  nor_520_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_sva(1)) OR (NOT((COMP_LOOP_acc_10_cse_10_1_sva(2))
      AND (COMP_LOOP_acc_10_cse_10_1_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_sva(4))
      AND (COMP_LOOP_acc_10_cse_10_1_sva(0)) AND (fsm_output(7)))));
  nor_521_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (fsm_output(7)));
  mux_1232_nl <= MUX_s_1_2_2(nor_520_nl, nor_521_nl, fsm_output(4));
  nor_522_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1110"))))
      OR nand_446_cse);
  nor_523_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (fsm_output(7)));
  mux_1231_nl <= MUX_s_1_2_2(nor_522_nl, nor_523_nl, fsm_output(4));
  mux_1233_nl <= MUX_s_1_2_2(mux_1232_nl, mux_1231_nl, fsm_output(0));
  and_351_nl <= (fsm_output(6)) AND mux_1233_nl;
  or_1751_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_266_cse;
  or_1749_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (fsm_output(7));
  mux_1229_nl <= MUX_s_1_2_2(or_1751_nl, or_1749_nl, fsm_output(4));
  or_1748_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"))
      OR nand_297_cse;
  or_1746_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (fsm_output(7));
  mux_1228_nl <= MUX_s_1_2_2(or_1748_nl, or_1746_nl, fsm_output(4));
  mux_1230_nl <= MUX_s_1_2_2(mux_1229_nl, mux_1228_nl, fsm_output(0));
  nor_524_nl <= NOT((fsm_output(6)) OR mux_1230_nl);
  mux_1234_nl <= MUX_s_1_2_2(and_351_nl, nor_524_nl, fsm_output(3));
  nand_477_nl <= NOT((fsm_output(5)) AND mux_1234_nl);
  nor_526_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1110"))))
      OR nand_448_cse);
  nor_527_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (fsm_output(7)));
  mux_1225_nl <= MUX_s_1_2_2(nor_526_nl, nor_527_nl, fsm_output(4));
  and_524_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(7));
  nor_529_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(7)));
  mux_1224_nl <= MUX_s_1_2_2(and_524_nl, nor_529_nl, fsm_output(4));
  and_352_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1224_nl;
  mux_1226_nl <= MUX_s_1_2_2(mux_1225_nl, and_352_nl, fsm_output(0));
  nand_168_nl <= NOT((fsm_output(6)) AND mux_1226_nl);
  nand_512_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND (fsm_output(7)));
  or_1735_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (fsm_output(7));
  mux_1222_nl <= MUX_s_1_2_2(nand_512_nl, or_1735_nl, fsm_output(4));
  nand_166_nl <= NOT(nor_98_cse AND mux_1221_cse);
  mux_1223_nl <= MUX_s_1_2_2(mux_1222_nl, nand_166_nl, fsm_output(0));
  or_1738_nl <= (fsm_output(6)) OR mux_1223_nl;
  mux_1227_nl <= MUX_s_1_2_2(nand_168_nl, or_1738_nl, fsm_output(3));
  or_2251_nl <= (fsm_output(5)) OR mux_1227_nl;
  mux_1235_nl <= MUX_s_1_2_2(nand_477_nl, or_2251_nl, fsm_output(2));
  vec_rsc_0_29_i_we_d_pff <= NOT(mux_1235_nl OR (fsm_output(1)));
  nor_515_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_516_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1249_nl <= MUX_s_1_2_2(nor_515_nl, nor_516_nl, fsm_output(0));
  and_348_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_1216_cse);
  and_349_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND (fsm_output(4)) AND (fsm_output(6)) AND (NOT (fsm_output(7)));
  and_523_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  nor_518_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1243_nl <= MUX_s_1_2_2(and_523_nl, nor_518_nl, fsm_output(4));
  mux_1244_nl <= MUX_s_1_2_2(and_349_nl, mux_1243_nl, fsm_output(3));
  mux_1248_nl <= MUX_s_1_2_2(and_348_nl, mux_1244_nl, fsm_output(0));
  mux_1250_nl <= MUX_s_1_2_2(mux_1249_nl, mux_1248_nl, fsm_output(5));
  or_1768_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)) OR nand_443_cse;
  nand_251_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("01")));
  mux_1240_nl <= MUX_s_1_2_2(or_1768_nl, nand_251_nl, fsm_output(4));
  nand_511_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1763_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1239_nl <= MUX_s_1_2_2(nand_511_nl, or_1763_nl, fsm_output(4));
  mux_1241_nl <= MUX_s_1_2_2(mux_1240_nl, mux_1239_nl, fsm_output(3));
  or_1762_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(1)) OR (NOT((COMP_LOOP_acc_10_cse_10_1_sva(2))
      AND (COMP_LOOP_acc_10_cse_10_1_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_sva(4))
      AND (COMP_LOOP_acc_10_cse_10_1_sva(0)) AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("11"))));
  nand_254_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_1237_nl <= MUX_s_1_2_2(or_1762_nl, nand_254_nl, fsm_output(4));
  nand_462_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  or_1758_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1236_nl <= MUX_s_1_2_2(nand_462_nl, or_1758_nl, fsm_output(4));
  mux_1238_nl <= MUX_s_1_2_2(mux_1237_nl, mux_1236_nl, fsm_output(3));
  mux_1242_nl <= MUX_s_1_2_2(mux_1241_nl, mux_1238_nl, fsm_output(0));
  nor_519_nl <= NOT((fsm_output(5)) OR mux_1242_nl);
  mux_1251_nl <= MUX_s_1_2_2(mux_1250_nl, nor_519_nl, fsm_output(2));
  vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1251_nl AND (fsm_output(1));
  and_529_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (fsm_output(7));
  nor_507_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(7)));
  mux_1263_nl <= MUX_s_1_2_2(and_529_nl, nor_507_nl, fsm_output(4));
  and_530_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (fsm_output(7));
  nor_509_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(7)));
  mux_1262_nl <= MUX_s_1_2_2(and_530_nl, nor_509_nl, fsm_output(4));
  mux_1264_nl <= MUX_s_1_2_2(mux_1263_nl, mux_1262_nl, fsm_output(0));
  and_347_nl <= (fsm_output(6)) AND mux_1264_nl;
  or_1796_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(0)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4
      DOWNTO 1)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(7))));
  or_1795_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(7));
  mux_1260_nl <= MUX_s_1_2_2(or_1796_nl, or_1795_nl, fsm_output(4));
  nand_510_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (fsm_output(7)));
  or_1792_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(7));
  mux_1259_nl <= MUX_s_1_2_2(nand_510_nl, or_1792_nl, fsm_output(4));
  mux_1261_nl <= MUX_s_1_2_2(mux_1260_nl, mux_1259_nl, fsm_output(0));
  nor_510_nl <= NOT((fsm_output(6)) OR mux_1261_nl);
  mux_1265_nl <= MUX_s_1_2_2(and_347_nl, nor_510_nl, fsm_output(3));
  nand_476_nl <= NOT((fsm_output(5)) AND mux_1265_nl);
  and_531_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (fsm_output(7));
  nor_513_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(7)));
  mux_1256_nl <= MUX_s_1_2_2(and_531_nl, nor_513_nl, fsm_output(4));
  nand_243_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(7)));
  nand_244_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(7))));
  mux_1255_nl <= MUX_s_1_2_2(nand_243_nl, nand_244_nl, fsm_output(4));
  nor_514_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1255_nl);
  mux_1257_nl <= MUX_s_1_2_2(mux_1256_nl, nor_514_nl, fsm_output(0));
  nand_173_nl <= NOT((fsm_output(6)) AND mux_1257_nl);
  or_1784_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4
      DOWNTO 1)=STD_LOGIC_VECTOR'("1111")) AND (fsm_output(7))));
  or_1783_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(7));
  mux_1253_nl <= MUX_s_1_2_2(or_1784_nl, or_1783_nl, fsm_output(4));
  or_1782_nl <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1190_cse;
  mux_1254_nl <= MUX_s_1_2_2(mux_1253_nl, or_1782_nl, fsm_output(0));
  or_1785_nl <= (fsm_output(6)) OR mux_1254_nl;
  mux_1258_nl <= MUX_s_1_2_2(nand_173_nl, or_1785_nl, fsm_output(3));
  or_2250_nl <= (fsm_output(5)) OR mux_1258_nl;
  mux_1266_nl <= MUX_s_1_2_2(nand_476_nl, or_2250_nl, fsm_output(2));
  vec_rsc_0_30_i_we_d_pff <= NOT(mux_1266_nl OR (fsm_output(1)));
  nor_500_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_501_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1280_nl <= MUX_s_1_2_2(nor_500_nl, nor_501_nl, fsm_output(0));
  nor_502_nl <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) OR mux_1278_cse);
  and_345_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (fsm_output(4)) AND (fsm_output(6)) AND (NOT (fsm_output(7)));
  and_522_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  nor_504_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1274_nl <= MUX_s_1_2_2(and_522_nl, nor_504_nl, fsm_output(4));
  mux_1275_nl <= MUX_s_1_2_2(and_345_nl, mux_1274_nl, fsm_output(3));
  mux_1279_nl <= MUX_s_1_2_2(nor_502_nl, mux_1275_nl, fsm_output(0));
  mux_1281_nl <= MUX_s_1_2_2(mux_1280_nl, mux_1279_nl, fsm_output(5));
  or_1815_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)) OR nand_443_cse;
  nand_231_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("01")));
  mux_1271_nl <= MUX_s_1_2_2(or_1815_nl, nand_231_nl, fsm_output(4));
  nand_509_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  or_1810_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("00"));
  mux_1270_nl <= MUX_s_1_2_2(nand_509_nl, or_1810_nl, fsm_output(4));
  mux_1272_nl <= MUX_s_1_2_2(mux_1271_nl, mux_1270_nl, fsm_output(3));
  or_1809_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))))
      OR nand_443_cse;
  nand_234_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_1268_nl <= MUX_s_1_2_2(or_1809_nl, nand_234_nl, fsm_output(4));
  nand_460_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  or_1804_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_1267_nl <= MUX_s_1_2_2(nand_460_nl, or_1804_nl, fsm_output(4));
  mux_1269_nl <= MUX_s_1_2_2(mux_1268_nl, mux_1267_nl, fsm_output(3));
  mux_1273_nl <= MUX_s_1_2_2(mux_1272_nl, mux_1269_nl, fsm_output(0));
  nor_505_nl <= NOT((fsm_output(5)) OR mux_1273_nl);
  mux_1282_nl <= MUX_s_1_2_2(mux_1281_nl, nor_505_nl, fsm_output(2));
  vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1282_nl AND (fsm_output(1));
  and_334_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(7));
  and_335_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (NOT (fsm_output(7)));
  mux_1294_nl <= MUX_s_1_2_2(and_334_nl, and_335_nl, fsm_output(4));
  and_336_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(7));
  and_337_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (NOT (fsm_output(7)));
  mux_1293_nl <= MUX_s_1_2_2(and_336_nl, and_337_nl, fsm_output(4));
  mux_1295_nl <= MUX_s_1_2_2(mux_1294_nl, mux_1293_nl, fsm_output(0));
  and_333_nl <= (fsm_output(6)) AND mux_1295_nl;
  nand_223_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(7)));
  nand_224_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (NOT (fsm_output(7))));
  mux_1291_nl <= MUX_s_1_2_2(nand_223_nl, nand_224_nl, fsm_output(4));
  nand_225_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(7)));
  nand_226_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (NOT (fsm_output(7))));
  mux_1290_nl <= MUX_s_1_2_2(nand_225_nl, nand_226_nl, fsm_output(4));
  mux_1292_nl <= MUX_s_1_2_2(mux_1291_nl, mux_1290_nl, fsm_output(0));
  nor_498_nl <= NOT((fsm_output(6)) OR mux_1292_nl);
  mux_1296_nl <= MUX_s_1_2_2(and_333_nl, nor_498_nl, fsm_output(3));
  nand_475_nl <= NOT((fsm_output(5)) AND mux_1296_nl);
  and_338_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(7));
  and_339_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (NOT (fsm_output(7)));
  mux_1287_nl <= MUX_s_1_2_2(and_338_nl, and_339_nl, fsm_output(4));
  and_341_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(7));
  and_342_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(7)));
  mux_1286_nl <= MUX_s_1_2_2(and_341_nl, and_342_nl, fsm_output(4));
  and_340_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND mux_1286_nl;
  mux_1288_nl <= MUX_s_1_2_2(mux_1287_nl, and_340_nl, fsm_output(0));
  nand_179_nl <= NOT((fsm_output(6)) AND mux_1288_nl);
  nand_227_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(7)));
  nand_228_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (NOT (fsm_output(7))));
  mux_1284_nl <= MUX_s_1_2_2(nand_227_nl, nand_228_nl, fsm_output(4));
  nand_177_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND mux_1221_cse);
  mux_1285_nl <= MUX_s_1_2_2(mux_1284_nl, nand_177_nl, fsm_output(0));
  or_1830_nl <= (fsm_output(6)) OR mux_1285_nl;
  mux_1289_nl <= MUX_s_1_2_2(nand_179_nl, or_1830_nl, fsm_output(3));
  or_2249_nl <= (fsm_output(5)) OR mux_1289_nl;
  mux_1297_nl <= MUX_s_1_2_2(nand_475_nl, or_2249_nl, fsm_output(2));
  vec_rsc_0_31_i_we_d_pff <= NOT(mux_1297_nl OR (fsm_output(1)));
  nor_494_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11111"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  nor_495_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_1311_nl <= MUX_s_1_2_2(nor_494_nl, nor_495_nl, fsm_output(0));
  and_329_nl <= (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT mux_1278_cse);
  and_330_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(4)) AND (fsm_output(6)) AND (NOT (fsm_output(7)));
  and_521_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  and_331_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("00"));
  mux_1305_nl <= MUX_s_1_2_2(and_521_nl, and_331_nl, fsm_output(4));
  mux_1306_nl <= MUX_s_1_2_2(and_330_nl, mux_1305_nl, fsm_output(3));
  mux_1310_nl <= MUX_s_1_2_2(and_329_nl, mux_1306_nl, fsm_output(0));
  mux_1312_nl <= MUX_s_1_2_2(mux_1311_nl, mux_1310_nl, fsm_output(5));
  or_1848_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm)) OR nand_443_cse;
  nand_214_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("01")));
  mux_1302_nl <= MUX_s_1_2_2(or_1848_nl, nand_214_nl, fsm_output(4));
  nand_508_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("10")));
  nand_216_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(fsm_output(7 DOWNTO
      6)=STD_LOGIC_VECTOR'("00")));
  mux_1301_nl <= MUX_s_1_2_2(nand_508_nl, nand_216_nl, fsm_output(4));
  mux_1303_nl <= MUX_s_1_2_2(mux_1302_nl, mux_1301_nl, fsm_output(3));
  nand_217_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")));
  nand_218_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  mux_1299_nl <= MUX_s_1_2_2(nand_217_nl, nand_218_nl, fsm_output(4));
  nand_458_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  nand_220_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("00")));
  mux_1298_nl <= MUX_s_1_2_2(nand_458_nl, nand_220_nl, fsm_output(4));
  mux_1300_nl <= MUX_s_1_2_2(mux_1299_nl, mux_1298_nl, fsm_output(3));
  mux_1304_nl <= MUX_s_1_2_2(mux_1303_nl, mux_1300_nl, fsm_output(0));
  nor_497_nl <= NOT((fsm_output(5)) OR mux_1304_nl);
  mux_1313_nl <= MUX_s_1_2_2(mux_1312_nl, nor_497_nl, fsm_output(2));
  vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1313_nl AND (fsm_output(1));
  twiddle_rsc_0_0_i_radr_d_pff <= MUX1HOT_v_5_7_2((z_out_8(6 DOWNTO 2)), (z_out_7(9
      DOWNTO 5)), (z_out_7(8 DOWNTO 4)), (COMP_LOOP_5_tmp_mul_idiv_sva(7 DOWNTO 3)),
      (COMP_LOOP_2_tmp_mul_idiv_sva(9 DOWNTO 5)), (COMP_LOOP_3_tmp_lshift_ncse_sva(8
      DOWNTO 4)), (COMP_LOOP_2_tmp_lshift_ncse_sva(9 DOWNTO 5)), STD_LOGIC_VECTOR'(
      and_dcpl_46 & COMP_LOOP_or_42_cse & and_dcpl_171 & and_dcpl_173 & and_dcpl_174
      & and_dcpl_176 & and_dcpl_177));
  nor_489_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(3)));
  nor_486_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(3))));
  nor_487_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(3))));
  mux_1318_nl <= MUX_s_1_2_2(nor_486_nl, nor_487_nl, fsm_output(0));
  nor_488_nl <= NOT(CONV_SL_1_1(z_out_8(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (fsm_output(3)));
  mux_1317_nl <= MUX_s_1_2_2(nor_488_nl, nor_489_cse, fsm_output(0));
  mux_1319_nl <= MUX_s_1_2_2(mux_1318_nl, mux_1317_nl, fsm_output(1));
  nor_490_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      (fsm_output(3)));
  mux_1315_nl <= MUX_s_1_2_2(nor_490_nl, nor_489_cse, fsm_output(0));
  nor_492_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)));
  nor_493_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(3)));
  mux_1314_nl <= MUX_s_1_2_2(nor_492_nl, nor_493_nl, fsm_output(0));
  mux_1316_nl <= MUX_s_1_2_2(mux_1315_nl, mux_1314_nl, fsm_output(1));
  mux_1320_nl <= MUX_s_1_2_2(mux_1319_nl, mux_1316_nl, fsm_output(2));
  twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1320_nl AND and_dcpl_179;
  twiddle_rsc_0_1_i_radr_d_pff <= z_out_7(9 DOWNTO 5);
  nor_483_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT and_316_cse));
  nor_484_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1322_nl <= MUX_s_1_2_2(nor_483_nl, nor_484_nl, fsm_output(3));
  or_1872_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001")) OR (NOT
      (fsm_output(1)));
  or_1870_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001")) OR (fsm_output(1));
  mux_1321_nl <= MUX_s_1_2_2(or_1872_nl, or_1870_nl, fsm_output(0));
  nor_485_nl <= NOT((fsm_output(3)) OR mux_1321_nl);
  mux_1323_nl <= MUX_s_1_2_2(mux_1322_nl, nor_485_nl, fsm_output(2));
  twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1323_nl AND and_dcpl_179;
  twiddle_rsc_0_2_i_radr_d_pff <= MUX_v_5_2_2((z_out_7(9 DOWNTO 5)), (z_out_7(8 DOWNTO
      4)), COMP_LOOP_tmp_or_35_cse);
  nor_480_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(3)));
  nor_479_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(3)));
  nor_477_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(3))));
  nor_478_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(3)));
  mux_1327_nl <= MUX_s_1_2_2(nor_477_nl, nor_478_nl, fsm_output(1));
  mux_1325_nl <= MUX_s_1_2_2(nor_479_cse, nor_480_cse, fsm_output(0));
  mux_1324_nl <= MUX_s_1_2_2(nor_480_cse, nor_479_cse, fsm_output(0));
  mux_1326_nl <= MUX_s_1_2_2(mux_1325_nl, mux_1324_nl, fsm_output(1));
  mux_1328_nl <= MUX_s_1_2_2(mux_1327_nl, mux_1326_nl, fsm_output(2));
  twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1328_nl AND and_dcpl_179;
  nor_474_nl <= NOT((z_out_7(3)) OR (z_out_7(4)) OR (NOT (z_out_7(0))) OR (z_out_7(2))
      OR not_tmp_618);
  nor_475_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1330_nl <= MUX_s_1_2_2(nor_474_nl, nor_475_nl, fsm_output(3));
  or_1886_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000")) OR not_tmp_617;
  or_1884_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011")) OR (fsm_output(1));
  mux_1329_nl <= MUX_s_1_2_2(or_1886_nl, or_1884_nl, fsm_output(0));
  nor_476_nl <= NOT((fsm_output(3)) OR mux_1329_nl);
  mux_1331_nl <= MUX_s_1_2_2(mux_1330_nl, nor_476_nl, fsm_output(2));
  twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1331_nl AND and_dcpl_179;
  twiddle_rsc_0_4_i_radr_d_pff <= MUX1HOT_v_5_6_2((z_out_7(9 DOWNTO 5)), (z_out_7(8
      DOWNTO 4)), (COMP_LOOP_5_tmp_mul_idiv_sva(7 DOWNTO 3)), (COMP_LOOP_2_tmp_mul_idiv_sva(9
      DOWNTO 5)), (COMP_LOOP_3_tmp_lshift_ncse_sva(8 DOWNTO 4)), (COMP_LOOP_2_tmp_lshift_ncse_sva(9
      DOWNTO 5)), STD_LOGIC_VECTOR'( COMP_LOOP_or_42_cse & and_dcpl_171 & and_dcpl_173
      & and_dcpl_174 & and_dcpl_176 & and_dcpl_177));
  nor_467_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(3))));
  nor_468_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(3))));
  mux_1335_nl <= MUX_s_1_2_2(nor_467_nl, nor_468_nl, fsm_output(0));
  nor_469_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(3)));
  mux_1336_nl <= MUX_s_1_2_2(mux_1335_nl, nor_469_nl, fsm_output(1));
  nor_470_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR
      (fsm_output(3)));
  nor_471_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(3)));
  mux_1333_nl <= MUX_s_1_2_2(nor_470_nl, nor_471_nl, fsm_output(0));
  nor_472_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)));
  nor_473_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(3)));
  mux_1332_nl <= MUX_s_1_2_2(nor_472_nl, nor_473_nl, fsm_output(0));
  mux_1334_nl <= MUX_s_1_2_2(mux_1333_nl, mux_1332_nl, fsm_output(1));
  mux_1337_nl <= MUX_s_1_2_2(mux_1336_nl, mux_1334_nl, fsm_output(2));
  twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1337_nl AND and_dcpl_179;
  nor_464_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT and_316_cse));
  nor_465_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1339_nl <= MUX_s_1_2_2(nor_464_nl, nor_465_nl, fsm_output(3));
  or_1902_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101")) OR (NOT
      (fsm_output(1)));
  or_1900_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101")) OR (fsm_output(1));
  mux_1338_nl <= MUX_s_1_2_2(or_1902_nl, or_1900_nl, fsm_output(0));
  nor_466_nl <= NOT((fsm_output(3)) OR mux_1338_nl);
  mux_1340_nl <= MUX_s_1_2_2(mux_1339_nl, nor_466_nl, fsm_output(2));
  twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1340_nl AND and_dcpl_179;
  nor_461_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(3)));
  nor_460_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(3)));
  nor_458_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(3))));
  nor_459_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(3)));
  mux_1344_nl <= MUX_s_1_2_2(nor_458_nl, nor_459_nl, fsm_output(1));
  mux_1342_nl <= MUX_s_1_2_2(nor_460_cse, nor_461_cse, fsm_output(0));
  mux_1341_nl <= MUX_s_1_2_2(nor_461_cse, nor_460_cse, fsm_output(0));
  mux_1343_nl <= MUX_s_1_2_2(mux_1342_nl, mux_1341_nl, fsm_output(1));
  mux_1345_nl <= MUX_s_1_2_2(mux_1344_nl, mux_1343_nl, fsm_output(2));
  twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1345_nl AND and_dcpl_179;
  nor_455_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00")) OR
      not_tmp_625);
  nor_456_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1347_nl <= MUX_s_1_2_2(nor_455_nl, nor_456_nl, fsm_output(3));
  or_1916_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("001")) OR not_tmp_617;
  or_1914_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111")) OR (fsm_output(1));
  mux_1346_nl <= MUX_s_1_2_2(or_1916_nl, or_1914_nl, fsm_output(0));
  nor_457_nl <= NOT((fsm_output(3)) OR mux_1346_nl);
  mux_1348_nl <= MUX_s_1_2_2(mux_1347_nl, nor_457_nl, fsm_output(2));
  twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1348_nl AND and_dcpl_179;
  nor_450_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(3)));
  nor_447_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(3))));
  nor_448_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(3))));
  mux_1353_nl <= MUX_s_1_2_2(nor_447_nl, nor_448_nl, fsm_output(0));
  nor_449_nl <= NOT(CONV_SL_1_1(z_out_8(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(3)));
  mux_1352_nl <= MUX_s_1_2_2(nor_449_nl, nor_450_cse, fsm_output(0));
  mux_1354_nl <= MUX_s_1_2_2(mux_1353_nl, mux_1352_nl, fsm_output(1));
  nor_451_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR
      (fsm_output(3)));
  mux_1350_nl <= MUX_s_1_2_2(nor_451_nl, nor_450_cse, fsm_output(0));
  nor_453_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)));
  nor_454_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(3)));
  mux_1349_nl <= MUX_s_1_2_2(nor_453_nl, nor_454_nl, fsm_output(0));
  mux_1351_nl <= MUX_s_1_2_2(mux_1350_nl, mux_1349_nl, fsm_output(1));
  mux_1355_nl <= MUX_s_1_2_2(mux_1354_nl, mux_1351_nl, fsm_output(2));
  twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1355_nl AND and_dcpl_179;
  nor_444_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT and_316_cse));
  nor_445_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1357_nl <= MUX_s_1_2_2(nor_444_nl, nor_445_nl, fsm_output(3));
  or_1933_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001")) OR (NOT
      (fsm_output(1)));
  or_1931_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001")) OR (fsm_output(1));
  mux_1356_nl <= MUX_s_1_2_2(or_1933_nl, or_1931_nl, fsm_output(0));
  nor_446_nl <= NOT((fsm_output(3)) OR mux_1356_nl);
  mux_1358_nl <= MUX_s_1_2_2(mux_1357_nl, nor_446_nl, fsm_output(2));
  twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1358_nl AND and_dcpl_179;
  nor_441_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(3)));
  nor_440_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(3)));
  nor_438_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(3))));
  nor_439_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(3)));
  mux_1362_nl <= MUX_s_1_2_2(nor_438_nl, nor_439_nl, fsm_output(1));
  mux_1360_nl <= MUX_s_1_2_2(nor_440_cse, nor_441_cse, fsm_output(0));
  mux_1359_nl <= MUX_s_1_2_2(nor_441_cse, nor_440_cse, fsm_output(0));
  mux_1361_nl <= MUX_s_1_2_2(mux_1360_nl, mux_1359_nl, fsm_output(1));
  mux_1363_nl <= MUX_s_1_2_2(mux_1362_nl, mux_1361_nl, fsm_output(2));
  twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1363_nl AND and_dcpl_179;
  nor_435_nl <= NOT((NOT (z_out_7(3))) OR (z_out_7(4)) OR (NOT (z_out_7(0))) OR (z_out_7(2))
      OR not_tmp_618);
  nor_436_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1365_nl <= MUX_s_1_2_2(nor_435_nl, nor_436_nl, fsm_output(3));
  or_1947_nl <= (z_out_7(2)) OR (z_out_7(4)) OR not_tmp_632;
  or_1945_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011")) OR (fsm_output(1));
  mux_1364_nl <= MUX_s_1_2_2(or_1947_nl, or_1945_nl, fsm_output(0));
  nor_437_nl <= NOT((fsm_output(3)) OR mux_1364_nl);
  mux_1366_nl <= MUX_s_1_2_2(mux_1365_nl, nor_437_nl, fsm_output(2));
  twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1366_nl AND and_dcpl_179;
  nor_428_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(3))));
  nor_429_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(3))));
  mux_1370_nl <= MUX_s_1_2_2(nor_428_nl, nor_429_nl, fsm_output(0));
  nor_430_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(3)));
  mux_1371_nl <= MUX_s_1_2_2(mux_1370_nl, nor_430_nl, fsm_output(1));
  nor_431_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR
      (fsm_output(3)));
  nor_432_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(3)));
  mux_1368_nl <= MUX_s_1_2_2(nor_431_nl, nor_432_nl, fsm_output(0));
  nor_433_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)));
  nor_434_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(3)));
  mux_1367_nl <= MUX_s_1_2_2(nor_433_nl, nor_434_nl, fsm_output(0));
  mux_1369_nl <= MUX_s_1_2_2(mux_1368_nl, mux_1367_nl, fsm_output(1));
  mux_1372_nl <= MUX_s_1_2_2(mux_1371_nl, mux_1369_nl, fsm_output(2));
  twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1372_nl AND and_dcpl_179;
  nor_425_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT and_316_cse));
  nor_426_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1374_nl <= MUX_s_1_2_2(nor_425_nl, nor_426_nl, fsm_output(3));
  or_1963_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101")) OR (NOT
      (fsm_output(1)));
  or_1961_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101")) OR (fsm_output(1));
  mux_1373_nl <= MUX_s_1_2_2(or_1963_nl, or_1961_nl, fsm_output(0));
  nor_427_nl <= NOT((fsm_output(3)) OR mux_1373_nl);
  mux_1375_nl <= MUX_s_1_2_2(mux_1374_nl, nor_427_nl, fsm_output(2));
  twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1375_nl AND and_dcpl_179;
  nor_422_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(3)));
  nor_421_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(3)));
  nor_419_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(3))));
  nor_420_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(3)));
  mux_1379_nl <= MUX_s_1_2_2(nor_419_nl, nor_420_nl, fsm_output(1));
  mux_1377_nl <= MUX_s_1_2_2(nor_421_cse, nor_422_cse, fsm_output(0));
  mux_1376_nl <= MUX_s_1_2_2(nor_422_cse, nor_421_cse, fsm_output(0));
  mux_1378_nl <= MUX_s_1_2_2(mux_1377_nl, mux_1376_nl, fsm_output(1));
  mux_1380_nl <= MUX_s_1_2_2(mux_1379_nl, mux_1378_nl, fsm_output(2));
  twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1380_nl AND and_dcpl_179;
  nor_416_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("01")) OR
      not_tmp_625);
  nor_417_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1382_nl <= MUX_s_1_2_2(nor_416_nl, nor_417_nl, fsm_output(3));
  or_1977_nl <= (NOT (z_out_7(2))) OR (z_out_7(4)) OR not_tmp_632;
  or_1975_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111")) OR (fsm_output(1));
  mux_1381_nl <= MUX_s_1_2_2(or_1977_nl, or_1975_nl, fsm_output(0));
  nor_418_nl <= NOT((fsm_output(3)) OR mux_1381_nl);
  mux_1383_nl <= MUX_s_1_2_2(mux_1382_nl, nor_418_nl, fsm_output(2));
  twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1383_nl AND and_dcpl_179;
  nor_411_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(3)));
  nor_408_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_204_cse);
  nor_409_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_205_cse);
  mux_1388_nl <= MUX_s_1_2_2(nor_408_nl, nor_409_nl, fsm_output(0));
  nor_410_nl <= NOT(CONV_SL_1_1(z_out_8(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (fsm_output(3)));
  mux_1387_nl <= MUX_s_1_2_2(nor_410_nl, nor_411_cse, fsm_output(0));
  mux_1389_nl <= MUX_s_1_2_2(mux_1388_nl, mux_1387_nl, fsm_output(1));
  nor_412_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR
      (fsm_output(3)));
  mux_1385_nl <= MUX_s_1_2_2(nor_412_nl, nor_411_cse, fsm_output(0));
  nor_414_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)));
  nor_415_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(3)));
  mux_1384_nl <= MUX_s_1_2_2(nor_414_nl, nor_415_nl, fsm_output(0));
  mux_1386_nl <= MUX_s_1_2_2(mux_1385_nl, mux_1384_nl, fsm_output(1));
  mux_1390_nl <= MUX_s_1_2_2(mux_1389_nl, mux_1386_nl, fsm_output(2));
  twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1390_nl AND and_dcpl_179;
  nor_405_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT and_316_cse));
  nor_406_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1392_nl <= MUX_s_1_2_2(nor_405_nl, nor_406_nl, fsm_output(3));
  or_1994_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001")) OR (NOT
      (fsm_output(1)));
  or_1992_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001")) OR (fsm_output(1));
  mux_1391_nl <= MUX_s_1_2_2(or_1994_nl, or_1992_nl, fsm_output(0));
  nor_407_nl <= NOT((fsm_output(3)) OR mux_1391_nl);
  mux_1393_nl <= MUX_s_1_2_2(mux_1392_nl, nor_407_nl, fsm_output(2));
  twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1393_nl AND and_dcpl_179;
  nor_402_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(3)));
  nor_401_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(3)));
  nor_399_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(3))));
  nor_400_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(3)));
  mux_1397_nl <= MUX_s_1_2_2(nor_399_nl, nor_400_nl, fsm_output(1));
  mux_1395_nl <= MUX_s_1_2_2(nor_401_cse, nor_402_cse, fsm_output(0));
  mux_1394_nl <= MUX_s_1_2_2(nor_402_cse, nor_401_cse, fsm_output(0));
  mux_1396_nl <= MUX_s_1_2_2(mux_1395_nl, mux_1394_nl, fsm_output(1));
  mux_1398_nl <= MUX_s_1_2_2(mux_1397_nl, mux_1396_nl, fsm_output(2));
  twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1398_nl AND and_dcpl_179;
  nor_396_nl <= NOT((z_out_7(3)) OR (NOT (z_out_7(4))) OR (NOT (z_out_7(0))) OR (z_out_7(2))
      OR not_tmp_618);
  nor_397_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1400_nl <= MUX_s_1_2_2(nor_396_nl, nor_397_nl, fsm_output(3));
  or_2008_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("100")) OR not_tmp_617;
  or_2006_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011")) OR (fsm_output(1));
  mux_1399_nl <= MUX_s_1_2_2(or_2008_nl, or_2006_nl, fsm_output(0));
  nor_398_nl <= NOT((fsm_output(3)) OR mux_1399_nl);
  mux_1401_nl <= MUX_s_1_2_2(mux_1400_nl, nor_398_nl, fsm_output(2));
  twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1401_nl AND and_dcpl_179;
  nor_389_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_204_cse);
  nor_390_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_205_cse);
  mux_1405_nl <= MUX_s_1_2_2(nor_389_nl, nor_390_nl, fsm_output(0));
  nor_391_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(3)));
  mux_1406_nl <= MUX_s_1_2_2(mux_1405_nl, nor_391_nl, fsm_output(1));
  nor_392_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR
      (fsm_output(3)));
  nor_393_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(3)));
  mux_1403_nl <= MUX_s_1_2_2(nor_392_nl, nor_393_nl, fsm_output(0));
  nor_394_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)));
  nor_395_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(3)));
  mux_1402_nl <= MUX_s_1_2_2(nor_394_nl, nor_395_nl, fsm_output(0));
  mux_1404_nl <= MUX_s_1_2_2(mux_1403_nl, mux_1402_nl, fsm_output(1));
  mux_1407_nl <= MUX_s_1_2_2(mux_1406_nl, mux_1404_nl, fsm_output(2));
  twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1407_nl AND and_dcpl_179;
  nor_386_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT and_316_cse));
  nor_387_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1409_nl <= MUX_s_1_2_2(nor_386_nl, nor_387_nl, fsm_output(3));
  or_2024_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101")) OR (NOT
      (fsm_output(1)));
  or_2022_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101")) OR (fsm_output(1));
  mux_1408_nl <= MUX_s_1_2_2(or_2024_nl, or_2022_nl, fsm_output(0));
  nor_388_nl <= NOT((fsm_output(3)) OR mux_1408_nl);
  mux_1410_nl <= MUX_s_1_2_2(mux_1409_nl, nor_388_nl, fsm_output(2));
  twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1410_nl AND and_dcpl_179;
  nor_383_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(3)));
  nor_382_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(3)));
  nor_380_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(3))));
  nor_381_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(3)));
  mux_1414_nl <= MUX_s_1_2_2(nor_380_nl, nor_381_nl, fsm_output(1));
  mux_1412_nl <= MUX_s_1_2_2(nor_382_cse, nor_383_cse, fsm_output(0));
  mux_1411_nl <= MUX_s_1_2_2(nor_383_cse, nor_382_cse, fsm_output(0));
  mux_1413_nl <= MUX_s_1_2_2(mux_1412_nl, mux_1411_nl, fsm_output(1));
  mux_1415_nl <= MUX_s_1_2_2(mux_1414_nl, mux_1413_nl, fsm_output(2));
  twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1415_nl AND and_dcpl_179;
  nor_377_nl <= NOT((z_out_7(3)) OR (NOT((z_out_7(4)) AND (z_out_7(0)) AND (z_out_7(2))
      AND (z_out_7(1)) AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")))));
  nor_378_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1417_nl <= MUX_s_1_2_2(nor_377_nl, nor_378_nl, fsm_output(3));
  or_2038_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("101")) OR not_tmp_617;
  or_2036_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111")) OR (fsm_output(1));
  mux_1416_nl <= MUX_s_1_2_2(or_2038_nl, or_2036_nl, fsm_output(0));
  nor_379_nl <= NOT((fsm_output(3)) OR mux_1416_nl);
  mux_1418_nl <= MUX_s_1_2_2(mux_1417_nl, nor_379_nl, fsm_output(2));
  twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1418_nl AND and_dcpl_179;
  nor_372_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(3)));
  nor_369_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)))));
  nor_370_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)))));
  mux_1423_nl <= MUX_s_1_2_2(nor_369_nl, nor_370_nl, fsm_output(0));
  nor_371_nl <= NOT(CONV_SL_1_1(z_out_8(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (fsm_output(3)));
  mux_1422_nl <= MUX_s_1_2_2(nor_371_nl, nor_372_cse, fsm_output(0));
  mux_1424_nl <= MUX_s_1_2_2(mux_1423_nl, mux_1422_nl, fsm_output(1));
  nor_373_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR
      (fsm_output(3)));
  mux_1420_nl <= MUX_s_1_2_2(nor_373_nl, nor_372_cse, fsm_output(0));
  nor_375_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)));
  nor_376_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(3)));
  mux_1419_nl <= MUX_s_1_2_2(nor_375_nl, nor_376_nl, fsm_output(0));
  mux_1421_nl <= MUX_s_1_2_2(mux_1420_nl, mux_1419_nl, fsm_output(1));
  mux_1425_nl <= MUX_s_1_2_2(mux_1424_nl, mux_1421_nl, fsm_output(2));
  twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1425_nl AND and_dcpl_179;
  nor_366_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT and_316_cse));
  nor_367_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1427_nl <= MUX_s_1_2_2(nor_366_nl, nor_367_nl, fsm_output(3));
  or_2054_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001")) OR (NOT
      (fsm_output(1)));
  or_2052_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001")) OR (fsm_output(1));
  mux_1426_nl <= MUX_s_1_2_2(or_2054_nl, or_2052_nl, fsm_output(0));
  nor_368_nl <= NOT((fsm_output(3)) OR mux_1426_nl);
  mux_1428_nl <= MUX_s_1_2_2(mux_1427_nl, nor_368_nl, fsm_output(2));
  twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1428_nl AND and_dcpl_179;
  nor_363_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(3)));
  nor_362_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(3)));
  nor_360_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(3))));
  nor_361_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(3)));
  mux_1432_nl <= MUX_s_1_2_2(nor_360_nl, nor_361_nl, fsm_output(1));
  mux_1430_nl <= MUX_s_1_2_2(nor_362_cse, nor_363_cse, fsm_output(0));
  mux_1429_nl <= MUX_s_1_2_2(nor_363_cse, nor_362_cse, fsm_output(0));
  mux_1431_nl <= MUX_s_1_2_2(mux_1430_nl, mux_1429_nl, fsm_output(1));
  mux_1433_nl <= MUX_s_1_2_2(mux_1432_nl, mux_1431_nl, fsm_output(2));
  twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1433_nl AND and_dcpl_179;
  nor_357_nl <= NOT((NOT((z_out_7(3)) AND (z_out_7(4)) AND (z_out_7(0)) AND (NOT
      (z_out_7(2))))) OR not_tmp_618);
  nor_358_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1435_nl <= MUX_s_1_2_2(nor_357_nl, nor_358_nl, fsm_output(3));
  or_2067_nl <= (z_out_7(2)) OR (NOT((z_out_7(4)) AND (z_out_7(3)) AND (z_out_7(0))
      AND (z_out_7(1)) AND (fsm_output(1))));
  or_2066_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011")) OR (fsm_output(1));
  mux_1434_nl <= MUX_s_1_2_2(or_2067_nl, or_2066_nl, fsm_output(0));
  nor_359_nl <= NOT((fsm_output(3)) OR mux_1434_nl);
  mux_1436_nl <= MUX_s_1_2_2(mux_1435_nl, nor_359_nl, fsm_output(2));
  twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1436_nl AND and_dcpl_179;
  nor_351_nl <= NOT((COMP_LOOP_3_tmp_lshift_ncse_sva(0)) OR (NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(3
      DOWNTO 1)=STD_LOGIC_VECTOR'("111")) AND (fsm_output(3)))));
  nor_352_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)))));
  mux_1440_nl <= MUX_s_1_2_2(nor_351_nl, nor_352_nl, fsm_output(0));
  nor_353_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(3)));
  mux_1441_nl <= MUX_s_1_2_2(mux_1440_nl, nor_353_nl, fsm_output(1));
  nor_354_nl <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR
      (fsm_output(3)));
  nor_355_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(3)));
  mux_1438_nl <= MUX_s_1_2_2(nor_354_nl, nor_355_nl, fsm_output(0));
  and_328_nl <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (fsm_output(3)));
  nor_356_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(3)));
  mux_1437_nl <= MUX_s_1_2_2(and_328_nl, nor_356_nl, fsm_output(0));
  mux_1439_nl <= MUX_s_1_2_2(mux_1438_nl, mux_1437_nl, fsm_output(1));
  mux_1442_nl <= MUX_s_1_2_2(mux_1441_nl, mux_1439_nl, fsm_output(2));
  twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1442_nl AND and_dcpl_179;
  and_327_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101")) AND and_316_cse;
  nor_349_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  mux_1444_nl <= MUX_s_1_2_2(and_327_nl, nor_349_nl, fsm_output(3));
  nand_474_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND (fsm_output(1)));
  or_2080_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101")) OR (fsm_output(1));
  mux_1443_nl <= MUX_s_1_2_2(nand_474_nl, or_2080_nl, fsm_output(0));
  nor_350_nl <= NOT((fsm_output(3)) OR mux_1443_nl);
  mux_1445_nl <= MUX_s_1_2_2(mux_1444_nl, nor_350_nl, fsm_output(2));
  twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1445_nl AND and_dcpl_179;
  nor_347_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(3)));
  and_325_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND (NOT
      (fsm_output(3)));
  and_323_nl <= (NOT (fsm_output(0))) AND CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (fsm_output(3));
  and_324_nl <= (fsm_output(0)) AND CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (NOT (fsm_output(3)));
  mux_1449_nl <= MUX_s_1_2_2(and_323_nl, and_324_nl, fsm_output(1));
  mux_1447_nl <= MUX_s_1_2_2(and_325_cse, nor_347_cse, fsm_output(0));
  mux_1446_nl <= MUX_s_1_2_2(nor_347_cse, and_325_cse, fsm_output(0));
  mux_1448_nl <= MUX_s_1_2_2(mux_1447_nl, mux_1446_nl, fsm_output(1));
  mux_1450_nl <= MUX_s_1_2_2(mux_1449_nl, mux_1448_nl, fsm_output(2));
  twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1450_nl AND and_dcpl_179;
  and_321_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111")) AND CONV_SL_1_1(fsm_output(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_322_nl <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111")) AND CONV_SL_1_1(fsm_output(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("00"));
  mux_1452_nl <= MUX_s_1_2_2(and_321_nl, and_322_nl, fsm_output(3));
  nand_192_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(1)));
  nand_193_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (NOT (fsm_output(1))));
  mux_1451_nl <= MUX_s_1_2_2(nand_192_nl, nand_193_nl, fsm_output(0));
  nor_346_nl <= NOT((fsm_output(3)) OR mux_1451_nl);
  mux_1453_nl <= MUX_s_1_2_2(mux_1452_nl, nor_346_nl, fsm_output(2));
  twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_1453_nl AND and_dcpl_179;
  and_dcpl_334 <= (fsm_output(6)) AND (fsm_output(7)) AND (fsm_output(1)) AND (fsm_output(0))
      AND and_dcpl_29 AND (NOT (fsm_output(2))) AND (fsm_output(5));
  and_dcpl_347 <= nor_1025_cse AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND and_dcpl_29 AND and_dcpl_28;
  and_dcpl_353 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("00")) AND
      and_dcpl_31;
  and_605_cse <= and_dcpl_353 AND and_dcpl_29 AND (NOT (fsm_output(2))) AND (fsm_output(5));
  and_609_cse <= and_dcpl_353 AND and_479_cse AND and_dcpl_35;
  and_dcpl_365 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")) AND
      and_dcpl_31;
  and_614_cse <= and_dcpl_365 AND and_479_cse AND and_dcpl_28;
  and_617_cse <= and_dcpl_365 AND and_dcpl_59 AND and_dcpl_35;
  and_dcpl_372 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")) AND
      and_dcpl_31;
  and_621_cse <= and_dcpl_372 AND and_dcpl_59 AND and_dcpl_28;
  and_624_cse <= and_dcpl_372 AND and_dcpl_69 AND and_dcpl_35;
  and_628_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")) AND
      and_dcpl_31 AND and_dcpl_69 AND and_dcpl_28;
  and_dcpl_419 <= nor_1025_cse AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_420 <= and_dcpl_419 AND and_dcpl_30;
  and_dcpl_422 <= nor_1025_cse AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_423 <= and_dcpl_422 AND and_dcpl_30;
  and_dcpl_425 <= and_dcpl_29 AND (fsm_output(2)) AND (NOT (fsm_output(5)));
  and_dcpl_428 <= nor_1025_cse AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))
      AND and_dcpl_425;
  and_dcpl_429 <= and_dcpl_419 AND and_dcpl_425;
  and_dcpl_433 <= nor_1025_cse AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("00"));
  and_dcpl_434 <= and_dcpl_433 AND CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("01"))
      AND and_dcpl_28;
  and_dcpl_435 <= and_dcpl_433 AND and_dcpl_425;
  and_dcpl_436 <= and_dcpl_422 AND and_dcpl_425;
  and_dcpl_448 <= and_dcpl_33 AND and_dcpl_59 AND and_dcpl_28;
  and_dcpl_452 <= and_dcpl_33 AND and_dcpl_69 AND and_dcpl_35;
  and_dcpl_456 <= and_dcpl_365 AND and_dcpl_69 AND and_dcpl_28;
  and_dcpl_458 <= and_dcpl_365 AND and_dcpl_29 AND and_dcpl_35;
  and_dcpl_461 <= and_dcpl_372 AND and_dcpl_30;
  and_dcpl_465 <= and_dcpl_372 AND and_479_cse AND and_dcpl_50;
  and_dcpl_468 <= and_dcpl_372 AND and_479_cse AND (NOT (fsm_output(2))) AND (fsm_output(5));
  and_dcpl_472 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")) AND
      and_dcpl_31 AND and_dcpl_59 AND and_dcpl_50;
  and_dcpl_479 <= and_dcpl_353 AND and_dcpl_29 AND (fsm_output(2)) AND (NOT (fsm_output(5)));
  or_tmp_2098 <= (NOT (fsm_output(7))) OR (fsm_output(5)) OR (NOT or_212_cse);
  mux_1600_nl <= MUX_s_1_2_2(or_212_cse, (NOT or_212_cse), fsm_output(5));
  nand_520_nl <= NOT((fsm_output(7)) AND mux_1600_nl);
  mux_tmp_1564 <= MUX_s_1_2_2(nand_520_nl, or_tmp_2098, fsm_output(2));
  COMP_LOOP_or_33_itm <= and_605_cse OR and_609_cse OR and_614_cse OR and_617_cse
      OR and_621_cse OR and_624_cse OR and_628_cse;
  COMP_LOOP_tmp_or_71_itm <= and_dcpl_435 OR and_dcpl_436;
  COMP_LOOP_tmp_or_54_ssc <= and_dcpl_428 OR and_dcpl_429 OR and_dcpl_434;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((and_dcpl_33 AND and_dcpl_30) OR STAGE_LOOP_i_3_0_sva_mx0c1) = '1' )
          THEN
        STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "1010"), z_out_4,
            STAGE_LOOP_i_3_0_sva_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_1019_nl, mux_320_nl, fsm_output(5))) = '1' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_vec_rsc_triosy_0_31_obj_ld_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        COMP_LOOP_1_tmp_mul_idiv_sva_1_0 <= STD_LOGIC_VECTOR'( "00");
        COMP_LOOP_3_tmp_mul_idiv_sva_3_0 <= STD_LOGIC_VECTOR'( "0000");
      ELSE
        reg_vec_rsc_triosy_0_31_obj_ld_cse <= and_464_cse AND CONV_SL_1_1(fsm_output(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100100")) AND (NOT (z_out_2(4)));
        reg_ensig_cgo_cse <= mux_1462_rmff;
        COMP_LOOP_1_tmp_mul_idiv_sva_1_0 <= z_out_8(1 DOWNTO 0);
        COMP_LOOP_3_tmp_mul_idiv_sva_3_0 <= z_out_7(3 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      tmp_21_sva_2 <= twiddle_rsc_0_2_i_q_d;
      tmp_21_sva_6 <= twiddle_rsc_0_6_i_q_d;
      tmp_21_sva_11 <= MUX_v_64_2_2(twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_30_i_q_d,
          and_dcpl_176);
      tmp_21_sva_13 <= MUX_v_64_2_2(twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_6_i_q_d,
          and_dcpl_176);
      tmp_21_sva_14 <= MUX_v_64_2_2(twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_10_i_q_d,
          and_dcpl_176);
      tmp_21_sva_15 <= MUX_v_64_2_2(twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_14_i_q_d,
          and_dcpl_176);
      tmp_21_sva_17 <= MUX_v_64_2_2(twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d,
          and_dcpl_176);
      tmp_21_sva_18 <= twiddle_rsc_0_18_i_q_d;
      tmp_21_sva_22 <= twiddle_rsc_0_22_i_q_d;
      tmp_21_sva_26 <= twiddle_rsc_0_26_i_q_d;
      tmp_21_sva_30 <= twiddle_rsc_0_30_i_q_d;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_j_10_0_sva_9_0 <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (VEC_LOOP_j_10_0_sva_9_0_mx0c0 OR (and_dcpl_82 AND and_dcpl_104)) =
          '1' ) THEN
        VEC_LOOP_j_10_0_sva_9_0 <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"),
            (z_out_3(9 DOWNTO 0)), VEC_LOOP_j_not_1_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_1160_nl, and_nl, fsm_output(5))) = '1' ) THEN
        STAGE_LOOP_lshift_psp_sva <= z_out;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_1604_nl, mux_1603_nl, fsm_output(1))) = '1' ) THEN
        COMP_LOOP_k_10_3_sva_6_0 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), reg_COMP_LOOP_k_10_3_ftd,
            nand_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva <= COMP_LOOP_1_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_psp_sva <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_5_tmp_mul_idiv_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_5_tmp_mul_idiv_sva <= z_out_7(7 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm <= z_out_3(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_1_tmp_acc_cse_sva <= z_out_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_625_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_126_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_377_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_128_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_129_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_130_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_6_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_132_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_133_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_134_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_10_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_136_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_12_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_13_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_14_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_140_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_141_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_142_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_18_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_144_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_20_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_21_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_22_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_23_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_24_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_25_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_26_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_27_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_28_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_29_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_30_itm <= '0';
      ELSIF ( mux_1489_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_625_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
        COMP_LOOP_COMP_LOOP_and_126_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
        COMP_LOOP_COMP_LOOP_and_377_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
        COMP_LOOP_COMP_LOOP_and_128_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
        COMP_LOOP_COMP_LOOP_and_129_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
        COMP_LOOP_COMP_LOOP_and_130_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
        COMP_LOOP_COMP_LOOP_and_6_itm <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO
            0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("00"));
        COMP_LOOP_COMP_LOOP_and_132_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
        COMP_LOOP_COMP_LOOP_and_133_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
        COMP_LOOP_COMP_LOOP_and_134_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
        COMP_LOOP_COMP_LOOP_and_10_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(0)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1))
            OR (VEC_LOOP_j_10_0_sva_9_0(2))));
        COMP_LOOP_COMP_LOOP_and_136_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
        COMP_LOOP_COMP_LOOP_and_12_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(0)) AND (VEC_LOOP_j_10_0_sva_9_0(2))
            AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1))
            OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_13_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(0)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1))
            OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_14_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(0)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (NOT (COMP_LOOP_acc_psp_sva_mx0w0(1)));
        COMP_LOOP_COMP_LOOP_and_140_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10001"));
        COMP_LOOP_COMP_LOOP_and_141_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10010"));
        COMP_LOOP_COMP_LOOP_and_142_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10011"));
        COMP_LOOP_COMP_LOOP_and_18_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(1)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0))
            OR (VEC_LOOP_j_10_0_sva_9_0(2))));
        COMP_LOOP_COMP_LOOP_and_144_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10101"));
        COMP_LOOP_COMP_LOOP_and_20_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(1)) AND (VEC_LOOP_j_10_0_sva_9_0(2))
            AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0))
            OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_21_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(1)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0))
            OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_22_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(1)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (NOT (COMP_LOOP_acc_psp_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_23_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("000"));
        COMP_LOOP_COMP_LOOP_and_24_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("001"));
        COMP_LOOP_COMP_LOOP_and_25_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("010"));
        COMP_LOOP_COMP_LOOP_and_26_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("011"));
        COMP_LOOP_COMP_LOOP_and_27_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("100"));
        COMP_LOOP_COMP_LOOP_and_28_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("101"));
        COMP_LOOP_COMP_LOOP_and_29_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("110"));
        COMP_LOOP_COMP_LOOP_and_30_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_1459, mux_1492_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_6_sva <= COMP_LOOP_acc_1_cse_6_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_1497_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_4_sva <= COMP_LOOP_acc_1_cse_4_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_1499_nl AND nor_1025_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_1500_nl AND nor_1025_cse)) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_2_sva <= COMP_LOOP_2_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(mux_1502_nl AND nor_1025_cse)) = '1' ) THEN
        COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_3_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_5_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_5_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_126_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_126_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_127_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_127_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_157_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_157_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_129_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_129_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_159_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_159_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_160_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_160_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_161_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_161_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_133_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_133_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_163_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_163_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_164_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_164_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_165_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_165_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_166_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_166_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_167_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_167_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_168_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_168_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_169_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_169_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_140_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_nor_140_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_171_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_171_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_172_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_172_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_173_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_173_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_174_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_174_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_175_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_175_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_176_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_176_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_177_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_177_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_178_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_178_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_179_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_179_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_180_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_180_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_181_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_181_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_182_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_182_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_183_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_183_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_184_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_184_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_185_itm <= '0';
      ELSIF ( and_dcpl_252 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_185_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (mux_1505_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 1)) + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "01")),
            9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_3_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_1507_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_3_sva <= COMP_LOOP_3_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_1509_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm <= COMP_LOOP_acc_12_nl(8);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_9_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_9_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_226_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_nor_226_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_227_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_nor_227_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_281_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_281_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_229_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_nor_229_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_283_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_283_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_284_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_284_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_285_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_285_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_233_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_nor_233_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_287_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_287_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_288_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_288_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_289_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_289_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_290_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_290_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_291_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_291_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_292_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_292_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_293_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_293_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_240_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_nor_240_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_295_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_295_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_296_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_296_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_297_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_297_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_298_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_298_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_299_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_299_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_300_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_300_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_301_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_301_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_302_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_302_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_303_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_303_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_304_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_304_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_305_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_305_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_306_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_306_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_307_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_307_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_308_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_308_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_309_itm <= '0';
      ELSIF ( and_dcpl_256 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_309_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_1511_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_4_sva <= COMP_LOOP_4_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_1513_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_5_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_13_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_13_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_326_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_nor_326_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_327_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_nor_327_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_405_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_405_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_329_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_nor_329_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_407_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_407_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_408_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_408_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_409_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_409_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_333_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_nor_333_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_411_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_411_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_412_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_412_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_413_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_413_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_414_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_414_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_415_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_415_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_416_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_416_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_417_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_417_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_340_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_nor_340_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_419_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_419_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_420_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_420_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_421_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_421_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_422_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_422_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_423_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_423_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_424_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_424_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_425_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_425_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_426_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_426_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_427_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_427_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_428_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_428_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_429_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_429_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_430_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_430_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_431_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_431_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_432_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_432_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_433_itm <= '0';
      ELSIF ( and_dcpl_259 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_433_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (MUX_s_1_2_2(mux_1518_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 2)) + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & '1'), 8));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_5_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_1520_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_acc_10_cse_10_1_5_sva <= COMP_LOOP_5_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_1523_nl, (fsm_output(7)), fsm_output(5))) = '1' ) THEN
        COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_6_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_17_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_17_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_426_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_nor_426_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_427_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_nor_427_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_529_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_529_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_429_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_nor_429_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_531_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_531_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_532_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_532_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_533_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_533_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_433_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_nor_433_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_535_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_535_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_536_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_536_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_537_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_537_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_538_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_538_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_539_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_539_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_540_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_540_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_541_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_541_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_440_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_nor_440_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_543_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_543_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_544_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_544_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_545_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_545_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_546_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_546_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_547_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_547_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_548_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_548_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_549_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_549_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_550_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_550_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_551_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_551_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_552_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_552_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_553_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_553_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_554_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_554_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_555_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_555_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_556_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_556_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_557_itm <= '0';
      ELSIF ( and_dcpl_260 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_557_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm <= '0';
      ELSIF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_itm <= '0';
      ELSIF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_itm <= CONV_SL_1_1(z_out_7(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_itm <= '0';
      ELSIF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_itm <= CONV_SL_1_1(z_out_7(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_itm <= '0';
      ELSIF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_itm <= CONV_SL_1_1(z_out_7(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_itm <= '0';
      ELSIF ( or_dcpl_84 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_itm <= CONV_SL_1_1(z_out_7(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_1459, and_491_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_6_sva <= COMP_LOOP_6_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_tmp_1459, mux_1528_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_7_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_21_itm <= '0';
        COMP_LOOP_nor_526_itm <= '0';
        COMP_LOOP_nor_527_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_653_itm <= '0';
        COMP_LOOP_nor_529_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_655_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_656_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_657_itm <= '0';
        COMP_LOOP_nor_533_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_659_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_660_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_661_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_662_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_663_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_664_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_665_itm <= '0';
        COMP_LOOP_nor_540_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_667_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_668_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_669_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_670_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_671_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_672_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_673_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_674_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_675_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_676_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_677_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_678_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_679_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_680_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_681_itm <= '0';
      ELSIF ( mux_1531_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_21_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_nor_526_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_527_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_653_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
        COMP_LOOP_nor_529_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_655_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
        COMP_LOOP_COMP_LOOP_and_656_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
        COMP_LOOP_COMP_LOOP_and_657_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
        COMP_LOOP_nor_533_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_659_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
        COMP_LOOP_COMP_LOOP_and_660_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
        COMP_LOOP_COMP_LOOP_and_661_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
        COMP_LOOP_COMP_LOOP_and_662_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01100"));
        COMP_LOOP_COMP_LOOP_and_663_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
        COMP_LOOP_COMP_LOOP_and_664_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01110"));
        COMP_LOOP_COMP_LOOP_and_665_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
        COMP_LOOP_nor_540_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_COMP_LOOP_and_667_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10001"));
        COMP_LOOP_COMP_LOOP_and_668_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10010"));
        COMP_LOOP_COMP_LOOP_and_669_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10011"));
        COMP_LOOP_COMP_LOOP_and_670_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10100"));
        COMP_LOOP_COMP_LOOP_and_671_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10101"));
        COMP_LOOP_COMP_LOOP_and_672_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10110"));
        COMP_LOOP_COMP_LOOP_and_673_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
        COMP_LOOP_COMP_LOOP_and_674_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11000"));
        COMP_LOOP_COMP_LOOP_and_675_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11001"));
        COMP_LOOP_COMP_LOOP_and_676_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11010"));
        COMP_LOOP_COMP_LOOP_and_677_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
        COMP_LOOP_COMP_LOOP_and_678_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11100"));
        COMP_LOOP_COMP_LOOP_and_679_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
        COMP_LOOP_COMP_LOOP_and_680_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
        COMP_LOOP_COMP_LOOP_and_681_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (MUX_s_1_2_2(mux_1532_nl, and_464_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 1)) + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "11")),
            9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_7_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2((NOT or_tmp_2048), and_464_cse, or_162_nl)) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_7_sva <= COMP_LOOP_7_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_1536_itm = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm <= COMP_LOOP_acc_15_nl(7);
        reg_COMP_LOOP_k_10_3_ftd <= z_out_2(6 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_25_itm <= '0';
        COMP_LOOP_nor_626_itm <= '0';
        COMP_LOOP_nor_627_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_777_itm <= '0';
        COMP_LOOP_nor_629_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_779_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_780_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_781_itm <= '0';
        COMP_LOOP_nor_633_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_783_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_784_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_785_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_786_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_787_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_788_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_789_itm <= '0';
        COMP_LOOP_nor_640_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_791_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_792_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_793_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_794_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_795_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_796_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_797_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_798_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_799_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_800_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_801_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_802_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_803_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_804_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_805_itm <= '0';
      ELSIF ( mux_1538_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_25_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_nor_626_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_627_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_777_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
        COMP_LOOP_nor_629_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_779_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
        COMP_LOOP_COMP_LOOP_and_780_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
        COMP_LOOP_COMP_LOOP_and_781_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
        COMP_LOOP_nor_633_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_783_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
        COMP_LOOP_COMP_LOOP_and_784_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
        COMP_LOOP_COMP_LOOP_and_785_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
        COMP_LOOP_COMP_LOOP_and_786_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01100"));
        COMP_LOOP_COMP_LOOP_and_787_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
        COMP_LOOP_COMP_LOOP_and_788_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01110"));
        COMP_LOOP_COMP_LOOP_and_789_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
        COMP_LOOP_nor_640_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_COMP_LOOP_and_791_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10001"));
        COMP_LOOP_COMP_LOOP_and_792_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10010"));
        COMP_LOOP_COMP_LOOP_and_793_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10011"));
        COMP_LOOP_COMP_LOOP_and_794_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10100"));
        COMP_LOOP_COMP_LOOP_and_795_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10101"));
        COMP_LOOP_COMP_LOOP_and_796_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10110"));
        COMP_LOOP_COMP_LOOP_and_797_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
        COMP_LOOP_COMP_LOOP_and_798_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11000"));
        COMP_LOOP_COMP_LOOP_and_799_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11001"));
        COMP_LOOP_COMP_LOOP_and_800_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11010"));
        COMP_LOOP_COMP_LOOP_and_801_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
        COMP_LOOP_COMP_LOOP_and_802_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11100"));
        COMP_LOOP_COMP_LOOP_and_803_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
        COMP_LOOP_COMP_LOOP_and_804_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
        COMP_LOOP_COMP_LOOP_and_805_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_717, and_305_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "111")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_717, and_464_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_sva <= COMP_LOOP_8_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(not_tmp_717, and_304_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_1_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_29_itm <= '0';
        COMP_LOOP_nor_726_itm <= '0';
        COMP_LOOP_nor_727_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_901_itm <= '0';
        COMP_LOOP_nor_729_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_903_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_904_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_905_itm <= '0';
        COMP_LOOP_nor_733_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_907_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_908_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_909_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_910_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_911_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_912_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_913_itm <= '0';
        COMP_LOOP_nor_740_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_915_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_916_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_917_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_918_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_919_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_920_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_921_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_922_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_923_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_924_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_925_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_926_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_927_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_928_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_929_itm <= '0';
      ELSIF ( mux_1543_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_29_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_nor_726_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_727_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_901_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00011"));
        COMP_LOOP_nor_729_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_903_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00101"));
        COMP_LOOP_COMP_LOOP_and_904_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00110"));
        COMP_LOOP_COMP_LOOP_and_905_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("00111"));
        COMP_LOOP_nor_733_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_907_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01001"));
        COMP_LOOP_COMP_LOOP_and_908_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01010"));
        COMP_LOOP_COMP_LOOP_and_909_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01011"));
        COMP_LOOP_COMP_LOOP_and_910_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01100"));
        COMP_LOOP_COMP_LOOP_and_911_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01101"));
        COMP_LOOP_COMP_LOOP_and_912_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01110"));
        COMP_LOOP_COMP_LOOP_and_913_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
        COMP_LOOP_nor_740_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_COMP_LOOP_and_915_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10001"));
        COMP_LOOP_COMP_LOOP_and_916_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10010"));
        COMP_LOOP_COMP_LOOP_and_917_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10011"));
        COMP_LOOP_COMP_LOOP_and_918_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10100"));
        COMP_LOOP_COMP_LOOP_and_919_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10101"));
        COMP_LOOP_COMP_LOOP_and_920_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10110"));
        COMP_LOOP_COMP_LOOP_and_921_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
        COMP_LOOP_COMP_LOOP_and_922_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11000"));
        COMP_LOOP_COMP_LOOP_and_923_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11001"));
        COMP_LOOP_COMP_LOOP_and_924_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11010"));
        COMP_LOOP_COMP_LOOP_and_925_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
        COMP_LOOP_COMP_LOOP_and_926_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11100"));
        COMP_LOOP_COMP_LOOP_and_927_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
        COMP_LOOP_COMP_LOOP_and_928_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
        COMP_LOOP_COMP_LOOP_and_929_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_33_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_35_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_36_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_37_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_39_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_40_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_41_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_42_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_43_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_44_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_45_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_47_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & and_dcpl_49 & and_dcpl_171 & COMP_LOOP_or_59_cse
            & and_dcpl_173));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm <= '0';
        COMP_LOOP_tmp_nor_1_itm <= '0';
        COMP_LOOP_tmp_nor_14_itm <= '0';
        COMP_LOOP_tmp_nor_3_itm <= '0';
        COMP_LOOP_tmp_nor_42_itm <= '0';
        COMP_LOOP_tmp_nor_49_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_12_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_48_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & COMP_LOOP_or_59_cse & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_49_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & COMP_LOOP_or_59_cse & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_50_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & COMP_LOOP_or_59_cse & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_51_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & COMP_LOOP_or_59_cse & and_dcpl_173));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_52_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & COMP_LOOP_or_59_cse & and_dcpl_173));
        COMP_LOOP_tmp_nor_1_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_26_nl, COMP_LOOP_tmp_nor_1_cse,
            COMP_LOOP_tmp_nor_35_cse, COMP_LOOP_tmp_nor_101_cse, STD_LOGIC_VECTOR'(
            and_dcpl_46 & and_dcpl_49 & COMP_LOOP_or_41_cse & and_dcpl_176));
        COMP_LOOP_tmp_nor_14_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_27_nl, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse,
            COMP_LOOP_tmp_nor_1_cse, COMP_LOOP_tmp_nor_105_cse, STD_LOGIC_VECTOR'(
            and_dcpl_46 & and_dcpl_49 & COMP_LOOP_or_41_cse & and_dcpl_176));
        COMP_LOOP_tmp_nor_3_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_nor_29_nl, COMP_LOOP_tmp_nor_101_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & COMP_LOOP_or_39_cse & and_dcpl_176));
        COMP_LOOP_tmp_nor_42_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_nor_33_nl, COMP_LOOP_tmp_nor_105_cse,
            COMP_LOOP_tmp_nor_35_cse, STD_LOGIC_VECTOR'( and_dcpl_46 & COMP_LOOP_or_39_cse
            & and_dcpl_176));
        COMP_LOOP_tmp_nor_49_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_40_nl, COMP_LOOP_tmp_nor_35_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse, COMP_LOOP_tmp_nor_1_cse, STD_LOGIC_VECTOR'(
            and_dcpl_46 & and_dcpl_49 & COMP_LOOP_or_41_cse & and_dcpl_176));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_17_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_53_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_54_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_55_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_56_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_57_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_58_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_59_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_60_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_61_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse, STD_LOGIC_VECTOR'( and_dcpl_46
            & and_dcpl_49 & and_dcpl_172 & and_dcpl_174));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_nor_1_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse,
            STD_LOGIC_VECTOR'( and_dcpl_46 & COMP_LOOP_or_42_cse & and_dcpl_174));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_mux1h_itm_mx0c0 OR COMP_LOOP_tmp_mux1h_itm_mx0c1 OR COMP_LOOP_tmp_mux1h_itm_mx0c2
          OR COMP_LOOP_tmp_mux1h_itm_mx0c3) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_itm <= MUX1HOT_v_64_4_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_8_i_q_d,
            twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_24_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_mux1h_itm_mx0c0
            & COMP_LOOP_tmp_mux1h_itm_mx0c1 & COMP_LOOP_tmp_mux1h_itm_mx0c2 & COMP_LOOP_tmp_mux1h_itm_mx0c3));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_2_tmp_mul_idiv_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( COMP_LOOP_or_39_cse = '1' ) THEN
        COMP_LOOP_2_tmp_mul_idiv_sva <= z_out_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_2_tmp_lshift_ncse_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (and_dcpl_49 OR and_dcpl_176) = '1' ) THEN
        COMP_LOOP_2_tmp_lshift_ncse_sva <= MUX_v_10_2_2(z_out_1, z_out_7, and_dcpl_176);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_49 OR and_dcpl_171 OR and_dcpl_278 OR and_dcpl_176 OR COMP_LOOP_1_acc_8_itm_mx0c4
          OR and_dcpl_54 OR and_dcpl_222 OR and_dcpl_58 OR and_dcpl_226 OR and_dcpl_65
          OR and_dcpl_229 OR and_dcpl_68 OR and_dcpl_232 OR and_dcpl_75 OR and_dcpl_234
          OR and_dcpl_78 OR and_dcpl_236 OR and_dcpl_83 OR and_dcpl_238) = '1' )
          THEN
        COMP_LOOP_1_acc_8_itm <= MUX1HOT_v_64_36_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
            vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
            vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
            vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
            vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, vec_rsc_0_16_i_q_d, vec_rsc_0_17_i_q_d,
            vec_rsc_0_18_i_q_d, vec_rsc_0_19_i_q_d, vec_rsc_0_20_i_q_d, vec_rsc_0_21_i_q_d,
            vec_rsc_0_22_i_q_d, vec_rsc_0_23_i_q_d, vec_rsc_0_24_i_q_d, vec_rsc_0_25_i_q_d,
            vec_rsc_0_26_i_q_d, vec_rsc_0_27_i_q_d, vec_rsc_0_28_i_q_d, vec_rsc_0_29_i_q_d,
            vec_rsc_0_30_i_q_d, vec_rsc_0_31_i_q_d, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_acc_17_nl),
            64)), twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_26_i_q_d, COMP_LOOP_1_modulo_dev_cmp_return_rsc_z,
            STD_LOGIC_VECTOR'( COMP_LOOP_or_nl & COMP_LOOP_or_1_nl & COMP_LOOP_or_2_nl
            & COMP_LOOP_or_3_nl & COMP_LOOP_or_4_nl & COMP_LOOP_or_5_nl & COMP_LOOP_or_6_nl
            & COMP_LOOP_or_7_nl & COMP_LOOP_or_8_nl & COMP_LOOP_or_9_nl & COMP_LOOP_or_10_nl
            & COMP_LOOP_or_11_nl & COMP_LOOP_or_12_nl & COMP_LOOP_or_13_nl & COMP_LOOP_or_14_nl
            & COMP_LOOP_or_15_nl & COMP_LOOP_or_16_nl & COMP_LOOP_or_17_nl & COMP_LOOP_or_18_nl
            & COMP_LOOP_or_19_nl & COMP_LOOP_or_20_nl & COMP_LOOP_or_21_nl & COMP_LOOP_or_22_nl
            & COMP_LOOP_or_23_nl & COMP_LOOP_or_24_nl & COMP_LOOP_or_25_nl & COMP_LOOP_or_26_nl
            & COMP_LOOP_or_27_nl & COMP_LOOP_or_28_nl & COMP_LOOP_or_29_nl & COMP_LOOP_or_30_nl
            & COMP_LOOP_or_31_nl & COMP_LOOP_or_36_itm & and_dcpl_278 & and_dcpl_176
            & COMP_LOOP_1_acc_8_itm_mx0c4));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_3_tmp_lshift_ncse_sva <= STD_LOGIC_VECTOR'( "000000000");
        COMP_LOOP_tmp_nor_25_itm <= '0';
        COMP_LOOP_tmp_nor_26_itm <= '0';
        COMP_LOOP_tmp_nor_28_itm <= '0';
        COMP_LOOP_tmp_nor_31_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_35_cse = '1' ) THEN
        COMP_LOOP_3_tmp_lshift_ncse_sva <= MUX_v_9_2_2((z_out_1(8 DOWNTO 0)), (z_out_7(8
            DOWNTO 0)), and_dcpl_174);
        COMP_LOOP_tmp_nor_25_itm <= COMP_LOOP_tmp_nor_78_cse;
        COMP_LOOP_tmp_nor_26_itm <= COMP_LOOP_tmp_nor_79_cse;
        COMP_LOOP_tmp_nor_28_itm <= COMP_LOOP_tmp_nor_81_cse;
        COMP_LOOP_tmp_nor_31_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_294_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_1_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
            twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d,
            twiddle_rsc_0_5_i_q_d, twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d,
            twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_9_i_q_d, twiddle_rsc_0_10_i_q_d,
            twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_13_i_q_d,
            twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_16_i_q_d,
            twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_19_i_q_d,
            twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_21_i_q_d, twiddle_rsc_0_22_i_q_d,
            twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_25_i_q_d,
            twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_27_i_q_d, twiddle_rsc_0_28_i_q_d,
            twiddle_rsc_0_29_i_q_d, twiddle_rsc_0_30_i_q_d, twiddle_rsc_0_31_i_q_d,
            STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_127_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl & COMP_LOOP_tmp_and_128_nl & COMP_LOOP_tmp_and_129_nl
            & COMP_LOOP_tmp_and_130_nl & COMP_LOOP_tmp_and_131_nl & COMP_LOOP_tmp_and_132_nl
            & COMP_LOOP_tmp_and_133_nl & COMP_LOOP_tmp_and_134_nl & COMP_LOOP_tmp_and_135_nl
            & COMP_LOOP_tmp_and_136_nl & COMP_LOOP_tmp_and_137_nl & COMP_LOOP_tmp_and_138_nl
            & COMP_LOOP_tmp_and_139_nl & COMP_LOOP_tmp_and_140_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_nl
            & COMP_LOOP_tmp_and_141_nl & COMP_LOOP_tmp_and_142_nl & COMP_LOOP_tmp_and_143_nl
            & COMP_LOOP_tmp_and_144_nl & COMP_LOOP_tmp_and_145_nl & COMP_LOOP_tmp_and_146_nl
            & COMP_LOOP_tmp_and_147_nl & COMP_LOOP_tmp_and_148_nl & COMP_LOOP_tmp_and_149_nl
            & COMP_LOOP_tmp_and_150_nl & COMP_LOOP_tmp_and_151_nl & COMP_LOOP_tmp_and_152_nl
            & COMP_LOOP_tmp_and_153_nl & COMP_LOOP_tmp_and_154_nl & COMP_LOOP_tmp_and_155_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( nor_1119_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_2_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_2_i_q_d,
            twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_8_i_q_d,
            twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_14_i_q_d,
            twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_20_i_q_d,
            twiddle_rsc_0_22_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_26_i_q_d,
            twiddle_rsc_0_28_i_q_d, twiddle_rsc_0_30_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_115_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_nl
            & COMP_LOOP_tmp_and_116_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_nl &
            COMP_LOOP_tmp_and_117_nl & COMP_LOOP_tmp_and_118_nl & COMP_LOOP_tmp_and_119_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_nl & COMP_LOOP_tmp_and_120_nl &
            COMP_LOOP_tmp_and_121_nl & COMP_LOOP_tmp_and_122_nl & COMP_LOOP_tmp_and_123_nl
            & COMP_LOOP_tmp_and_124_nl & COMP_LOOP_tmp_and_125_nl & COMP_LOOP_tmp_and_126_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( nor_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_3_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
            twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d,
            twiddle_rsc_0_5_i_q_d, twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d,
            twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_9_i_q_d, twiddle_rsc_0_10_i_q_d,
            twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_13_i_q_d,
            twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_16_i_q_d,
            twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_19_i_q_d,
            twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_21_i_q_d, twiddle_rsc_0_22_i_q_d,
            twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_25_i_q_d,
            twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_27_i_q_d, twiddle_rsc_0_28_i_q_d,
            twiddle_rsc_0_29_i_q_d, twiddle_rsc_0_30_i_q_d, twiddle_rsc_0_31_i_q_d,
            STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_83_nl & COMP_LOOP_tmp_and_84_nl
            & COMP_LOOP_tmp_and_85_nl & COMP_LOOP_tmp_and_86_nl & COMP_LOOP_tmp_and_87_nl
            & COMP_LOOP_tmp_and_88_nl & COMP_LOOP_tmp_and_89_nl & COMP_LOOP_tmp_and_90_nl
            & COMP_LOOP_tmp_and_91_nl & COMP_LOOP_tmp_and_92_nl & COMP_LOOP_tmp_and_93_nl
            & COMP_LOOP_tmp_and_94_nl & COMP_LOOP_tmp_and_95_nl & COMP_LOOP_tmp_and_96_nl
            & COMP_LOOP_tmp_and_97_nl & COMP_LOOP_tmp_and_98_nl & COMP_LOOP_tmp_and_99_nl
            & COMP_LOOP_tmp_and_100_nl & COMP_LOOP_tmp_and_101_nl & COMP_LOOP_tmp_and_102_nl
            & COMP_LOOP_tmp_and_103_nl & COMP_LOOP_tmp_and_104_nl & COMP_LOOP_tmp_and_105_nl
            & COMP_LOOP_tmp_and_106_nl & COMP_LOOP_tmp_and_107_nl & COMP_LOOP_tmp_and_108_nl
            & COMP_LOOP_tmp_and_109_nl & COMP_LOOP_tmp_and_110_nl & COMP_LOOP_tmp_and_111_nl
            & COMP_LOOP_tmp_and_112_nl & COMP_LOOP_tmp_and_113_nl & COMP_LOOP_tmp_and_114_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_40_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse;
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_cse, and_dcpl_176);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse, and_dcpl_176);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_cse, and_dcpl_176);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_cse, and_dcpl_176);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_cse, and_dcpl_176);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_cse, and_dcpl_176);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_cse, and_dcpl_176);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_cse, and_dcpl_176);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_cse, and_dcpl_176);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( nor_1117_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_4_itm <= MUX1HOT_v_64_8_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_4_i_q_d,
            twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_16_i_q_d,
            twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_28_i_q_d,
            STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_78_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_nl & COMP_LOOP_tmp_and_79_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_nl
            & COMP_LOOP_tmp_and_80_nl & COMP_LOOP_tmp_and_81_nl & COMP_LOOP_tmp_and_82_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (((NOT((COMP_LOOP_2_tmp_lshift_ncse_sva(0)) AND COMP_LOOP_tmp_nor_42_itm))
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm OR and_dcpl_278 OR and_dcpl_176)
          AND mux_1585_nl) = '1' ) THEN
        tmp_21_sva_1 <= MUX1HOT_v_64_33_2(twiddle_rsc_0_1_i_q_d, twiddle_rsc_0_22_i_q_d,
            twiddle_rsc_0_0_i_q_d, tmp_21_sva_2, tmp_21_sva_3, twiddle_rsc_0_4_i_q_d,
            tmp_21_sva_5, tmp_21_sva_6, tmp_21_sva_7, twiddle_rsc_0_8_i_q_d, tmp_21_sva_9,
            COMP_LOOP_1_acc_8_itm, tmp_21_sva_11, twiddle_rsc_0_12_i_q_d, tmp_21_sva_13,
            tmp_21_sva_14, tmp_21_sva_15, twiddle_rsc_0_16_i_q_d, tmp_21_sva_17,
            tmp_21_sva_18, tmp_21_sva_19, twiddle_rsc_0_20_i_q_d, tmp_21_sva_21,
            tmp_21_sva_22, tmp_21_sva_23, twiddle_rsc_0_24_i_q_d, tmp_21_sva_25,
            tmp_21_sva_26, tmp_21_sva_27, twiddle_rsc_0_28_i_q_d, tmp_21_sva_29,
            tmp_21_sva_30, tmp_21_sva_31, STD_LOGIC_VECTOR'( and_dcpl_278 & and_dcpl_176
            & COMP_LOOP_tmp_and_47_nl & COMP_LOOP_tmp_and_48_nl & COMP_LOOP_tmp_and_49_nl
            & COMP_LOOP_tmp_and_50_nl & COMP_LOOP_tmp_and_51_nl & COMP_LOOP_tmp_and_52_nl
            & COMP_LOOP_tmp_and_53_nl & COMP_LOOP_tmp_and_54_nl & COMP_LOOP_tmp_and_55_nl
            & COMP_LOOP_tmp_and_56_nl & COMP_LOOP_tmp_and_57_nl & COMP_LOOP_tmp_and_58_nl
            & COMP_LOOP_tmp_and_59_nl & COMP_LOOP_tmp_and_60_nl & COMP_LOOP_tmp_and_61_nl
            & COMP_LOOP_tmp_and_62_nl & COMP_LOOP_tmp_and_63_nl & COMP_LOOP_tmp_and_64_nl
            & COMP_LOOP_tmp_and_65_nl & COMP_LOOP_tmp_and_66_nl & COMP_LOOP_tmp_and_67_nl
            & COMP_LOOP_tmp_and_68_nl & COMP_LOOP_tmp_and_69_nl & COMP_LOOP_tmp_and_70_nl
            & COMP_LOOP_tmp_and_71_nl & COMP_LOOP_tmp_and_72_nl & COMP_LOOP_tmp_and_73_nl
            & COMP_LOOP_tmp_and_74_nl & COMP_LOOP_tmp_and_75_nl & COMP_LOOP_tmp_and_76_nl
            & COMP_LOOP_tmp_and_77_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm)
          = '1' ) THEN
        tmp_21_sva_3 <= twiddle_rsc_0_3_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm)
          = '1' ) THEN
        tmp_21_sva_5 <= twiddle_rsc_0_5_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm)
          = '1' ) THEN
        tmp_21_sva_7 <= twiddle_rsc_0_7_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm)
          = '1' ) THEN
        tmp_21_sva_9 <= twiddle_rsc_0_9_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm)
          = '1' ) THEN
        tmp_21_sva_19 <= twiddle_rsc_0_19_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm)
          = '1' ) THEN
        tmp_21_sva_21 <= twiddle_rsc_0_21_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm)
          = '1' ) THEN
        tmp_21_sva_23 <= twiddle_rsc_0_23_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm)
          = '1' ) THEN
        tmp_21_sva_25 <= twiddle_rsc_0_25_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm)
          = '1' ) THEN
        tmp_21_sva_27 <= twiddle_rsc_0_27_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm)
          = '1' ) THEN
        tmp_21_sva_29 <= twiddle_rsc_0_29_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm)
          = '1' ) THEN
        tmp_21_sva_31 <= twiddle_rsc_0_31_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm <= '0';
      ELSIF ( or_dcpl_109 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm <= '0';
      ELSIF ( or_dcpl_109 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_1592_tmp = '1' ) THEN
        COMP_LOOP_tmp_mux1h_5_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_0_i_q_d, tmp_21_sva_1,
            tmp_21_sva_2, tmp_21_sva_3, twiddle_rsc_0_4_i_q_d, tmp_21_sva_5, tmp_21_sva_6,
            tmp_21_sva_7, twiddle_rsc_0_8_i_q_d, tmp_21_sva_9, COMP_LOOP_1_acc_8_itm,
            tmp_21_sva_11, twiddle_rsc_0_12_i_q_d, tmp_21_sva_13, tmp_21_sva_14,
            tmp_21_sva_15, twiddle_rsc_0_16_i_q_d, tmp_21_sva_17, tmp_21_sva_18,
            tmp_21_sva_19, twiddle_rsc_0_20_i_q_d, tmp_21_sva_21, tmp_21_sva_22,
            tmp_21_sva_23, twiddle_rsc_0_24_i_q_d, tmp_21_sva_25, tmp_21_sva_26,
            tmp_21_sva_27, twiddle_rsc_0_28_i_q_d, tmp_21_sva_29, tmp_21_sva_30,
            tmp_21_sva_31, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_15_nl & COMP_LOOP_tmp_and_16_nl
            & COMP_LOOP_tmp_and_17_nl & COMP_LOOP_tmp_and_18_nl & COMP_LOOP_tmp_and_19_nl
            & COMP_LOOP_tmp_and_20_nl & COMP_LOOP_tmp_and_21_nl & COMP_LOOP_tmp_and_22_nl
            & COMP_LOOP_tmp_and_23_nl & COMP_LOOP_tmp_and_24_nl & COMP_LOOP_tmp_and_25_nl
            & COMP_LOOP_tmp_and_26_nl & COMP_LOOP_tmp_and_27_nl & COMP_LOOP_tmp_and_28_nl
            & COMP_LOOP_tmp_and_29_nl & COMP_LOOP_tmp_and_30_nl & COMP_LOOP_tmp_and_31_nl
            & COMP_LOOP_tmp_and_32_nl & COMP_LOOP_tmp_and_33_nl & COMP_LOOP_tmp_and_34_nl
            & COMP_LOOP_tmp_and_35_nl & COMP_LOOP_tmp_and_36_nl & COMP_LOOP_tmp_and_37_nl
            & COMP_LOOP_tmp_and_38_nl & COMP_LOOP_tmp_and_39_nl & COMP_LOOP_tmp_and_40_nl
            & COMP_LOOP_tmp_and_41_nl & COMP_LOOP_tmp_and_42_nl & COMP_LOOP_tmp_and_43_nl
            & COMP_LOOP_tmp_and_44_nl & COMP_LOOP_tmp_and_45_nl & COMP_LOOP_tmp_and_46_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (((NOT((COMP_LOOP_3_tmp_lshift_ncse_sva(0)) AND COMP_LOOP_tmp_nor_25_itm))
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_119_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_121_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_125_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm OR and_dcpl_176) AND mux_1597_nl)
          = '1' ) THEN
        COMP_LOOP_tmp_mux1h_6_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_0_i_q_d,
            twiddle_rsc_0_4_i_q_d, tmp_21_sva_13, twiddle_rsc_0_8_i_q_d, tmp_21_sva_14,
            twiddle_rsc_0_12_i_q_d, tmp_21_sva_15, twiddle_rsc_0_16_i_q_d, tmp_21_sva_17,
            twiddle_rsc_0_20_i_q_d, tmp_21_sva_1, twiddle_rsc_0_24_i_q_d, COMP_LOOP_1_acc_8_itm,
            twiddle_rsc_0_28_i_q_d, tmp_21_sva_11, STD_LOGIC_VECTOR'( and_dcpl_176
            & COMP_LOOP_tmp_and_nl & COMP_LOOP_tmp_and_1_nl & COMP_LOOP_tmp_and_2_nl
            & COMP_LOOP_tmp_and_3_nl & COMP_LOOP_tmp_and_4_nl & COMP_LOOP_tmp_and_5_nl
            & COMP_LOOP_tmp_and_6_nl & COMP_LOOP_tmp_and_7_nl & COMP_LOOP_tmp_and_8_nl
            & COMP_LOOP_tmp_and_9_nl & COMP_LOOP_tmp_and_10_nl & COMP_LOOP_tmp_and_11_nl
            & COMP_LOOP_tmp_and_12_nl & COMP_LOOP_tmp_and_13_nl & COMP_LOOP_tmp_and_14_nl));
      END IF;
    END IF;
  END PROCESS;
  nor_1019_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(0))
      OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(7)));
  mux_320_nl <= MUX_s_1_2_2(and_33_cse, nor_tmp_95, fsm_output(2));
  VEC_LOOP_j_not_1_nl <= NOT VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  nor_1160_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(1))
      OR (fsm_output(6)) OR (fsm_output(7)));
  and_nl <= or_220_cse AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  nor_1021_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(7)));
  and_451_nl <= (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(7));
  mux_312_nl <= MUX_s_1_2_2(nor_1021_nl, and_451_nl, fsm_output(5));
  nand_nl <= NOT(mux_312_nl AND and_dcpl_244 AND nor_1023_cse);
  or_2285_nl <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(4))
      OR (fsm_output(3));
  mux_1604_nl <= MUX_s_1_2_2(or_2285_nl, mux_tmp_1564, fsm_output(6));
  or_2284_nl <= (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(4)) OR (fsm_output(3));
  or_nl <= (NOT (fsm_output(7))) OR (fsm_output(5));
  mux_nl <= MUX_s_1_2_2(or_tmp_2098, or_nl, fsm_output(2));
  mux_1602_nl <= MUX_s_1_2_2(mux_tmp_1564, mux_nl, fsm_output(0));
  mux_1603_nl <= MUX_s_1_2_2(or_2284_nl, mux_1602_nl, fsm_output(6));
  mux_1492_nl <= MUX_s_1_2_2(mux_tmp_1456, and_491_cse, fsm_output(2));
  mux_1496_nl <= MUX_s_1_2_2(and_tmp_11, and_485_cse, fsm_output(2));
  mux_1497_nl <= MUX_s_1_2_2(not_tmp_692, mux_1496_nl, fsm_output(5));
  and_260_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND or_32_cse;
  mux_1498_nl <= MUX_s_1_2_2(and_260_nl, and_479_cse, fsm_output(2));
  mux_1499_nl <= MUX_s_1_2_2(or_tmp_2057, (NOT mux_1498_nl), fsm_output(5));
  mux_1500_nl <= MUX_s_1_2_2(or_tmp_2057, (NOT and_479_cse), fsm_output(5));
  COMP_LOOP_3_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & STD_LOGIC_VECTOR'( "010")), 10), 11) + SIGNED'( "00000000001"), 11));
  and_310_nl <= (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(1));
  mux_1501_nl <= MUX_s_1_2_2(and_310_nl, and_479_cse, fsm_output(2));
  mux_1502_nl <= MUX_s_1_2_2(or_tmp_2057, (NOT mux_1501_nl), fsm_output(5));
  mux_1504_nl <= MUX_s_1_2_2(mux_tmp_1468, and_tmp_11, fsm_output(2));
  mux_1505_nl <= MUX_s_1_2_2(mux_1504_nl, (fsm_output(6)), fsm_output(5));
  mux_1506_nl <= MUX_s_1_2_2(mux_tmp_1468, and_485_cse, fsm_output(2));
  mux_1507_nl <= MUX_s_1_2_2(mux_1506_nl, (fsm_output(6)), fsm_output(5));
  COMP_LOOP_acc_12_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 3)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & '0'), 8), 9) + UNSIGNED'( "000000001"), 9));
  mux_1508_nl <= MUX_s_1_2_2(mux_tmp_1468, and_tmp_13, fsm_output(2));
  mux_1509_nl <= MUX_s_1_2_2(mux_1508_nl, (fsm_output(6)), fsm_output(5));
  mux_1511_nl <= MUX_s_1_2_2(not_tmp_692, and_485_cse, fsm_output(5));
  COMP_LOOP_5_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & STD_LOGIC_VECTOR'( "100")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_1512_nl <= MUX_s_1_2_2(and_tmp_13, and_485_cse, fsm_output(2));
  mux_1513_nl <= MUX_s_1_2_2(not_tmp_692, mux_1512_nl, fsm_output(5));
  mux_1518_nl <= MUX_s_1_2_2(mux_tmp_1482, mux_tmp_1456, fsm_output(2));
  mux_1520_nl <= MUX_s_1_2_2(mux_tmp_1482, and_491_cse, fsm_output(2));
  COMP_LOOP_6_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & STD_LOGIC_VECTOR'( "101")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_1523_nl <= MUX_s_1_2_2(mux_tmp_1482, mux_tmp_1487, fsm_output(2));
  COMP_LOOP_7_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & STD_LOGIC_VECTOR'( "110")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_1528_nl <= MUX_s_1_2_2(mux_tmp_1487, and_491_cse, fsm_output(2));
  mux_1532_nl <= MUX_s_1_2_2(mux_tmp_1452, nor_tmp_95, fsm_output(2));
  or_162_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("0000"));
  COMP_LOOP_acc_15_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 4)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0),
      7), 8) + UNSIGNED'( "00000001"), 8));
  and_305_nl <= (CONV_SL_1_1(fsm_output(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  COMP_LOOP_1_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(z_out_2 & STD_LOGIC_VECTOR'(
      "000")) + SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10 DOWNTO 1)))) + SIGNED'(
      "00000000001"), 11));
  and_304_nl <= (CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  COMP_LOOP_COMP_LOOP_and_33_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("00011"));
  COMP_LOOP_COMP_LOOP_and_35_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("00101"));
  COMP_LOOP_COMP_LOOP_and_36_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("00110"));
  COMP_LOOP_COMP_LOOP_and_37_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("00111"));
  COMP_LOOP_COMP_LOOP_and_39_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("01001"));
  COMP_LOOP_COMP_LOOP_and_40_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("01010"));
  COMP_LOOP_COMP_LOOP_and_41_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("01011"));
  COMP_LOOP_COMP_LOOP_and_42_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("01100"));
  COMP_LOOP_COMP_LOOP_and_43_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("01101"));
  COMP_LOOP_COMP_LOOP_and_44_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("01110"));
  COMP_LOOP_COMP_LOOP_and_45_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("01111"));
  COMP_LOOP_COMP_LOOP_and_47_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("10001"));
  COMP_LOOP_COMP_LOOP_and_48_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("10010"));
  COMP_LOOP_COMP_LOOP_and_49_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("10011"));
  COMP_LOOP_COMP_LOOP_and_50_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("10100"));
  COMP_LOOP_COMP_LOOP_and_51_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("10101"));
  COMP_LOOP_COMP_LOOP_and_52_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("10110"));
  COMP_LOOP_nor_26_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
  COMP_LOOP_nor_27_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(3))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_29_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(3))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_33_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(2))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_40_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
  COMP_LOOP_COMP_LOOP_and_53_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("10111"));
  COMP_LOOP_COMP_LOOP_and_54_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("11000"));
  COMP_LOOP_COMP_LOOP_and_55_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("11001"));
  COMP_LOOP_COMP_LOOP_and_56_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("11010"));
  COMP_LOOP_COMP_LOOP_and_57_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("11011"));
  COMP_LOOP_COMP_LOOP_and_58_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("11100"));
  COMP_LOOP_COMP_LOOP_and_59_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("11101"));
  COMP_LOOP_COMP_LOOP_and_60_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("11110"));
  COMP_LOOP_COMP_LOOP_and_61_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO
      0)=STD_LOGIC_VECTOR'("11111"));
  COMP_LOOP_COMP_LOOP_nor_1_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
  COMP_LOOP_COMP_LOOP_mux_2_nl <= MUX_v_64_2_2(COMP_LOOP_1_acc_8_itm, z_out_9, COMP_LOOP_or_33_itm);
  COMP_LOOP_acc_17_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_385_cse)
      + UNSIGNED(COMP_LOOP_COMP_LOOP_mux_2_nl), 64));
  COMP_LOOP_or_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm AND and_dcpl_49) OR
      (COMP_LOOP_COMP_LOOP_and_30_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_29_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_28_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_27_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_26_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_25_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_24_itm AND and_dcpl_83);
  COMP_LOOP_or_1_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(0)) AND COMP_LOOP_tmp_nor_1_itm
      AND and_dcpl_49) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_29_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_28_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_27_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_26_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_25_itm AND and_dcpl_83);
  COMP_LOOP_or_2_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(1)) AND COMP_LOOP_tmp_nor_14_itm
      AND and_dcpl_49) OR (COMP_LOOP_COMP_LOOP_and_625_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_29_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_28_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_27_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_26_itm AND and_dcpl_83);
  COMP_LOOP_or_3_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_126_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_625_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_29_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_28_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_27_itm AND and_dcpl_83);
  COMP_LOOP_or_4_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(2)) AND COMP_LOOP_tmp_nor_3_itm
      AND and_dcpl_49) OR (COMP_LOOP_COMP_LOOP_and_377_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_126_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_625_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_29_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_28_itm AND and_dcpl_83);
  COMP_LOOP_or_5_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_128_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_377_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_126_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_625_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_29_itm AND and_dcpl_83);
  COMP_LOOP_or_6_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_129_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_128_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_377_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_126_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_625_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_dcpl_83);
  COMP_LOOP_or_7_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_130_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_129_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_128_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_377_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_126_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_625_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_83);
  COMP_LOOP_or_8_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(3)) AND COMP_LOOP_tmp_nor_42_itm
      AND and_dcpl_49) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_130_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_129_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_128_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_377_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_126_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_625_itm AND and_dcpl_83);
  COMP_LOOP_or_9_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_132_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_130_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_129_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_128_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_377_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_126_itm AND and_dcpl_83);
  COMP_LOOP_or_10_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_133_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_132_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_130_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_129_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_128_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_377_itm AND and_dcpl_83);
  COMP_LOOP_or_11_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_134_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_133_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_132_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_130_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_129_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_128_itm AND and_dcpl_83);
  COMP_LOOP_or_12_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_134_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_133_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_132_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_130_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_129_itm AND and_dcpl_83);
  COMP_LOOP_or_13_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_136_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_134_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_133_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_132_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_130_itm AND and_dcpl_83);
  COMP_LOOP_or_14_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_136_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_134_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_133_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_132_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_83);
  COMP_LOOP_or_15_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_136_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_134_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_133_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_132_itm AND and_dcpl_83);
  COMP_LOOP_or_16_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(4)) AND COMP_LOOP_tmp_nor_49_itm
      AND and_dcpl_49) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_136_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_134_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_133_itm AND and_dcpl_83);
  COMP_LOOP_or_17_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_140_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_136_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_134_itm AND and_dcpl_83);
  COMP_LOOP_or_18_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_141_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_140_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_136_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_83);
  COMP_LOOP_or_19_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_142_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_141_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_140_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_136_itm AND and_dcpl_83);
  COMP_LOOP_or_20_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_18_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_142_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_141_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_140_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_83);
  COMP_LOOP_or_21_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_144_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_18_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_142_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_141_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_140_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_83);
  COMP_LOOP_or_22_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_20_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_144_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_18_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_142_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_141_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_140_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_83);
  COMP_LOOP_or_23_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_21_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_20_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_144_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_18_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_142_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_141_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_140_itm AND and_dcpl_83);
  COMP_LOOP_or_24_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_22_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_21_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_20_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_144_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_18_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_142_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_141_itm AND and_dcpl_83);
  COMP_LOOP_or_25_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_23_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_22_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_21_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_20_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_144_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_18_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_142_itm AND and_dcpl_83);
  COMP_LOOP_or_26_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_24_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_23_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_22_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_21_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_20_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_144_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_18_itm AND and_dcpl_83);
  COMP_LOOP_or_27_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_25_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_24_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_23_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_22_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_21_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_20_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_144_itm AND and_dcpl_83);
  COMP_LOOP_or_28_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_26_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_25_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_24_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_23_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_22_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_21_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_20_itm AND and_dcpl_83);
  COMP_LOOP_or_29_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_27_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_26_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_25_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_24_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_23_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_22_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_21_itm AND and_dcpl_83);
  COMP_LOOP_or_30_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_28_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_27_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_26_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_25_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_24_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_23_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_22_itm AND and_dcpl_83);
  COMP_LOOP_or_31_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm AND and_dcpl_49)
      OR (COMP_LOOP_COMP_LOOP_and_29_itm AND and_dcpl_54) OR (COMP_LOOP_COMP_LOOP_and_28_itm
      AND and_dcpl_58) OR (COMP_LOOP_COMP_LOOP_and_27_itm AND and_dcpl_65) OR (COMP_LOOP_COMP_LOOP_and_26_itm
      AND and_dcpl_68) OR (COMP_LOOP_COMP_LOOP_and_25_itm AND and_dcpl_75) OR (COMP_LOOP_COMP_LOOP_and_24_itm
      AND and_dcpl_78) OR (COMP_LOOP_COMP_LOOP_and_23_itm AND and_dcpl_83);
  COMP_LOOP_tmp_and_127_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(0)) AND COMP_LOOP_tmp_nor_49_itm
      AND (NOT and_294_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(1)) AND COMP_LOOP_tmp_nor_1_itm
      AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_128_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_129_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_130_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_131_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_132_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_133_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_134_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_135_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_136_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_137_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_138_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_139_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_140_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(4)) AND
      COMP_LOOP_tmp_nor_14_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_141_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_142_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_143_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_144_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_145_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_146_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_147_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_148_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_149_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_150_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_151_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_152_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_153_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_154_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_155_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm AND (NOT and_294_tmp);
  COMP_LOOP_tmp_and_115_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_3_0(0))
      AND COMP_LOOP_tmp_nor_25_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_3_0(1))
      AND COMP_LOOP_tmp_nor_26_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_116_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_3_0(2))
      AND COMP_LOOP_tmp_nor_28_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_117_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_118_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_119_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_3_0(3))
      AND COMP_LOOP_tmp_nor_31_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_120_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_121_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_122_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_123_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_124_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_125_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_126_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm AND (NOT nor_1119_tmp);
  COMP_LOOP_tmp_and_83_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_84_nl <= and_1_cse AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_85_nl <= and_4_cse AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_86_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_87_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_88_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_89_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_90_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_91_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_92_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_93_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_94_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_95_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_96_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_97_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_98_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_99_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_165 AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_100_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_101_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_102_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_103_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_104_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_105_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_106_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_107_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_108_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_109_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_110_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_111_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_112_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_113_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_114_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm AND (NOT nor_tmp);
  COMP_LOOP_tmp_and_78_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm AND (NOT nor_1117_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_nl <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("001")) AND (NOT nor_1117_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_nl <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("010")) AND (NOT nor_1117_tmp);
  COMP_LOOP_tmp_and_79_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_itm AND (NOT nor_1117_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_nl <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("100")) AND (NOT nor_1117_tmp);
  COMP_LOOP_tmp_and_80_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_itm AND (NOT nor_1117_tmp);
  COMP_LOOP_tmp_and_81_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_itm AND (NOT nor_1117_tmp);
  COMP_LOOP_tmp_and_82_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_itm AND (NOT nor_1117_tmp);
  COMP_LOOP_tmp_and_47_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_48_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_rgt AND and_298_m1c;
  COMP_LOOP_tmp_and_49_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_50_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_rgt AND and_298_m1c;
  COMP_LOOP_tmp_and_51_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_52_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_53_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_54_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_rgt AND and_298_m1c;
  COMP_LOOP_tmp_and_55_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_56_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_57_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_58_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_59_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_60_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_61_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_62_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_rgt AND and_298_m1c;
  COMP_LOOP_tmp_and_63_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_64_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_65_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_66_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_67_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_68_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_69_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_70_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_71_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_72_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_73_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_74_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_75_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_76_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm AND and_298_m1c;
  COMP_LOOP_tmp_and_77_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm AND and_298_m1c;
  nor_337_nl <= NOT(((fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(1))) OR
      CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  mux_1583_nl <= MUX_s_1_2_2(nor_337_nl, and_449_cse, fsm_output(4));
  mux_1582_nl <= MUX_s_1_2_2((NOT or_tmp_2075), and_464_cse, fsm_output(4));
  mux_1584_nl <= MUX_s_1_2_2(mux_1583_nl, mux_1582_nl, fsm_output(2));
  mux_1585_nl <= MUX_s_1_2_2(mux_1584_nl, and_464_cse, fsm_output(5));
  COMP_LOOP_tmp_and_15_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_16_nl <= and_1_cse AND mux_1592_tmp;
  COMP_LOOP_tmp_and_17_nl <= and_4_cse AND mux_1592_tmp;
  COMP_LOOP_tmp_and_18_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_19_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_169 AND mux_1592_tmp;
  COMP_LOOP_tmp_and_20_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_21_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_22_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_23_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_167 AND mux_1592_tmp;
  COMP_LOOP_tmp_and_24_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_25_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_26_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_27_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_28_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_29_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_30_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_31_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_165 AND mux_1592_tmp;
  COMP_LOOP_tmp_and_32_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_33_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_34_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_35_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_36_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_37_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_38_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_39_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_40_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_111_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_41_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_112_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_42_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_113_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_43_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_114_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_44_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_115_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_45_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_46_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_117_itm AND mux_1592_tmp;
  COMP_LOOP_tmp_and_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_1_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_119_rgt AND and_dcpl_177;
  COMP_LOOP_tmp_and_2_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_3_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_121_rgt AND and_dcpl_177;
  COMP_LOOP_tmp_and_4_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_122_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_5_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_123_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_6_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_124_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_7_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_125_rgt AND and_dcpl_177;
  COMP_LOOP_tmp_and_8_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_126_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_9_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_127_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_10_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_128_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_11_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_129_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_12_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_130_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_13_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_131_itm AND and_dcpl_177;
  COMP_LOOP_tmp_and_14_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_itm AND and_dcpl_177;
  mux_1594_nl <= MUX_s_1_2_2(mux_189_cse, and_464_cse, and_496_cse);
  mux_1595_nl <= MUX_s_1_2_2(mux_1594_nl, and_464_cse, fsm_output(4));
  mux_217_nl <= MUX_s_1_2_2(mux_189_cse, and_464_cse, or_212_cse);
  mux_1596_nl <= MUX_s_1_2_2(mux_1595_nl, mux_217_nl, fsm_output(2));
  and_478_nl <= (and_479_cse OR (fsm_output(6))) AND (fsm_output(7));
  mux_1597_nl <= MUX_s_1_2_2(mux_1596_nl, and_478_nl, fsm_output(5));
  and_755_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11")) AND and_dcpl_31
      AND and_dcpl_29 AND (fsm_output(2)) AND (fsm_output(5));
  COMP_LOOP_mux_382_nl <= MUX_v_7_2_2(COMP_LOOP_k_10_3_sva_6_0, (STD_LOGIC_VECTOR'(
      "001") & (NOT z_out_4)), and_755_nl);
  z_out_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_382_nl),
      8) + UNSIGNED'( "00000001"), 8));
  COMP_LOOP_mux_383_nl <= MUX_v_11_2_2(('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))), STAGE_LOOP_lshift_psp_sva, and_dcpl_334);
  COMP_LOOP_COMP_LOOP_nand_1_nl <= NOT(and_dcpl_334 AND (NOT(nor_1025_cse AND CONV_SL_1_1(fsm_output(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("10")) AND and_dcpl_29 AND and_dcpl_28)));
  COMP_LOOP_mux_384_nl <= MUX_v_10_2_2((COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'(
      "001")), VEC_LOOP_j_10_0_sva_9_0, and_dcpl_334);
  acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_383_nl & COMP_LOOP_COMP_LOOP_nand_1_nl)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_384_nl & '1'), 11), 12),
      12));
  z_out_3 <= acc_1_nl(11 DOWNTO 1);
  STAGE_LOOP_mux_4_nl <= MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, (NOT STAGE_LOOP_i_3_0_sva),
      and_dcpl_347);
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_mux_4_nl) + UNSIGNED('1'
      & (NOT and_dcpl_347) & STD_LOGIC_VECTOR'( "11")), 4));
  COMP_LOOP_mux_385_cse <= MUX_v_64_2_2(z_out_9, COMP_LOOP_1_acc_8_itm, COMP_LOOP_or_33_itm);
  COMP_LOOP_tmp_nor_135_cse <= NOT(and_dcpl_420 OR and_dcpl_435 OR and_dcpl_436);
  COMP_LOOP_tmp_mux_21_nl <= MUX_s_1_2_2((z_out_1(9)), (COMP_LOOP_2_tmp_lshift_ncse_sva(9)),
      COMP_LOOP_tmp_or_54_ssc);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_nl <= COMP_LOOP_tmp_mux_21_nl AND COMP_LOOP_tmp_nor_135_cse;
  COMP_LOOP_tmp_or_76_nl <= and_dcpl_423 OR and_dcpl_435;
  COMP_LOOP_tmp_mux1h_94_nl <= MUX1HOT_v_9_4_2(('0' & (z_out(7 DOWNTO 0))), (z_out_1(8
      DOWNTO 0)), (COMP_LOOP_2_tmp_lshift_ncse_sva(8 DOWNTO 0)), COMP_LOOP_3_tmp_lshift_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_420 & COMP_LOOP_tmp_or_76_nl & COMP_LOOP_tmp_or_54_ssc
      & and_dcpl_436));
  COMP_LOOP_tmp_and_161_nl <= (COMP_LOOP_k_10_3_sva_6_0(6)) AND COMP_LOOP_tmp_nor_135_cse;
  COMP_LOOP_tmp_or_77_nl <= and_dcpl_423 OR and_dcpl_428 OR and_dcpl_429 OR and_dcpl_434;
  COMP_LOOP_tmp_mux1h_95_nl <= MUX1HOT_v_6_3_2(('0' & (COMP_LOOP_k_10_3_sva_6_0(6
      DOWNTO 2))), (COMP_LOOP_k_10_3_sva_6_0(5 DOWNTO 0)), (COMP_LOOP_k_10_3_sva_6_0(6
      DOWNTO 1)), STD_LOGIC_VECTOR'( and_dcpl_420 & COMP_LOOP_tmp_or_77_nl & COMP_LOOP_tmp_or_71_itm));
  COMP_LOOP_tmp_COMP_LOOP_tmp_mux_18_nl <= MUX_s_1_2_2((COMP_LOOP_k_10_3_sva_6_0(1)),
      (COMP_LOOP_k_10_3_sva_6_0(0)), COMP_LOOP_tmp_or_71_itm);
  COMP_LOOP_tmp_or_78_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_mux_18_nl AND (NOT(and_dcpl_423
      OR and_dcpl_428))) OR and_dcpl_429 OR and_dcpl_434;
  COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl <= ((COMP_LOOP_k_10_3_sva_6_0(0)) AND (NOT(and_dcpl_423
      OR and_dcpl_429 OR and_dcpl_435))) OR and_dcpl_428 OR and_dcpl_434 OR and_dcpl_436;
  z_out_7 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_nl
      & COMP_LOOP_tmp_mux1h_94_nl) * UNSIGNED(COMP_LOOP_tmp_and_161_nl & COMP_LOOP_tmp_mux1h_95_nl
      & COMP_LOOP_tmp_or_78_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl & '1')), 10));
  and_756_nl <= nor_1025_cse AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND and_dcpl_30;
  COMP_LOOP_tmp_mux1h_96_nl <= MUX1HOT_v_64_9_2((STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000")
      & (z_out_1(6 DOWNTO 0))), COMP_LOOP_tmp_mux1h_itm, COMP_LOOP_tmp_mux1h_1_itm,
      COMP_LOOP_tmp_mux1h_2_itm, COMP_LOOP_tmp_mux1h_3_itm, COMP_LOOP_tmp_mux1h_4_itm,
      COMP_LOOP_tmp_mux1h_5_itm, COMP_LOOP_tmp_mux1h_6_itm, tmp_21_sva_1, STD_LOGIC_VECTOR'(
      and_756_nl & and_dcpl_448 & and_dcpl_452 & and_dcpl_456 & and_dcpl_458 & and_dcpl_461
      & and_dcpl_465 & and_dcpl_468 & and_dcpl_472));
  COMP_LOOP_tmp_or_79_nl <= and_dcpl_448 OR and_dcpl_452 OR and_dcpl_456 OR and_dcpl_458
      OR and_dcpl_461 OR and_dcpl_465 OR and_dcpl_468 OR and_dcpl_472;
  COMP_LOOP_tmp_mux_22_nl <= MUX_v_64_2_2((STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000")
      & COMP_LOOP_k_10_3_sva_6_0), COMP_LOOP_1_modulo_dev_cmp_return_rsc_z, COMP_LOOP_tmp_or_79_nl);
  z_out_8 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(COMP_LOOP_tmp_mux1h_96_nl)
      * UNSIGNED(COMP_LOOP_tmp_mux_22_nl)), 64));
  COMP_LOOP_mux1h_657_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_nor_itm, COMP_LOOP_COMP_LOOP_nor_5_itm,
      COMP_LOOP_COMP_LOOP_nor_9_itm, COMP_LOOP_COMP_LOOP_nor_13_itm, COMP_LOOP_COMP_LOOP_nor_17_itm,
      COMP_LOOP_COMP_LOOP_nor_21_itm, COMP_LOOP_COMP_LOOP_nor_25_itm, COMP_LOOP_COMP_LOOP_nor_29_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_COMP_LOOP_and_930_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(0)) AND COMP_LOOP_nor_126_itm;
  COMP_LOOP_COMP_LOOP_and_931_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(0)) AND COMP_LOOP_nor_226_itm;
  COMP_LOOP_COMP_LOOP_and_932_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(0)) AND COMP_LOOP_nor_326_itm;
  COMP_LOOP_COMP_LOOP_and_933_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) AND COMP_LOOP_nor_426_itm;
  COMP_LOOP_COMP_LOOP_and_934_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(0)) AND COMP_LOOP_nor_526_itm;
  COMP_LOOP_COMP_LOOP_and_935_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) AND COMP_LOOP_nor_626_itm;
  COMP_LOOP_COMP_LOOP_and_936_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(0)) AND COMP_LOOP_nor_726_itm;
  COMP_LOOP_mux1h_658_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_625_itm, COMP_LOOP_COMP_LOOP_and_930_nl,
      COMP_LOOP_COMP_LOOP_and_931_nl, COMP_LOOP_COMP_LOOP_and_932_nl, COMP_LOOP_COMP_LOOP_and_933_nl,
      COMP_LOOP_COMP_LOOP_and_934_nl, COMP_LOOP_COMP_LOOP_and_935_nl, COMP_LOOP_COMP_LOOP_and_936_nl,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_COMP_LOOP_and_937_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(1)) AND COMP_LOOP_nor_127_itm;
  COMP_LOOP_COMP_LOOP_and_938_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(1)) AND COMP_LOOP_nor_227_itm;
  COMP_LOOP_COMP_LOOP_and_939_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(1)) AND COMP_LOOP_nor_327_itm;
  COMP_LOOP_COMP_LOOP_and_940_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) AND COMP_LOOP_nor_427_itm;
  COMP_LOOP_COMP_LOOP_and_941_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(1)) AND COMP_LOOP_nor_527_itm;
  COMP_LOOP_COMP_LOOP_and_942_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) AND COMP_LOOP_nor_627_itm;
  COMP_LOOP_COMP_LOOP_and_943_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(1)) AND COMP_LOOP_nor_727_itm;
  COMP_LOOP_mux1h_659_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_126_itm, COMP_LOOP_COMP_LOOP_and_937_nl,
      COMP_LOOP_COMP_LOOP_and_938_nl, COMP_LOOP_COMP_LOOP_and_939_nl, COMP_LOOP_COMP_LOOP_and_940_nl,
      COMP_LOOP_COMP_LOOP_and_941_nl, COMP_LOOP_COMP_LOOP_and_942_nl, COMP_LOOP_COMP_LOOP_and_943_nl,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_660_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_377_itm, COMP_LOOP_COMP_LOOP_and_157_itm,
      COMP_LOOP_COMP_LOOP_and_281_itm, COMP_LOOP_COMP_LOOP_and_405_itm, COMP_LOOP_COMP_LOOP_and_529_itm,
      COMP_LOOP_COMP_LOOP_and_653_itm, COMP_LOOP_COMP_LOOP_and_777_itm, COMP_LOOP_COMP_LOOP_and_901_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_COMP_LOOP_and_944_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(2)) AND COMP_LOOP_nor_129_itm;
  COMP_LOOP_COMP_LOOP_and_945_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(2)) AND COMP_LOOP_nor_229_itm;
  COMP_LOOP_COMP_LOOP_and_946_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(2)) AND COMP_LOOP_nor_329_itm;
  COMP_LOOP_COMP_LOOP_and_947_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(2)) AND COMP_LOOP_nor_429_itm;
  COMP_LOOP_COMP_LOOP_and_948_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(2)) AND COMP_LOOP_nor_529_itm;
  COMP_LOOP_COMP_LOOP_and_949_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(2)) AND COMP_LOOP_nor_629_itm;
  COMP_LOOP_COMP_LOOP_and_950_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(2)) AND COMP_LOOP_nor_729_itm;
  COMP_LOOP_mux1h_661_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_128_itm, COMP_LOOP_COMP_LOOP_and_944_nl,
      COMP_LOOP_COMP_LOOP_and_945_nl, COMP_LOOP_COMP_LOOP_and_946_nl, COMP_LOOP_COMP_LOOP_and_947_nl,
      COMP_LOOP_COMP_LOOP_and_948_nl, COMP_LOOP_COMP_LOOP_and_949_nl, COMP_LOOP_COMP_LOOP_and_950_nl,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_662_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_129_itm, COMP_LOOP_COMP_LOOP_and_159_itm,
      COMP_LOOP_COMP_LOOP_and_283_itm, COMP_LOOP_COMP_LOOP_and_407_itm, COMP_LOOP_COMP_LOOP_and_531_itm,
      COMP_LOOP_COMP_LOOP_and_655_itm, COMP_LOOP_COMP_LOOP_and_779_itm, COMP_LOOP_COMP_LOOP_and_903_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_663_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_130_itm, COMP_LOOP_COMP_LOOP_and_160_itm,
      COMP_LOOP_COMP_LOOP_and_284_itm, COMP_LOOP_COMP_LOOP_and_408_itm, COMP_LOOP_COMP_LOOP_and_532_itm,
      COMP_LOOP_COMP_LOOP_and_656_itm, COMP_LOOP_COMP_LOOP_and_780_itm, COMP_LOOP_COMP_LOOP_and_904_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_664_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_6_itm, COMP_LOOP_COMP_LOOP_and_161_itm,
      COMP_LOOP_COMP_LOOP_and_285_itm, COMP_LOOP_COMP_LOOP_and_409_itm, COMP_LOOP_COMP_LOOP_and_533_itm,
      COMP_LOOP_COMP_LOOP_and_657_itm, COMP_LOOP_COMP_LOOP_and_781_itm, COMP_LOOP_COMP_LOOP_and_905_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_COMP_LOOP_and_951_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(3)) AND COMP_LOOP_nor_133_itm;
  COMP_LOOP_COMP_LOOP_and_952_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(3)) AND COMP_LOOP_nor_233_itm;
  COMP_LOOP_COMP_LOOP_and_953_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(3)) AND COMP_LOOP_nor_333_itm;
  COMP_LOOP_COMP_LOOP_and_954_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) AND COMP_LOOP_nor_433_itm;
  COMP_LOOP_COMP_LOOP_and_955_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(3)) AND COMP_LOOP_nor_533_itm;
  COMP_LOOP_COMP_LOOP_and_956_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(3)) AND COMP_LOOP_nor_633_itm;
  COMP_LOOP_COMP_LOOP_and_957_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(3)) AND COMP_LOOP_nor_733_itm;
  COMP_LOOP_mux1h_665_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_132_itm, COMP_LOOP_COMP_LOOP_and_951_nl,
      COMP_LOOP_COMP_LOOP_and_952_nl, COMP_LOOP_COMP_LOOP_and_953_nl, COMP_LOOP_COMP_LOOP_and_954_nl,
      COMP_LOOP_COMP_LOOP_and_955_nl, COMP_LOOP_COMP_LOOP_and_956_nl, COMP_LOOP_COMP_LOOP_and_957_nl,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_666_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_133_itm, COMP_LOOP_COMP_LOOP_and_163_itm,
      COMP_LOOP_COMP_LOOP_and_287_itm, COMP_LOOP_COMP_LOOP_and_411_itm, COMP_LOOP_COMP_LOOP_and_535_itm,
      COMP_LOOP_COMP_LOOP_and_659_itm, COMP_LOOP_COMP_LOOP_and_783_itm, COMP_LOOP_COMP_LOOP_and_907_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_667_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_134_itm, COMP_LOOP_COMP_LOOP_and_164_itm,
      COMP_LOOP_COMP_LOOP_and_288_itm, COMP_LOOP_COMP_LOOP_and_412_itm, COMP_LOOP_COMP_LOOP_and_536_itm,
      COMP_LOOP_COMP_LOOP_and_660_itm, COMP_LOOP_COMP_LOOP_and_784_itm, COMP_LOOP_COMP_LOOP_and_908_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_668_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_10_itm, COMP_LOOP_COMP_LOOP_and_165_itm,
      COMP_LOOP_COMP_LOOP_and_289_itm, COMP_LOOP_COMP_LOOP_and_413_itm, COMP_LOOP_COMP_LOOP_and_537_itm,
      COMP_LOOP_COMP_LOOP_and_661_itm, COMP_LOOP_COMP_LOOP_and_785_itm, COMP_LOOP_COMP_LOOP_and_909_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_669_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_136_itm, COMP_LOOP_COMP_LOOP_and_166_itm,
      COMP_LOOP_COMP_LOOP_and_290_itm, COMP_LOOP_COMP_LOOP_and_414_itm, COMP_LOOP_COMP_LOOP_and_538_itm,
      COMP_LOOP_COMP_LOOP_and_662_itm, COMP_LOOP_COMP_LOOP_and_786_itm, COMP_LOOP_COMP_LOOP_and_910_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_670_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_12_itm, COMP_LOOP_COMP_LOOP_and_167_itm,
      COMP_LOOP_COMP_LOOP_and_291_itm, COMP_LOOP_COMP_LOOP_and_415_itm, COMP_LOOP_COMP_LOOP_and_539_itm,
      COMP_LOOP_COMP_LOOP_and_663_itm, COMP_LOOP_COMP_LOOP_and_787_itm, COMP_LOOP_COMP_LOOP_and_911_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_671_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_13_itm, COMP_LOOP_COMP_LOOP_and_168_itm,
      COMP_LOOP_COMP_LOOP_and_292_itm, COMP_LOOP_COMP_LOOP_and_416_itm, COMP_LOOP_COMP_LOOP_and_540_itm,
      COMP_LOOP_COMP_LOOP_and_664_itm, COMP_LOOP_COMP_LOOP_and_788_itm, COMP_LOOP_COMP_LOOP_and_912_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_672_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_14_itm, COMP_LOOP_COMP_LOOP_and_169_itm,
      COMP_LOOP_COMP_LOOP_and_293_itm, COMP_LOOP_COMP_LOOP_and_417_itm, COMP_LOOP_COMP_LOOP_and_541_itm,
      COMP_LOOP_COMP_LOOP_and_665_itm, COMP_LOOP_COMP_LOOP_and_789_itm, COMP_LOOP_COMP_LOOP_and_913_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_COMP_LOOP_and_958_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(4)) AND COMP_LOOP_nor_140_itm;
  COMP_LOOP_COMP_LOOP_and_959_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(4)) AND COMP_LOOP_nor_240_itm;
  COMP_LOOP_COMP_LOOP_and_960_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(4)) AND COMP_LOOP_nor_340_itm;
  COMP_LOOP_COMP_LOOP_and_961_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(4)) AND COMP_LOOP_nor_440_itm;
  COMP_LOOP_COMP_LOOP_and_962_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(4)) AND COMP_LOOP_nor_540_itm;
  COMP_LOOP_COMP_LOOP_and_963_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(4)) AND COMP_LOOP_nor_640_itm;
  COMP_LOOP_COMP_LOOP_and_964_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(4)) AND COMP_LOOP_nor_740_itm;
  COMP_LOOP_mux1h_673_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_140_itm, COMP_LOOP_COMP_LOOP_and_958_nl,
      COMP_LOOP_COMP_LOOP_and_959_nl, COMP_LOOP_COMP_LOOP_and_960_nl, COMP_LOOP_COMP_LOOP_and_961_nl,
      COMP_LOOP_COMP_LOOP_and_962_nl, COMP_LOOP_COMP_LOOP_and_963_nl, COMP_LOOP_COMP_LOOP_and_964_nl,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_674_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_141_itm, COMP_LOOP_COMP_LOOP_and_171_itm,
      COMP_LOOP_COMP_LOOP_and_295_itm, COMP_LOOP_COMP_LOOP_and_419_itm, COMP_LOOP_COMP_LOOP_and_543_itm,
      COMP_LOOP_COMP_LOOP_and_667_itm, COMP_LOOP_COMP_LOOP_and_791_itm, COMP_LOOP_COMP_LOOP_and_915_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_675_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_142_itm, COMP_LOOP_COMP_LOOP_and_172_itm,
      COMP_LOOP_COMP_LOOP_and_296_itm, COMP_LOOP_COMP_LOOP_and_420_itm, COMP_LOOP_COMP_LOOP_and_544_itm,
      COMP_LOOP_COMP_LOOP_and_668_itm, COMP_LOOP_COMP_LOOP_and_792_itm, COMP_LOOP_COMP_LOOP_and_916_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_676_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_18_itm, COMP_LOOP_COMP_LOOP_and_173_itm,
      COMP_LOOP_COMP_LOOP_and_297_itm, COMP_LOOP_COMP_LOOP_and_421_itm, COMP_LOOP_COMP_LOOP_and_545_itm,
      COMP_LOOP_COMP_LOOP_and_669_itm, COMP_LOOP_COMP_LOOP_and_793_itm, COMP_LOOP_COMP_LOOP_and_917_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_677_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_144_itm, COMP_LOOP_COMP_LOOP_and_174_itm,
      COMP_LOOP_COMP_LOOP_and_298_itm, COMP_LOOP_COMP_LOOP_and_422_itm, COMP_LOOP_COMP_LOOP_and_546_itm,
      COMP_LOOP_COMP_LOOP_and_670_itm, COMP_LOOP_COMP_LOOP_and_794_itm, COMP_LOOP_COMP_LOOP_and_918_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_678_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_20_itm, COMP_LOOP_COMP_LOOP_and_175_itm,
      COMP_LOOP_COMP_LOOP_and_299_itm, COMP_LOOP_COMP_LOOP_and_423_itm, COMP_LOOP_COMP_LOOP_and_547_itm,
      COMP_LOOP_COMP_LOOP_and_671_itm, COMP_LOOP_COMP_LOOP_and_795_itm, COMP_LOOP_COMP_LOOP_and_919_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_679_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_21_itm, COMP_LOOP_COMP_LOOP_and_176_itm,
      COMP_LOOP_COMP_LOOP_and_300_itm, COMP_LOOP_COMP_LOOP_and_424_itm, COMP_LOOP_COMP_LOOP_and_548_itm,
      COMP_LOOP_COMP_LOOP_and_672_itm, COMP_LOOP_COMP_LOOP_and_796_itm, COMP_LOOP_COMP_LOOP_and_920_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_680_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_22_itm, COMP_LOOP_COMP_LOOP_and_177_itm,
      COMP_LOOP_COMP_LOOP_and_301_itm, COMP_LOOP_COMP_LOOP_and_425_itm, COMP_LOOP_COMP_LOOP_and_549_itm,
      COMP_LOOP_COMP_LOOP_and_673_itm, COMP_LOOP_COMP_LOOP_and_797_itm, COMP_LOOP_COMP_LOOP_and_921_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_681_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_23_itm, COMP_LOOP_COMP_LOOP_and_178_itm,
      COMP_LOOP_COMP_LOOP_and_302_itm, COMP_LOOP_COMP_LOOP_and_426_itm, COMP_LOOP_COMP_LOOP_and_550_itm,
      COMP_LOOP_COMP_LOOP_and_674_itm, COMP_LOOP_COMP_LOOP_and_798_itm, COMP_LOOP_COMP_LOOP_and_922_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_682_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_24_itm, COMP_LOOP_COMP_LOOP_and_179_itm,
      COMP_LOOP_COMP_LOOP_and_303_itm, COMP_LOOP_COMP_LOOP_and_427_itm, COMP_LOOP_COMP_LOOP_and_551_itm,
      COMP_LOOP_COMP_LOOP_and_675_itm, COMP_LOOP_COMP_LOOP_and_799_itm, COMP_LOOP_COMP_LOOP_and_923_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_683_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_25_itm, COMP_LOOP_COMP_LOOP_and_180_itm,
      COMP_LOOP_COMP_LOOP_and_304_itm, COMP_LOOP_COMP_LOOP_and_428_itm, COMP_LOOP_COMP_LOOP_and_552_itm,
      COMP_LOOP_COMP_LOOP_and_676_itm, COMP_LOOP_COMP_LOOP_and_800_itm, COMP_LOOP_COMP_LOOP_and_924_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_684_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_26_itm, COMP_LOOP_COMP_LOOP_and_181_itm,
      COMP_LOOP_COMP_LOOP_and_305_itm, COMP_LOOP_COMP_LOOP_and_429_itm, COMP_LOOP_COMP_LOOP_and_553_itm,
      COMP_LOOP_COMP_LOOP_and_677_itm, COMP_LOOP_COMP_LOOP_and_801_itm, COMP_LOOP_COMP_LOOP_and_925_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_685_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_27_itm, COMP_LOOP_COMP_LOOP_and_182_itm,
      COMP_LOOP_COMP_LOOP_and_306_itm, COMP_LOOP_COMP_LOOP_and_430_itm, COMP_LOOP_COMP_LOOP_and_554_itm,
      COMP_LOOP_COMP_LOOP_and_678_itm, COMP_LOOP_COMP_LOOP_and_802_itm, COMP_LOOP_COMP_LOOP_and_926_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_686_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_28_itm, COMP_LOOP_COMP_LOOP_and_183_itm,
      COMP_LOOP_COMP_LOOP_and_307_itm, COMP_LOOP_COMP_LOOP_and_431_itm, COMP_LOOP_COMP_LOOP_and_555_itm,
      COMP_LOOP_COMP_LOOP_and_679_itm, COMP_LOOP_COMP_LOOP_and_803_itm, COMP_LOOP_COMP_LOOP_and_927_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_687_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_29_itm, COMP_LOOP_COMP_LOOP_and_184_itm,
      COMP_LOOP_COMP_LOOP_and_308_itm, COMP_LOOP_COMP_LOOP_and_432_itm, COMP_LOOP_COMP_LOOP_and_556_itm,
      COMP_LOOP_COMP_LOOP_and_680_itm, COMP_LOOP_COMP_LOOP_and_804_itm, COMP_LOOP_COMP_LOOP_and_928_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  COMP_LOOP_mux1h_688_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_30_itm, COMP_LOOP_COMP_LOOP_and_185_itm,
      COMP_LOOP_COMP_LOOP_and_309_itm, COMP_LOOP_COMP_LOOP_and_433_itm, COMP_LOOP_COMP_LOOP_and_557_itm,
      COMP_LOOP_COMP_LOOP_and_681_itm, COMP_LOOP_COMP_LOOP_and_805_itm, COMP_LOOP_COMP_LOOP_and_929_itm,
      STD_LOGIC_VECTOR'( and_dcpl_479 & and_605_cse & and_609_cse & and_614_cse &
      and_617_cse & and_621_cse & and_624_cse & and_628_cse));
  z_out_9 <= MUX1HOT_v_64_32_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d, vec_rsc_0_2_i_q_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d, vec_rsc_0_6_i_q_d,
      vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d, vec_rsc_0_14_i_q_d,
      vec_rsc_0_15_i_q_d, vec_rsc_0_16_i_q_d, vec_rsc_0_17_i_q_d, vec_rsc_0_18_i_q_d,
      vec_rsc_0_19_i_q_d, vec_rsc_0_20_i_q_d, vec_rsc_0_21_i_q_d, vec_rsc_0_22_i_q_d,
      vec_rsc_0_23_i_q_d, vec_rsc_0_24_i_q_d, vec_rsc_0_25_i_q_d, vec_rsc_0_26_i_q_d,
      vec_rsc_0_27_i_q_d, vec_rsc_0_28_i_q_d, vec_rsc_0_29_i_q_d, vec_rsc_0_30_i_q_d,
      vec_rsc_0_31_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_mux1h_657_nl & COMP_LOOP_mux1h_658_nl
      & COMP_LOOP_mux1h_659_nl & COMP_LOOP_mux1h_660_nl & COMP_LOOP_mux1h_661_nl
      & COMP_LOOP_mux1h_662_nl & COMP_LOOP_mux1h_663_nl & COMP_LOOP_mux1h_664_nl
      & COMP_LOOP_mux1h_665_nl & COMP_LOOP_mux1h_666_nl & COMP_LOOP_mux1h_667_nl
      & COMP_LOOP_mux1h_668_nl & COMP_LOOP_mux1h_669_nl & COMP_LOOP_mux1h_670_nl
      & COMP_LOOP_mux1h_671_nl & COMP_LOOP_mux1h_672_nl & COMP_LOOP_mux1h_673_nl
      & COMP_LOOP_mux1h_674_nl & COMP_LOOP_mux1h_675_nl & COMP_LOOP_mux1h_676_nl
      & COMP_LOOP_mux1h_677_nl & COMP_LOOP_mux1h_678_nl & COMP_LOOP_mux1h_679_nl
      & COMP_LOOP_mux1h_680_nl & COMP_LOOP_mux1h_681_nl & COMP_LOOP_mux1h_682_nl
      & COMP_LOOP_mux1h_683_nl & COMP_LOOP_mux1h_684_nl & COMP_LOOP_mux1h_685_nl
      & COMP_LOOP_mux1h_686_nl & COMP_LOOP_mux1h_687_nl & COMP_LOOP_mux1h_688_nl));
END v13;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_0_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_we : OUT STD_LOGIC;
    vec_rsc_0_0_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_0_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_1_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_we : OUT STD_LOGIC;
    vec_rsc_0_1_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_1_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_2_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_we : OUT STD_LOGIC;
    vec_rsc_0_2_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_2_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_3_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_we : OUT STD_LOGIC;
    vec_rsc_0_3_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_3_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_4_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_we : OUT STD_LOGIC;
    vec_rsc_0_4_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_4_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_5_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_we : OUT STD_LOGIC;
    vec_rsc_0_5_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_5_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_6_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_we : OUT STD_LOGIC;
    vec_rsc_0_6_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_6_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_7_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_we : OUT STD_LOGIC;
    vec_rsc_0_7_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_7_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_0_8_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_8_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_we : OUT STD_LOGIC;
    vec_rsc_0_8_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_8_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_0_9_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_9_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_we : OUT STD_LOGIC;
    vec_rsc_0_9_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_9_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_0_10_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_10_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_we : OUT STD_LOGIC;
    vec_rsc_0_10_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_10_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_0_11_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_11_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_we : OUT STD_LOGIC;
    vec_rsc_0_11_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_11_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_0_12_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_12_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_we : OUT STD_LOGIC;
    vec_rsc_0_12_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_12_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_0_13_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_13_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_we : OUT STD_LOGIC;
    vec_rsc_0_13_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_13_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_0_14_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_14_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_we : OUT STD_LOGIC;
    vec_rsc_0_14_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_14_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_0_15_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_15_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_we : OUT STD_LOGIC;
    vec_rsc_0_15_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_15_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    vec_rsc_0_16_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_16_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_16_we : OUT STD_LOGIC;
    vec_rsc_0_16_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_16_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    vec_rsc_0_17_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_17_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_17_we : OUT STD_LOGIC;
    vec_rsc_0_17_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_17_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    vec_rsc_0_18_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_18_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_18_we : OUT STD_LOGIC;
    vec_rsc_0_18_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_18_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    vec_rsc_0_19_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_19_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_19_we : OUT STD_LOGIC;
    vec_rsc_0_19_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_19_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    vec_rsc_0_20_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_20_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_20_we : OUT STD_LOGIC;
    vec_rsc_0_20_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_20_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    vec_rsc_0_21_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_21_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_21_we : OUT STD_LOGIC;
    vec_rsc_0_21_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_21_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    vec_rsc_0_22_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_22_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_22_we : OUT STD_LOGIC;
    vec_rsc_0_22_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_22_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    vec_rsc_0_23_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_23_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_23_we : OUT STD_LOGIC;
    vec_rsc_0_23_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_23_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    vec_rsc_0_24_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_24_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_24_we : OUT STD_LOGIC;
    vec_rsc_0_24_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_24_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    vec_rsc_0_25_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_25_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_25_we : OUT STD_LOGIC;
    vec_rsc_0_25_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_25_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    vec_rsc_0_26_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_26_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_26_we : OUT STD_LOGIC;
    vec_rsc_0_26_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_26_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    vec_rsc_0_27_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_27_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_27_we : OUT STD_LOGIC;
    vec_rsc_0_27_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_27_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    vec_rsc_0_28_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_28_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_28_we : OUT STD_LOGIC;
    vec_rsc_0_28_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_28_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    vec_rsc_0_29_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_29_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_29_we : OUT STD_LOGIC;
    vec_rsc_0_29_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_29_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    vec_rsc_0_30_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_30_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_30_we : OUT STD_LOGIC;
    vec_rsc_0_30_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_30_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    vec_rsc_0_31_wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_31_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_31_we : OUT STD_LOGIC;
    vec_rsc_0_31_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    vec_rsc_0_31_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_0_0_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_0_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_0_1_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_1_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_0_2_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_2_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_0_3_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_3_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_0_4_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_4_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_0_5_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_5_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_0_6_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_6_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_0_7_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_7_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_0_8_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_8_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_0_9_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_9_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_0_10_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_10_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_0_11_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_11_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_0_12_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_12_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_0_13_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_13_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_0_14_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_14_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_0_15_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_15_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_rsc_0_16_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_16_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    twiddle_rsc_0_17_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_17_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    twiddle_rsc_0_18_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_18_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    twiddle_rsc_0_19_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_19_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    twiddle_rsc_0_20_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_20_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    twiddle_rsc_0_21_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_21_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    twiddle_rsc_0_22_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_22_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    twiddle_rsc_0_23_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_23_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    twiddle_rsc_0_24_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_24_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    twiddle_rsc_0_25_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_25_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    twiddle_rsc_0_26_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_26_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    twiddle_rsc_0_27_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_27_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    twiddle_rsc_0_28_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_28_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    twiddle_rsc_0_29_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_29_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    twiddle_rsc_0_30_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_30_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    twiddle_rsc_0_31_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_0_31_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_31_lz : OUT STD_LOGIC
  );
END inPlaceNTT_DIF;

ARCHITECTURE v13 OF inPlaceNTT_DIF IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_d_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr_d_iff : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr_d_iff : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_16_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_17_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_18_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_19_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_20_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_21_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_22_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_23_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_24_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_25_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_26_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_27_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_28_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_29_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_30_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_31_i_we_d_iff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_radr_d_iff : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_radr_d_iff : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr_d_iff : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr_d_iff : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_8_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_9_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_10_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_11_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_12_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_13_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_14_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_15_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_16_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_17_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_18_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_19_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_20_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_21_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_22_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_23_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_24_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_25_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_26_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_27_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_28_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_29_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_30_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_31_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_wadr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_wadr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_0_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_1_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_2_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_3_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_4_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_5_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_6_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_7_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_8_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_9_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_10_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_11_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_12_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_13_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_14_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_15_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_16_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_16_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_16_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_16_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_17_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_17_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_17_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_17_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_18_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_18_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_18_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_18_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_19_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_19_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_19_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_19_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_20_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_20_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_20_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_20_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_21_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_21_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_21_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_21_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_22_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_22_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_22_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_22_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_23_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_23_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_23_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_23_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_24_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_24_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_24_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_24_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_25_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_25_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_25_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_25_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_26_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_26_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_26_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_26_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_27_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_27_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_27_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_27_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_28_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_28_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_28_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_28_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_29_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_29_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_29_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_29_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_30_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_30_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_30_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_30_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_31_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_31_i_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsc_0_31_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_31_i_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_16_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_17_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_18_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_19_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_20_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_21_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_22_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_23_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_24_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_25_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_26_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_27_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_28_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_29_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_30_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_31_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_16_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_17_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_18_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_19_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_20_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_21_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_22_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_23_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_24_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_25_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_26_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_27_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_28_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_29_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_30_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_31_lz : OUT STD_LOGIC;
      vec_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      vec_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      vec_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_1_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_2_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_3_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_4_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_5_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_6_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_7_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_8_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_9_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_10_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_11_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_12_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_13_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_14_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_15_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_16_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_17_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_18_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_19_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_20_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_21_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_22_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_23_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_24_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_25_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_26_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_27_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_28_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_29_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_30_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_31_i_we_d_pff : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_rsc_0_1_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_rsc_0_2_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_rsc_0_4_i_radr_d_pff : OUT STD_LOGIC_VECTOR (4 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff : STD_LOGIC_VECTOR (4
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff : STD_LOGIC_VECTOR (4
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d_pff : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff : STD_LOGIC_VECTOR
      (4 DOWNTO 0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_0_i_q,
      radr => vec_rsc_0_0_i_radr,
      we => vec_rsc_0_0_we,
      d => vec_rsc_0_0_i_d,
      wadr => vec_rsc_0_0_i_wadr,
      d_d => vec_rsc_0_0_i_d_d,
      q_d => vec_rsc_0_0_i_q_d_1,
      radr_d => vec_rsc_0_0_i_radr_d,
      wadr_d => vec_rsc_0_0_i_wadr_d,
      we_d => vec_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_0_i_q <= vec_rsc_0_0_q;
  vec_rsc_0_0_radr <= vec_rsc_0_0_i_radr;
  vec_rsc_0_0_d <= vec_rsc_0_0_i_d;
  vec_rsc_0_0_wadr <= vec_rsc_0_0_i_wadr;
  vec_rsc_0_0_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_0_i_q_d <= vec_rsc_0_0_i_q_d_1;
  vec_rsc_0_0_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_0_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_1_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_1_i_q,
      radr => vec_rsc_0_1_i_radr,
      we => vec_rsc_0_1_we,
      d => vec_rsc_0_1_i_d,
      wadr => vec_rsc_0_1_i_wadr,
      d_d => vec_rsc_0_1_i_d_d,
      q_d => vec_rsc_0_1_i_q_d_1,
      radr_d => vec_rsc_0_1_i_radr_d,
      wadr_d => vec_rsc_0_1_i_wadr_d,
      we_d => vec_rsc_0_1_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_1_i_q <= vec_rsc_0_1_q;
  vec_rsc_0_1_radr <= vec_rsc_0_1_i_radr;
  vec_rsc_0_1_d <= vec_rsc_0_1_i_d;
  vec_rsc_0_1_wadr <= vec_rsc_0_1_i_wadr;
  vec_rsc_0_1_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_1_i_q_d <= vec_rsc_0_1_i_q_d_1;
  vec_rsc_0_1_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_1_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_2_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_2_i_q,
      radr => vec_rsc_0_2_i_radr,
      we => vec_rsc_0_2_we,
      d => vec_rsc_0_2_i_d,
      wadr => vec_rsc_0_2_i_wadr,
      d_d => vec_rsc_0_2_i_d_d,
      q_d => vec_rsc_0_2_i_q_d_1,
      radr_d => vec_rsc_0_2_i_radr_d,
      wadr_d => vec_rsc_0_2_i_wadr_d,
      we_d => vec_rsc_0_2_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_2_i_q <= vec_rsc_0_2_q;
  vec_rsc_0_2_radr <= vec_rsc_0_2_i_radr;
  vec_rsc_0_2_d <= vec_rsc_0_2_i_d;
  vec_rsc_0_2_wadr <= vec_rsc_0_2_i_wadr;
  vec_rsc_0_2_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_2_i_q_d <= vec_rsc_0_2_i_q_d_1;
  vec_rsc_0_2_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_2_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_3_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_3_i_q,
      radr => vec_rsc_0_3_i_radr,
      we => vec_rsc_0_3_we,
      d => vec_rsc_0_3_i_d,
      wadr => vec_rsc_0_3_i_wadr,
      d_d => vec_rsc_0_3_i_d_d,
      q_d => vec_rsc_0_3_i_q_d_1,
      radr_d => vec_rsc_0_3_i_radr_d,
      wadr_d => vec_rsc_0_3_i_wadr_d,
      we_d => vec_rsc_0_3_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_3_i_q <= vec_rsc_0_3_q;
  vec_rsc_0_3_radr <= vec_rsc_0_3_i_radr;
  vec_rsc_0_3_d <= vec_rsc_0_3_i_d;
  vec_rsc_0_3_wadr <= vec_rsc_0_3_i_wadr;
  vec_rsc_0_3_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_3_i_q_d <= vec_rsc_0_3_i_q_d_1;
  vec_rsc_0_3_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_3_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_4_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_4_i_q,
      radr => vec_rsc_0_4_i_radr,
      we => vec_rsc_0_4_we,
      d => vec_rsc_0_4_i_d,
      wadr => vec_rsc_0_4_i_wadr,
      d_d => vec_rsc_0_4_i_d_d,
      q_d => vec_rsc_0_4_i_q_d_1,
      radr_d => vec_rsc_0_4_i_radr_d,
      wadr_d => vec_rsc_0_4_i_wadr_d,
      we_d => vec_rsc_0_4_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_4_i_q <= vec_rsc_0_4_q;
  vec_rsc_0_4_radr <= vec_rsc_0_4_i_radr;
  vec_rsc_0_4_d <= vec_rsc_0_4_i_d;
  vec_rsc_0_4_wadr <= vec_rsc_0_4_i_wadr;
  vec_rsc_0_4_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_4_i_q_d <= vec_rsc_0_4_i_q_d_1;
  vec_rsc_0_4_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_4_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_5_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_5_i_q,
      radr => vec_rsc_0_5_i_radr,
      we => vec_rsc_0_5_we,
      d => vec_rsc_0_5_i_d,
      wadr => vec_rsc_0_5_i_wadr,
      d_d => vec_rsc_0_5_i_d_d,
      q_d => vec_rsc_0_5_i_q_d_1,
      radr_d => vec_rsc_0_5_i_radr_d,
      wadr_d => vec_rsc_0_5_i_wadr_d,
      we_d => vec_rsc_0_5_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_5_i_q <= vec_rsc_0_5_q;
  vec_rsc_0_5_radr <= vec_rsc_0_5_i_radr;
  vec_rsc_0_5_d <= vec_rsc_0_5_i_d;
  vec_rsc_0_5_wadr <= vec_rsc_0_5_i_wadr;
  vec_rsc_0_5_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_5_i_q_d <= vec_rsc_0_5_i_q_d_1;
  vec_rsc_0_5_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_5_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_6_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_6_i_q,
      radr => vec_rsc_0_6_i_radr,
      we => vec_rsc_0_6_we,
      d => vec_rsc_0_6_i_d,
      wadr => vec_rsc_0_6_i_wadr,
      d_d => vec_rsc_0_6_i_d_d,
      q_d => vec_rsc_0_6_i_q_d_1,
      radr_d => vec_rsc_0_6_i_radr_d,
      wadr_d => vec_rsc_0_6_i_wadr_d,
      we_d => vec_rsc_0_6_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_6_i_q <= vec_rsc_0_6_q;
  vec_rsc_0_6_radr <= vec_rsc_0_6_i_radr;
  vec_rsc_0_6_d <= vec_rsc_0_6_i_d;
  vec_rsc_0_6_wadr <= vec_rsc_0_6_i_wadr;
  vec_rsc_0_6_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_6_i_q_d <= vec_rsc_0_6_i_q_d_1;
  vec_rsc_0_6_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_6_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_7_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_7_i_q,
      radr => vec_rsc_0_7_i_radr,
      we => vec_rsc_0_7_we,
      d => vec_rsc_0_7_i_d,
      wadr => vec_rsc_0_7_i_wadr,
      d_d => vec_rsc_0_7_i_d_d,
      q_d => vec_rsc_0_7_i_q_d_1,
      radr_d => vec_rsc_0_7_i_radr_d,
      wadr_d => vec_rsc_0_7_i_wadr_d,
      we_d => vec_rsc_0_7_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_7_i_q <= vec_rsc_0_7_q;
  vec_rsc_0_7_radr <= vec_rsc_0_7_i_radr;
  vec_rsc_0_7_d <= vec_rsc_0_7_i_d;
  vec_rsc_0_7_wadr <= vec_rsc_0_7_i_wadr;
  vec_rsc_0_7_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_7_i_q_d <= vec_rsc_0_7_i_q_d_1;
  vec_rsc_0_7_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_7_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_8_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_8_i_q,
      radr => vec_rsc_0_8_i_radr,
      we => vec_rsc_0_8_we,
      d => vec_rsc_0_8_i_d,
      wadr => vec_rsc_0_8_i_wadr,
      d_d => vec_rsc_0_8_i_d_d,
      q_d => vec_rsc_0_8_i_q_d_1,
      radr_d => vec_rsc_0_8_i_radr_d,
      wadr_d => vec_rsc_0_8_i_wadr_d,
      we_d => vec_rsc_0_8_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_8_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_8_i_q <= vec_rsc_0_8_q;
  vec_rsc_0_8_radr <= vec_rsc_0_8_i_radr;
  vec_rsc_0_8_d <= vec_rsc_0_8_i_d;
  vec_rsc_0_8_wadr <= vec_rsc_0_8_i_wadr;
  vec_rsc_0_8_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_8_i_q_d <= vec_rsc_0_8_i_q_d_1;
  vec_rsc_0_8_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_8_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_9_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_9_i_q,
      radr => vec_rsc_0_9_i_radr,
      we => vec_rsc_0_9_we,
      d => vec_rsc_0_9_i_d,
      wadr => vec_rsc_0_9_i_wadr,
      d_d => vec_rsc_0_9_i_d_d,
      q_d => vec_rsc_0_9_i_q_d_1,
      radr_d => vec_rsc_0_9_i_radr_d,
      wadr_d => vec_rsc_0_9_i_wadr_d,
      we_d => vec_rsc_0_9_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_9_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_9_i_q <= vec_rsc_0_9_q;
  vec_rsc_0_9_radr <= vec_rsc_0_9_i_radr;
  vec_rsc_0_9_d <= vec_rsc_0_9_i_d;
  vec_rsc_0_9_wadr <= vec_rsc_0_9_i_wadr;
  vec_rsc_0_9_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_9_i_q_d <= vec_rsc_0_9_i_q_d_1;
  vec_rsc_0_9_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_9_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_10_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_10_i_q,
      radr => vec_rsc_0_10_i_radr,
      we => vec_rsc_0_10_we,
      d => vec_rsc_0_10_i_d,
      wadr => vec_rsc_0_10_i_wadr,
      d_d => vec_rsc_0_10_i_d_d,
      q_d => vec_rsc_0_10_i_q_d_1,
      radr_d => vec_rsc_0_10_i_radr_d,
      wadr_d => vec_rsc_0_10_i_wadr_d,
      we_d => vec_rsc_0_10_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_10_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_10_i_q <= vec_rsc_0_10_q;
  vec_rsc_0_10_radr <= vec_rsc_0_10_i_radr;
  vec_rsc_0_10_d <= vec_rsc_0_10_i_d;
  vec_rsc_0_10_wadr <= vec_rsc_0_10_i_wadr;
  vec_rsc_0_10_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_10_i_q_d <= vec_rsc_0_10_i_q_d_1;
  vec_rsc_0_10_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_10_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_11_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_11_i_q,
      radr => vec_rsc_0_11_i_radr,
      we => vec_rsc_0_11_we,
      d => vec_rsc_0_11_i_d,
      wadr => vec_rsc_0_11_i_wadr,
      d_d => vec_rsc_0_11_i_d_d,
      q_d => vec_rsc_0_11_i_q_d_1,
      radr_d => vec_rsc_0_11_i_radr_d,
      wadr_d => vec_rsc_0_11_i_wadr_d,
      we_d => vec_rsc_0_11_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_11_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_11_i_q <= vec_rsc_0_11_q;
  vec_rsc_0_11_radr <= vec_rsc_0_11_i_radr;
  vec_rsc_0_11_d <= vec_rsc_0_11_i_d;
  vec_rsc_0_11_wadr <= vec_rsc_0_11_i_wadr;
  vec_rsc_0_11_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_11_i_q_d <= vec_rsc_0_11_i_q_d_1;
  vec_rsc_0_11_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_11_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_12_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_12_i_q,
      radr => vec_rsc_0_12_i_radr,
      we => vec_rsc_0_12_we,
      d => vec_rsc_0_12_i_d,
      wadr => vec_rsc_0_12_i_wadr,
      d_d => vec_rsc_0_12_i_d_d,
      q_d => vec_rsc_0_12_i_q_d_1,
      radr_d => vec_rsc_0_12_i_radr_d,
      wadr_d => vec_rsc_0_12_i_wadr_d,
      we_d => vec_rsc_0_12_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_12_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_12_i_q <= vec_rsc_0_12_q;
  vec_rsc_0_12_radr <= vec_rsc_0_12_i_radr;
  vec_rsc_0_12_d <= vec_rsc_0_12_i_d;
  vec_rsc_0_12_wadr <= vec_rsc_0_12_i_wadr;
  vec_rsc_0_12_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_12_i_q_d <= vec_rsc_0_12_i_q_d_1;
  vec_rsc_0_12_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_12_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_13_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_13_i_q,
      radr => vec_rsc_0_13_i_radr,
      we => vec_rsc_0_13_we,
      d => vec_rsc_0_13_i_d,
      wadr => vec_rsc_0_13_i_wadr,
      d_d => vec_rsc_0_13_i_d_d,
      q_d => vec_rsc_0_13_i_q_d_1,
      radr_d => vec_rsc_0_13_i_radr_d,
      wadr_d => vec_rsc_0_13_i_wadr_d,
      we_d => vec_rsc_0_13_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_13_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_13_i_q <= vec_rsc_0_13_q;
  vec_rsc_0_13_radr <= vec_rsc_0_13_i_radr;
  vec_rsc_0_13_d <= vec_rsc_0_13_i_d;
  vec_rsc_0_13_wadr <= vec_rsc_0_13_i_wadr;
  vec_rsc_0_13_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_13_i_q_d <= vec_rsc_0_13_i_q_d_1;
  vec_rsc_0_13_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_13_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_14_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_14_i_q,
      radr => vec_rsc_0_14_i_radr,
      we => vec_rsc_0_14_we,
      d => vec_rsc_0_14_i_d,
      wadr => vec_rsc_0_14_i_wadr,
      d_d => vec_rsc_0_14_i_d_d,
      q_d => vec_rsc_0_14_i_q_d_1,
      radr_d => vec_rsc_0_14_i_radr_d,
      wadr_d => vec_rsc_0_14_i_wadr_d,
      we_d => vec_rsc_0_14_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_14_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_14_i_q <= vec_rsc_0_14_q;
  vec_rsc_0_14_radr <= vec_rsc_0_14_i_radr;
  vec_rsc_0_14_d <= vec_rsc_0_14_i_d;
  vec_rsc_0_14_wadr <= vec_rsc_0_14_i_wadr;
  vec_rsc_0_14_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_14_i_q_d <= vec_rsc_0_14_i_q_d_1;
  vec_rsc_0_14_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_14_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_15_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_15_i_q,
      radr => vec_rsc_0_15_i_radr,
      we => vec_rsc_0_15_we,
      d => vec_rsc_0_15_i_d,
      wadr => vec_rsc_0_15_i_wadr,
      d_d => vec_rsc_0_15_i_d_d,
      q_d => vec_rsc_0_15_i_q_d_1,
      radr_d => vec_rsc_0_15_i_radr_d,
      wadr_d => vec_rsc_0_15_i_wadr_d,
      we_d => vec_rsc_0_15_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_15_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_15_i_q <= vec_rsc_0_15_q;
  vec_rsc_0_15_radr <= vec_rsc_0_15_i_radr;
  vec_rsc_0_15_d <= vec_rsc_0_15_i_d;
  vec_rsc_0_15_wadr <= vec_rsc_0_15_i_wadr;
  vec_rsc_0_15_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_15_i_q_d <= vec_rsc_0_15_i_q_d_1;
  vec_rsc_0_15_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_15_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_16_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_16_i_q,
      radr => vec_rsc_0_16_i_radr,
      we => vec_rsc_0_16_we,
      d => vec_rsc_0_16_i_d,
      wadr => vec_rsc_0_16_i_wadr,
      d_d => vec_rsc_0_16_i_d_d,
      q_d => vec_rsc_0_16_i_q_d_1,
      radr_d => vec_rsc_0_16_i_radr_d,
      wadr_d => vec_rsc_0_16_i_wadr_d,
      we_d => vec_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_16_i_q <= vec_rsc_0_16_q;
  vec_rsc_0_16_radr <= vec_rsc_0_16_i_radr;
  vec_rsc_0_16_d <= vec_rsc_0_16_i_d;
  vec_rsc_0_16_wadr <= vec_rsc_0_16_i_wadr;
  vec_rsc_0_16_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_16_i_q_d <= vec_rsc_0_16_i_q_d_1;
  vec_rsc_0_16_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_16_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_17_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_17_i_q,
      radr => vec_rsc_0_17_i_radr,
      we => vec_rsc_0_17_we,
      d => vec_rsc_0_17_i_d,
      wadr => vec_rsc_0_17_i_wadr,
      d_d => vec_rsc_0_17_i_d_d,
      q_d => vec_rsc_0_17_i_q_d_1,
      radr_d => vec_rsc_0_17_i_radr_d,
      wadr_d => vec_rsc_0_17_i_wadr_d,
      we_d => vec_rsc_0_17_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_17_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_17_i_q <= vec_rsc_0_17_q;
  vec_rsc_0_17_radr <= vec_rsc_0_17_i_radr;
  vec_rsc_0_17_d <= vec_rsc_0_17_i_d;
  vec_rsc_0_17_wadr <= vec_rsc_0_17_i_wadr;
  vec_rsc_0_17_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_17_i_q_d <= vec_rsc_0_17_i_q_d_1;
  vec_rsc_0_17_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_17_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_18_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_18_i_q,
      radr => vec_rsc_0_18_i_radr,
      we => vec_rsc_0_18_we,
      d => vec_rsc_0_18_i_d,
      wadr => vec_rsc_0_18_i_wadr,
      d_d => vec_rsc_0_18_i_d_d,
      q_d => vec_rsc_0_18_i_q_d_1,
      radr_d => vec_rsc_0_18_i_radr_d,
      wadr_d => vec_rsc_0_18_i_wadr_d,
      we_d => vec_rsc_0_18_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_18_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_18_i_q <= vec_rsc_0_18_q;
  vec_rsc_0_18_radr <= vec_rsc_0_18_i_radr;
  vec_rsc_0_18_d <= vec_rsc_0_18_i_d;
  vec_rsc_0_18_wadr <= vec_rsc_0_18_i_wadr;
  vec_rsc_0_18_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_18_i_q_d <= vec_rsc_0_18_i_q_d_1;
  vec_rsc_0_18_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_18_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_19_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_19_i_q,
      radr => vec_rsc_0_19_i_radr,
      we => vec_rsc_0_19_we,
      d => vec_rsc_0_19_i_d,
      wadr => vec_rsc_0_19_i_wadr,
      d_d => vec_rsc_0_19_i_d_d,
      q_d => vec_rsc_0_19_i_q_d_1,
      radr_d => vec_rsc_0_19_i_radr_d,
      wadr_d => vec_rsc_0_19_i_wadr_d,
      we_d => vec_rsc_0_19_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_19_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_19_i_q <= vec_rsc_0_19_q;
  vec_rsc_0_19_radr <= vec_rsc_0_19_i_radr;
  vec_rsc_0_19_d <= vec_rsc_0_19_i_d;
  vec_rsc_0_19_wadr <= vec_rsc_0_19_i_wadr;
  vec_rsc_0_19_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_19_i_q_d <= vec_rsc_0_19_i_q_d_1;
  vec_rsc_0_19_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_19_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_20_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_20_i_q,
      radr => vec_rsc_0_20_i_radr,
      we => vec_rsc_0_20_we,
      d => vec_rsc_0_20_i_d,
      wadr => vec_rsc_0_20_i_wadr,
      d_d => vec_rsc_0_20_i_d_d,
      q_d => vec_rsc_0_20_i_q_d_1,
      radr_d => vec_rsc_0_20_i_radr_d,
      wadr_d => vec_rsc_0_20_i_wadr_d,
      we_d => vec_rsc_0_20_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_20_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_20_i_q <= vec_rsc_0_20_q;
  vec_rsc_0_20_radr <= vec_rsc_0_20_i_radr;
  vec_rsc_0_20_d <= vec_rsc_0_20_i_d;
  vec_rsc_0_20_wadr <= vec_rsc_0_20_i_wadr;
  vec_rsc_0_20_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_20_i_q_d <= vec_rsc_0_20_i_q_d_1;
  vec_rsc_0_20_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_20_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_21_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_21_i_q,
      radr => vec_rsc_0_21_i_radr,
      we => vec_rsc_0_21_we,
      d => vec_rsc_0_21_i_d,
      wadr => vec_rsc_0_21_i_wadr,
      d_d => vec_rsc_0_21_i_d_d,
      q_d => vec_rsc_0_21_i_q_d_1,
      radr_d => vec_rsc_0_21_i_radr_d,
      wadr_d => vec_rsc_0_21_i_wadr_d,
      we_d => vec_rsc_0_21_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_21_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_21_i_q <= vec_rsc_0_21_q;
  vec_rsc_0_21_radr <= vec_rsc_0_21_i_radr;
  vec_rsc_0_21_d <= vec_rsc_0_21_i_d;
  vec_rsc_0_21_wadr <= vec_rsc_0_21_i_wadr;
  vec_rsc_0_21_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_21_i_q_d <= vec_rsc_0_21_i_q_d_1;
  vec_rsc_0_21_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_21_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_22_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_22_i_q,
      radr => vec_rsc_0_22_i_radr,
      we => vec_rsc_0_22_we,
      d => vec_rsc_0_22_i_d,
      wadr => vec_rsc_0_22_i_wadr,
      d_d => vec_rsc_0_22_i_d_d,
      q_d => vec_rsc_0_22_i_q_d_1,
      radr_d => vec_rsc_0_22_i_radr_d,
      wadr_d => vec_rsc_0_22_i_wadr_d,
      we_d => vec_rsc_0_22_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_22_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_22_i_q <= vec_rsc_0_22_q;
  vec_rsc_0_22_radr <= vec_rsc_0_22_i_radr;
  vec_rsc_0_22_d <= vec_rsc_0_22_i_d;
  vec_rsc_0_22_wadr <= vec_rsc_0_22_i_wadr;
  vec_rsc_0_22_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_22_i_q_d <= vec_rsc_0_22_i_q_d_1;
  vec_rsc_0_22_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_22_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_23_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_23_i_q,
      radr => vec_rsc_0_23_i_radr,
      we => vec_rsc_0_23_we,
      d => vec_rsc_0_23_i_d,
      wadr => vec_rsc_0_23_i_wadr,
      d_d => vec_rsc_0_23_i_d_d,
      q_d => vec_rsc_0_23_i_q_d_1,
      radr_d => vec_rsc_0_23_i_radr_d,
      wadr_d => vec_rsc_0_23_i_wadr_d,
      we_d => vec_rsc_0_23_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_23_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_23_i_q <= vec_rsc_0_23_q;
  vec_rsc_0_23_radr <= vec_rsc_0_23_i_radr;
  vec_rsc_0_23_d <= vec_rsc_0_23_i_d;
  vec_rsc_0_23_wadr <= vec_rsc_0_23_i_wadr;
  vec_rsc_0_23_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_23_i_q_d <= vec_rsc_0_23_i_q_d_1;
  vec_rsc_0_23_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_23_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_24_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_24_i_q,
      radr => vec_rsc_0_24_i_radr,
      we => vec_rsc_0_24_we,
      d => vec_rsc_0_24_i_d,
      wadr => vec_rsc_0_24_i_wadr,
      d_d => vec_rsc_0_24_i_d_d,
      q_d => vec_rsc_0_24_i_q_d_1,
      radr_d => vec_rsc_0_24_i_radr_d,
      wadr_d => vec_rsc_0_24_i_wadr_d,
      we_d => vec_rsc_0_24_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_24_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_24_i_q <= vec_rsc_0_24_q;
  vec_rsc_0_24_radr <= vec_rsc_0_24_i_radr;
  vec_rsc_0_24_d <= vec_rsc_0_24_i_d;
  vec_rsc_0_24_wadr <= vec_rsc_0_24_i_wadr;
  vec_rsc_0_24_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_24_i_q_d <= vec_rsc_0_24_i_q_d_1;
  vec_rsc_0_24_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_24_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_25_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_25_i_q,
      radr => vec_rsc_0_25_i_radr,
      we => vec_rsc_0_25_we,
      d => vec_rsc_0_25_i_d,
      wadr => vec_rsc_0_25_i_wadr,
      d_d => vec_rsc_0_25_i_d_d,
      q_d => vec_rsc_0_25_i_q_d_1,
      radr_d => vec_rsc_0_25_i_radr_d,
      wadr_d => vec_rsc_0_25_i_wadr_d,
      we_d => vec_rsc_0_25_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_25_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_25_i_q <= vec_rsc_0_25_q;
  vec_rsc_0_25_radr <= vec_rsc_0_25_i_radr;
  vec_rsc_0_25_d <= vec_rsc_0_25_i_d;
  vec_rsc_0_25_wadr <= vec_rsc_0_25_i_wadr;
  vec_rsc_0_25_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_25_i_q_d <= vec_rsc_0_25_i_q_d_1;
  vec_rsc_0_25_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_25_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_26_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_26_i_q,
      radr => vec_rsc_0_26_i_radr,
      we => vec_rsc_0_26_we,
      d => vec_rsc_0_26_i_d,
      wadr => vec_rsc_0_26_i_wadr,
      d_d => vec_rsc_0_26_i_d_d,
      q_d => vec_rsc_0_26_i_q_d_1,
      radr_d => vec_rsc_0_26_i_radr_d,
      wadr_d => vec_rsc_0_26_i_wadr_d,
      we_d => vec_rsc_0_26_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_26_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_26_i_q <= vec_rsc_0_26_q;
  vec_rsc_0_26_radr <= vec_rsc_0_26_i_radr;
  vec_rsc_0_26_d <= vec_rsc_0_26_i_d;
  vec_rsc_0_26_wadr <= vec_rsc_0_26_i_wadr;
  vec_rsc_0_26_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_26_i_q_d <= vec_rsc_0_26_i_q_d_1;
  vec_rsc_0_26_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_26_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_27_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_27_i_q,
      radr => vec_rsc_0_27_i_radr,
      we => vec_rsc_0_27_we,
      d => vec_rsc_0_27_i_d,
      wadr => vec_rsc_0_27_i_wadr,
      d_d => vec_rsc_0_27_i_d_d,
      q_d => vec_rsc_0_27_i_q_d_1,
      radr_d => vec_rsc_0_27_i_radr_d,
      wadr_d => vec_rsc_0_27_i_wadr_d,
      we_d => vec_rsc_0_27_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_27_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_27_i_q <= vec_rsc_0_27_q;
  vec_rsc_0_27_radr <= vec_rsc_0_27_i_radr;
  vec_rsc_0_27_d <= vec_rsc_0_27_i_d;
  vec_rsc_0_27_wadr <= vec_rsc_0_27_i_wadr;
  vec_rsc_0_27_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_27_i_q_d <= vec_rsc_0_27_i_q_d_1;
  vec_rsc_0_27_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_27_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_28_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_28_i_q,
      radr => vec_rsc_0_28_i_radr,
      we => vec_rsc_0_28_we,
      d => vec_rsc_0_28_i_d,
      wadr => vec_rsc_0_28_i_wadr,
      d_d => vec_rsc_0_28_i_d_d,
      q_d => vec_rsc_0_28_i_q_d_1,
      radr_d => vec_rsc_0_28_i_radr_d,
      wadr_d => vec_rsc_0_28_i_wadr_d,
      we_d => vec_rsc_0_28_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_28_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_28_i_q <= vec_rsc_0_28_q;
  vec_rsc_0_28_radr <= vec_rsc_0_28_i_radr;
  vec_rsc_0_28_d <= vec_rsc_0_28_i_d;
  vec_rsc_0_28_wadr <= vec_rsc_0_28_i_wadr;
  vec_rsc_0_28_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_28_i_q_d <= vec_rsc_0_28_i_q_d_1;
  vec_rsc_0_28_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_28_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_29_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_29_i_q,
      radr => vec_rsc_0_29_i_radr,
      we => vec_rsc_0_29_we,
      d => vec_rsc_0_29_i_d,
      wadr => vec_rsc_0_29_i_wadr,
      d_d => vec_rsc_0_29_i_d_d,
      q_d => vec_rsc_0_29_i_q_d_1,
      radr_d => vec_rsc_0_29_i_radr_d,
      wadr_d => vec_rsc_0_29_i_wadr_d,
      we_d => vec_rsc_0_29_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_29_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_29_i_q <= vec_rsc_0_29_q;
  vec_rsc_0_29_radr <= vec_rsc_0_29_i_radr;
  vec_rsc_0_29_d <= vec_rsc_0_29_i_d;
  vec_rsc_0_29_wadr <= vec_rsc_0_29_i_wadr;
  vec_rsc_0_29_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_29_i_q_d <= vec_rsc_0_29_i_q_d_1;
  vec_rsc_0_29_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_29_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_30_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_30_i_q,
      radr => vec_rsc_0_30_i_radr,
      we => vec_rsc_0_30_we,
      d => vec_rsc_0_30_i_d,
      wadr => vec_rsc_0_30_i_wadr,
      d_d => vec_rsc_0_30_i_d_d,
      q_d => vec_rsc_0_30_i_q_d_1,
      radr_d => vec_rsc_0_30_i_radr_d,
      wadr_d => vec_rsc_0_30_i_wadr_d,
      we_d => vec_rsc_0_30_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_30_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_30_i_q <= vec_rsc_0_30_q;
  vec_rsc_0_30_radr <= vec_rsc_0_30_i_radr;
  vec_rsc_0_30_d <= vec_rsc_0_30_i_d;
  vec_rsc_0_30_wadr <= vec_rsc_0_30_i_wadr;
  vec_rsc_0_30_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_30_i_q_d <= vec_rsc_0_30_i_q_d_1;
  vec_rsc_0_30_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_30_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_31_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_5_64_32_32_64_1_gen
    PORT MAP(
      q => vec_rsc_0_31_i_q,
      radr => vec_rsc_0_31_i_radr,
      we => vec_rsc_0_31_we,
      d => vec_rsc_0_31_i_d,
      wadr => vec_rsc_0_31_i_wadr,
      d_d => vec_rsc_0_31_i_d_d,
      q_d => vec_rsc_0_31_i_q_d_1,
      radr_d => vec_rsc_0_31_i_radr_d,
      wadr_d => vec_rsc_0_31_i_wadr_d,
      we_d => vec_rsc_0_31_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_31_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_31_i_q <= vec_rsc_0_31_q;
  vec_rsc_0_31_radr <= vec_rsc_0_31_i_radr;
  vec_rsc_0_31_d <= vec_rsc_0_31_i_d;
  vec_rsc_0_31_wadr <= vec_rsc_0_31_i_wadr;
  vec_rsc_0_31_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_31_i_q_d <= vec_rsc_0_31_i_q_d_1;
  vec_rsc_0_31_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_31_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  twiddle_rsc_0_0_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_41_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_0_i_q,
      radr => twiddle_rsc_0_0_i_radr,
      q_d => twiddle_rsc_0_0_i_q_d_1,
      radr_d => twiddle_rsc_0_0_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_0_i_q <= twiddle_rsc_0_0_q;
  twiddle_rsc_0_0_radr <= twiddle_rsc_0_0_i_radr;
  twiddle_rsc_0_0_i_q_d <= twiddle_rsc_0_0_i_q_d_1;
  twiddle_rsc_0_0_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_1_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_42_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_1_i_q,
      radr => twiddle_rsc_0_1_i_radr,
      q_d => twiddle_rsc_0_1_i_q_d_1,
      radr_d => twiddle_rsc_0_1_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_1_i_q <= twiddle_rsc_0_1_q;
  twiddle_rsc_0_1_radr <= twiddle_rsc_0_1_i_radr;
  twiddle_rsc_0_1_i_q_d <= twiddle_rsc_0_1_i_q_d_1;
  twiddle_rsc_0_1_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_2_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_43_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_2_i_q,
      radr => twiddle_rsc_0_2_i_radr,
      q_d => twiddle_rsc_0_2_i_q_d_1,
      radr_d => twiddle_rsc_0_2_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_2_i_q <= twiddle_rsc_0_2_q;
  twiddle_rsc_0_2_radr <= twiddle_rsc_0_2_i_radr;
  twiddle_rsc_0_2_i_q_d <= twiddle_rsc_0_2_i_q_d_1;
  twiddle_rsc_0_2_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_3_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_44_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_3_i_q,
      radr => twiddle_rsc_0_3_i_radr,
      q_d => twiddle_rsc_0_3_i_q_d_1,
      radr_d => twiddle_rsc_0_3_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_3_i_q <= twiddle_rsc_0_3_q;
  twiddle_rsc_0_3_radr <= twiddle_rsc_0_3_i_radr;
  twiddle_rsc_0_3_i_q_d <= twiddle_rsc_0_3_i_q_d_1;
  twiddle_rsc_0_3_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_4_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_45_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_4_i_q,
      radr => twiddle_rsc_0_4_i_radr,
      q_d => twiddle_rsc_0_4_i_q_d_1,
      radr_d => twiddle_rsc_0_4_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_4_i_q <= twiddle_rsc_0_4_q;
  twiddle_rsc_0_4_radr <= twiddle_rsc_0_4_i_radr;
  twiddle_rsc_0_4_i_q_d <= twiddle_rsc_0_4_i_q_d_1;
  twiddle_rsc_0_4_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_5_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_46_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_5_i_q,
      radr => twiddle_rsc_0_5_i_radr,
      q_d => twiddle_rsc_0_5_i_q_d_1,
      radr_d => twiddle_rsc_0_5_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_5_i_q <= twiddle_rsc_0_5_q;
  twiddle_rsc_0_5_radr <= twiddle_rsc_0_5_i_radr;
  twiddle_rsc_0_5_i_q_d <= twiddle_rsc_0_5_i_q_d_1;
  twiddle_rsc_0_5_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_6_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_47_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_6_i_q,
      radr => twiddle_rsc_0_6_i_radr,
      q_d => twiddle_rsc_0_6_i_q_d_1,
      radr_d => twiddle_rsc_0_6_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_6_i_q <= twiddle_rsc_0_6_q;
  twiddle_rsc_0_6_radr <= twiddle_rsc_0_6_i_radr;
  twiddle_rsc_0_6_i_q_d <= twiddle_rsc_0_6_i_q_d_1;
  twiddle_rsc_0_6_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_7_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_48_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_7_i_q,
      radr => twiddle_rsc_0_7_i_radr,
      q_d => twiddle_rsc_0_7_i_q_d_1,
      radr_d => twiddle_rsc_0_7_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_7_i_q <= twiddle_rsc_0_7_q;
  twiddle_rsc_0_7_radr <= twiddle_rsc_0_7_i_radr;
  twiddle_rsc_0_7_i_q_d <= twiddle_rsc_0_7_i_q_d_1;
  twiddle_rsc_0_7_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_8_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_49_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_8_i_q,
      radr => twiddle_rsc_0_8_i_radr,
      q_d => twiddle_rsc_0_8_i_q_d_1,
      radr_d => twiddle_rsc_0_8_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_8_i_q <= twiddle_rsc_0_8_q;
  twiddle_rsc_0_8_radr <= twiddle_rsc_0_8_i_radr;
  twiddle_rsc_0_8_i_q_d <= twiddle_rsc_0_8_i_q_d_1;
  twiddle_rsc_0_8_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_9_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_50_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_9_i_q,
      radr => twiddle_rsc_0_9_i_radr,
      q_d => twiddle_rsc_0_9_i_q_d_1,
      radr_d => twiddle_rsc_0_9_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_9_i_q <= twiddle_rsc_0_9_q;
  twiddle_rsc_0_9_radr <= twiddle_rsc_0_9_i_radr;
  twiddle_rsc_0_9_i_q_d <= twiddle_rsc_0_9_i_q_d_1;
  twiddle_rsc_0_9_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_10_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_51_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_10_i_q,
      radr => twiddle_rsc_0_10_i_radr,
      q_d => twiddle_rsc_0_10_i_q_d_1,
      radr_d => twiddle_rsc_0_10_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_10_i_q <= twiddle_rsc_0_10_q;
  twiddle_rsc_0_10_radr <= twiddle_rsc_0_10_i_radr;
  twiddle_rsc_0_10_i_q_d <= twiddle_rsc_0_10_i_q_d_1;
  twiddle_rsc_0_10_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_11_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_52_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_11_i_q,
      radr => twiddle_rsc_0_11_i_radr,
      q_d => twiddle_rsc_0_11_i_q_d_1,
      radr_d => twiddle_rsc_0_11_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_11_i_q <= twiddle_rsc_0_11_q;
  twiddle_rsc_0_11_radr <= twiddle_rsc_0_11_i_radr;
  twiddle_rsc_0_11_i_q_d <= twiddle_rsc_0_11_i_q_d_1;
  twiddle_rsc_0_11_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_12_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_53_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_12_i_q,
      radr => twiddle_rsc_0_12_i_radr,
      q_d => twiddle_rsc_0_12_i_q_d_1,
      radr_d => twiddle_rsc_0_12_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_12_i_q <= twiddle_rsc_0_12_q;
  twiddle_rsc_0_12_radr <= twiddle_rsc_0_12_i_radr;
  twiddle_rsc_0_12_i_q_d <= twiddle_rsc_0_12_i_q_d_1;
  twiddle_rsc_0_12_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_13_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_54_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_13_i_q,
      radr => twiddle_rsc_0_13_i_radr,
      q_d => twiddle_rsc_0_13_i_q_d_1,
      radr_d => twiddle_rsc_0_13_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_13_i_q <= twiddle_rsc_0_13_q;
  twiddle_rsc_0_13_radr <= twiddle_rsc_0_13_i_radr;
  twiddle_rsc_0_13_i_q_d <= twiddle_rsc_0_13_i_q_d_1;
  twiddle_rsc_0_13_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_14_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_55_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_14_i_q,
      radr => twiddle_rsc_0_14_i_radr,
      q_d => twiddle_rsc_0_14_i_q_d_1,
      radr_d => twiddle_rsc_0_14_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_14_i_q <= twiddle_rsc_0_14_q;
  twiddle_rsc_0_14_radr <= twiddle_rsc_0_14_i_radr;
  twiddle_rsc_0_14_i_q_d <= twiddle_rsc_0_14_i_q_d_1;
  twiddle_rsc_0_14_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_15_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_56_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_15_i_q,
      radr => twiddle_rsc_0_15_i_radr,
      q_d => twiddle_rsc_0_15_i_q_d_1,
      radr_d => twiddle_rsc_0_15_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_15_i_q <= twiddle_rsc_0_15_q;
  twiddle_rsc_0_15_radr <= twiddle_rsc_0_15_i_radr;
  twiddle_rsc_0_15_i_q_d <= twiddle_rsc_0_15_i_q_d_1;
  twiddle_rsc_0_15_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_16_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_57_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_16_i_q,
      radr => twiddle_rsc_0_16_i_radr,
      q_d => twiddle_rsc_0_16_i_q_d_1,
      radr_d => twiddle_rsc_0_16_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_16_i_q <= twiddle_rsc_0_16_q;
  twiddle_rsc_0_16_radr <= twiddle_rsc_0_16_i_radr;
  twiddle_rsc_0_16_i_q_d <= twiddle_rsc_0_16_i_q_d_1;
  twiddle_rsc_0_16_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_17_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_58_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_17_i_q,
      radr => twiddle_rsc_0_17_i_radr,
      q_d => twiddle_rsc_0_17_i_q_d_1,
      radr_d => twiddle_rsc_0_17_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_17_i_q <= twiddle_rsc_0_17_q;
  twiddle_rsc_0_17_radr <= twiddle_rsc_0_17_i_radr;
  twiddle_rsc_0_17_i_q_d <= twiddle_rsc_0_17_i_q_d_1;
  twiddle_rsc_0_17_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_18_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_59_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_18_i_q,
      radr => twiddle_rsc_0_18_i_radr,
      q_d => twiddle_rsc_0_18_i_q_d_1,
      radr_d => twiddle_rsc_0_18_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_18_i_q <= twiddle_rsc_0_18_q;
  twiddle_rsc_0_18_radr <= twiddle_rsc_0_18_i_radr;
  twiddle_rsc_0_18_i_q_d <= twiddle_rsc_0_18_i_q_d_1;
  twiddle_rsc_0_18_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_19_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_60_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_19_i_q,
      radr => twiddle_rsc_0_19_i_radr,
      q_d => twiddle_rsc_0_19_i_q_d_1,
      radr_d => twiddle_rsc_0_19_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_19_i_q <= twiddle_rsc_0_19_q;
  twiddle_rsc_0_19_radr <= twiddle_rsc_0_19_i_radr;
  twiddle_rsc_0_19_i_q_d <= twiddle_rsc_0_19_i_q_d_1;
  twiddle_rsc_0_19_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_20_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_61_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_20_i_q,
      radr => twiddle_rsc_0_20_i_radr,
      q_d => twiddle_rsc_0_20_i_q_d_1,
      radr_d => twiddle_rsc_0_20_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_20_i_q <= twiddle_rsc_0_20_q;
  twiddle_rsc_0_20_radr <= twiddle_rsc_0_20_i_radr;
  twiddle_rsc_0_20_i_q_d <= twiddle_rsc_0_20_i_q_d_1;
  twiddle_rsc_0_20_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_21_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_62_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_21_i_q,
      radr => twiddle_rsc_0_21_i_radr,
      q_d => twiddle_rsc_0_21_i_q_d_1,
      radr_d => twiddle_rsc_0_21_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_21_i_q <= twiddle_rsc_0_21_q;
  twiddle_rsc_0_21_radr <= twiddle_rsc_0_21_i_radr;
  twiddle_rsc_0_21_i_q_d <= twiddle_rsc_0_21_i_q_d_1;
  twiddle_rsc_0_21_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_22_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_63_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_22_i_q,
      radr => twiddle_rsc_0_22_i_radr,
      q_d => twiddle_rsc_0_22_i_q_d_1,
      radr_d => twiddle_rsc_0_22_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_22_i_q <= twiddle_rsc_0_22_q;
  twiddle_rsc_0_22_radr <= twiddle_rsc_0_22_i_radr;
  twiddle_rsc_0_22_i_q_d <= twiddle_rsc_0_22_i_q_d_1;
  twiddle_rsc_0_22_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_23_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_64_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_23_i_q,
      radr => twiddle_rsc_0_23_i_radr,
      q_d => twiddle_rsc_0_23_i_q_d_1,
      radr_d => twiddle_rsc_0_23_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_23_i_q <= twiddle_rsc_0_23_q;
  twiddle_rsc_0_23_radr <= twiddle_rsc_0_23_i_radr;
  twiddle_rsc_0_23_i_q_d <= twiddle_rsc_0_23_i_q_d_1;
  twiddle_rsc_0_23_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_24_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_65_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_24_i_q,
      radr => twiddle_rsc_0_24_i_radr,
      q_d => twiddle_rsc_0_24_i_q_d_1,
      radr_d => twiddle_rsc_0_24_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_24_i_q <= twiddle_rsc_0_24_q;
  twiddle_rsc_0_24_radr <= twiddle_rsc_0_24_i_radr;
  twiddle_rsc_0_24_i_q_d <= twiddle_rsc_0_24_i_q_d_1;
  twiddle_rsc_0_24_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_25_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_66_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_25_i_q,
      radr => twiddle_rsc_0_25_i_radr,
      q_d => twiddle_rsc_0_25_i_q_d_1,
      radr_d => twiddle_rsc_0_25_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_25_i_q <= twiddle_rsc_0_25_q;
  twiddle_rsc_0_25_radr <= twiddle_rsc_0_25_i_radr;
  twiddle_rsc_0_25_i_q_d <= twiddle_rsc_0_25_i_q_d_1;
  twiddle_rsc_0_25_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_26_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_67_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_26_i_q,
      radr => twiddle_rsc_0_26_i_radr,
      q_d => twiddle_rsc_0_26_i_q_d_1,
      radr_d => twiddle_rsc_0_26_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_26_i_q <= twiddle_rsc_0_26_q;
  twiddle_rsc_0_26_radr <= twiddle_rsc_0_26_i_radr;
  twiddle_rsc_0_26_i_q_d <= twiddle_rsc_0_26_i_q_d_1;
  twiddle_rsc_0_26_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_27_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_68_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_27_i_q,
      radr => twiddle_rsc_0_27_i_radr,
      q_d => twiddle_rsc_0_27_i_q_d_1,
      radr_d => twiddle_rsc_0_27_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_27_i_q <= twiddle_rsc_0_27_q;
  twiddle_rsc_0_27_radr <= twiddle_rsc_0_27_i_radr;
  twiddle_rsc_0_27_i_q_d <= twiddle_rsc_0_27_i_q_d_1;
  twiddle_rsc_0_27_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_28_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_69_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_28_i_q,
      radr => twiddle_rsc_0_28_i_radr,
      q_d => twiddle_rsc_0_28_i_q_d_1,
      radr_d => twiddle_rsc_0_28_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_28_i_q <= twiddle_rsc_0_28_q;
  twiddle_rsc_0_28_radr <= twiddle_rsc_0_28_i_radr;
  twiddle_rsc_0_28_i_q_d <= twiddle_rsc_0_28_i_q_d_1;
  twiddle_rsc_0_28_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_29_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_70_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_29_i_q,
      radr => twiddle_rsc_0_29_i_radr,
      q_d => twiddle_rsc_0_29_i_q_d_1,
      radr_d => twiddle_rsc_0_29_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_29_i_q <= twiddle_rsc_0_29_q;
  twiddle_rsc_0_29_radr <= twiddle_rsc_0_29_i_radr;
  twiddle_rsc_0_29_i_q_d <= twiddle_rsc_0_29_i_q_d_1;
  twiddle_rsc_0_29_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_30_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_71_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_30_i_q,
      radr => twiddle_rsc_0_30_i_radr,
      q_d => twiddle_rsc_0_30_i_q_d_1,
      radr_d => twiddle_rsc_0_30_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_30_i_q <= twiddle_rsc_0_30_q;
  twiddle_rsc_0_30_radr <= twiddle_rsc_0_30_i_radr;
  twiddle_rsc_0_30_i_q_d <= twiddle_rsc_0_30_i_q_d_1;
  twiddle_rsc_0_30_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_31_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_72_5_64_32_32_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_31_i_q,
      radr => twiddle_rsc_0_31_i_radr,
      q_d => twiddle_rsc_0_31_i_q_d_1,
      radr_d => twiddle_rsc_0_31_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_31_i_q <= twiddle_rsc_0_31_q;
  twiddle_rsc_0_31_radr <= twiddle_rsc_0_31_i_radr;
  twiddle_rsc_0_31_i_q_d <= twiddle_rsc_0_31_i_q_d_1;
  twiddle_rsc_0_31_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  inPlaceNTT_DIF_core_inst : inPlaceNTT_DIF_core
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      vec_rsc_triosy_0_8_lz => vec_rsc_triosy_0_8_lz,
      vec_rsc_triosy_0_9_lz => vec_rsc_triosy_0_9_lz,
      vec_rsc_triosy_0_10_lz => vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz => vec_rsc_triosy_0_11_lz,
      vec_rsc_triosy_0_12_lz => vec_rsc_triosy_0_12_lz,
      vec_rsc_triosy_0_13_lz => vec_rsc_triosy_0_13_lz,
      vec_rsc_triosy_0_14_lz => vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz => vec_rsc_triosy_0_15_lz,
      vec_rsc_triosy_0_16_lz => vec_rsc_triosy_0_16_lz,
      vec_rsc_triosy_0_17_lz => vec_rsc_triosy_0_17_lz,
      vec_rsc_triosy_0_18_lz => vec_rsc_triosy_0_18_lz,
      vec_rsc_triosy_0_19_lz => vec_rsc_triosy_0_19_lz,
      vec_rsc_triosy_0_20_lz => vec_rsc_triosy_0_20_lz,
      vec_rsc_triosy_0_21_lz => vec_rsc_triosy_0_21_lz,
      vec_rsc_triosy_0_22_lz => vec_rsc_triosy_0_22_lz,
      vec_rsc_triosy_0_23_lz => vec_rsc_triosy_0_23_lz,
      vec_rsc_triosy_0_24_lz => vec_rsc_triosy_0_24_lz,
      vec_rsc_triosy_0_25_lz => vec_rsc_triosy_0_25_lz,
      vec_rsc_triosy_0_26_lz => vec_rsc_triosy_0_26_lz,
      vec_rsc_triosy_0_27_lz => vec_rsc_triosy_0_27_lz,
      vec_rsc_triosy_0_28_lz => vec_rsc_triosy_0_28_lz,
      vec_rsc_triosy_0_29_lz => vec_rsc_triosy_0_29_lz,
      vec_rsc_triosy_0_30_lz => vec_rsc_triosy_0_30_lz,
      vec_rsc_triosy_0_31_lz => vec_rsc_triosy_0_31_lz,
      p_rsc_dat => inPlaceNTT_DIF_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_triosy_0_8_lz => twiddle_rsc_triosy_0_8_lz,
      twiddle_rsc_triosy_0_9_lz => twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_triosy_0_10_lz => twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_triosy_0_11_lz => twiddle_rsc_triosy_0_11_lz,
      twiddle_rsc_triosy_0_12_lz => twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_triosy_0_13_lz => twiddle_rsc_triosy_0_13_lz,
      twiddle_rsc_triosy_0_14_lz => twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_triosy_0_15_lz => twiddle_rsc_triosy_0_15_lz,
      twiddle_rsc_triosy_0_16_lz => twiddle_rsc_triosy_0_16_lz,
      twiddle_rsc_triosy_0_17_lz => twiddle_rsc_triosy_0_17_lz,
      twiddle_rsc_triosy_0_18_lz => twiddle_rsc_triosy_0_18_lz,
      twiddle_rsc_triosy_0_19_lz => twiddle_rsc_triosy_0_19_lz,
      twiddle_rsc_triosy_0_20_lz => twiddle_rsc_triosy_0_20_lz,
      twiddle_rsc_triosy_0_21_lz => twiddle_rsc_triosy_0_21_lz,
      twiddle_rsc_triosy_0_22_lz => twiddle_rsc_triosy_0_22_lz,
      twiddle_rsc_triosy_0_23_lz => twiddle_rsc_triosy_0_23_lz,
      twiddle_rsc_triosy_0_24_lz => twiddle_rsc_triosy_0_24_lz,
      twiddle_rsc_triosy_0_25_lz => twiddle_rsc_triosy_0_25_lz,
      twiddle_rsc_triosy_0_26_lz => twiddle_rsc_triosy_0_26_lz,
      twiddle_rsc_triosy_0_27_lz => twiddle_rsc_triosy_0_27_lz,
      twiddle_rsc_triosy_0_28_lz => twiddle_rsc_triosy_0_28_lz,
      twiddle_rsc_triosy_0_29_lz => twiddle_rsc_triosy_0_29_lz,
      twiddle_rsc_triosy_0_30_lz => twiddle_rsc_triosy_0_30_lz,
      twiddle_rsc_triosy_0_31_lz => twiddle_rsc_triosy_0_31_lz,
      vec_rsc_0_0_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d,
      vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d,
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d,
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d,
      vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d,
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d,
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d,
      vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d,
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_8_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d,
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d,
      vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_10_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d,
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_11_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d,
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d,
      vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_13_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d,
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_14_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d,
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d,
      vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_16_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_16_i_q_d,
      vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_17_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_17_i_q_d,
      vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_18_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_18_i_q_d,
      vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_19_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_19_i_q_d,
      vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_20_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_20_i_q_d,
      vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_21_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_21_i_q_d,
      vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_22_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_22_i_q_d,
      vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_23_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_23_i_q_d,
      vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_24_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_24_i_q_d,
      vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_25_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_25_i_q_d,
      vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_26_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_26_i_q_d,
      vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_27_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_27_i_q_d,
      vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_28_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_28_i_q_d,
      vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_29_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_29_i_q_d,
      vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_30_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_30_i_q_d,
      vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_31_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_31_i_q_d,
      vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_0_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d,
      twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d,
      twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d,
      twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d,
      twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d,
      twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d,
      twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d,
      twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d,
      twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_8_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d,
      twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_9_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d,
      twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_10_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d,
      twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_11_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d,
      twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_12_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d,
      twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_13_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d,
      twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_14_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d,
      twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_15_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d,
      twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_16_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_16_i_q_d,
      twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_17_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_17_i_q_d,
      twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_18_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_18_i_q_d,
      twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_19_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_19_i_q_d,
      twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_20_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_20_i_q_d,
      twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_21_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_21_i_q_d,
      twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_22_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_22_i_q_d,
      twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_23_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_23_i_q_d,
      twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_24_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_24_i_q_d,
      twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_25_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_25_i_q_d,
      twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_26_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_26_i_q_d,
      twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_27_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_27_i_q_d,
      twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_28_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_28_i_q_d,
      twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_29_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_29_i_q_d,
      twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_30_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_30_i_q_d,
      twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_31_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_31_i_q_d,
      twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_d_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff,
      vec_rsc_0_0_i_radr_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff,
      vec_rsc_0_0_i_wadr_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff,
      vec_rsc_0_0_i_we_d_pff => vec_rsc_0_0_i_we_d_iff,
      vec_rsc_0_1_i_we_d_pff => vec_rsc_0_1_i_we_d_iff,
      vec_rsc_0_2_i_we_d_pff => vec_rsc_0_2_i_we_d_iff,
      vec_rsc_0_3_i_we_d_pff => vec_rsc_0_3_i_we_d_iff,
      vec_rsc_0_4_i_we_d_pff => vec_rsc_0_4_i_we_d_iff,
      vec_rsc_0_5_i_we_d_pff => vec_rsc_0_5_i_we_d_iff,
      vec_rsc_0_6_i_we_d_pff => vec_rsc_0_6_i_we_d_iff,
      vec_rsc_0_7_i_we_d_pff => vec_rsc_0_7_i_we_d_iff,
      vec_rsc_0_8_i_we_d_pff => vec_rsc_0_8_i_we_d_iff,
      vec_rsc_0_9_i_we_d_pff => vec_rsc_0_9_i_we_d_iff,
      vec_rsc_0_10_i_we_d_pff => vec_rsc_0_10_i_we_d_iff,
      vec_rsc_0_11_i_we_d_pff => vec_rsc_0_11_i_we_d_iff,
      vec_rsc_0_12_i_we_d_pff => vec_rsc_0_12_i_we_d_iff,
      vec_rsc_0_13_i_we_d_pff => vec_rsc_0_13_i_we_d_iff,
      vec_rsc_0_14_i_we_d_pff => vec_rsc_0_14_i_we_d_iff,
      vec_rsc_0_15_i_we_d_pff => vec_rsc_0_15_i_we_d_iff,
      vec_rsc_0_16_i_we_d_pff => vec_rsc_0_16_i_we_d_iff,
      vec_rsc_0_17_i_we_d_pff => vec_rsc_0_17_i_we_d_iff,
      vec_rsc_0_18_i_we_d_pff => vec_rsc_0_18_i_we_d_iff,
      vec_rsc_0_19_i_we_d_pff => vec_rsc_0_19_i_we_d_iff,
      vec_rsc_0_20_i_we_d_pff => vec_rsc_0_20_i_we_d_iff,
      vec_rsc_0_21_i_we_d_pff => vec_rsc_0_21_i_we_d_iff,
      vec_rsc_0_22_i_we_d_pff => vec_rsc_0_22_i_we_d_iff,
      vec_rsc_0_23_i_we_d_pff => vec_rsc_0_23_i_we_d_iff,
      vec_rsc_0_24_i_we_d_pff => vec_rsc_0_24_i_we_d_iff,
      vec_rsc_0_25_i_we_d_pff => vec_rsc_0_25_i_we_d_iff,
      vec_rsc_0_26_i_we_d_pff => vec_rsc_0_26_i_we_d_iff,
      vec_rsc_0_27_i_we_d_pff => vec_rsc_0_27_i_we_d_iff,
      vec_rsc_0_28_i_we_d_pff => vec_rsc_0_28_i_we_d_iff,
      vec_rsc_0_29_i_we_d_pff => vec_rsc_0_29_i_we_d_iff,
      vec_rsc_0_30_i_we_d_pff => vec_rsc_0_30_i_we_d_iff,
      vec_rsc_0_31_i_we_d_pff => vec_rsc_0_31_i_we_d_iff,
      twiddle_rsc_0_0_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d_pff,
      twiddle_rsc_0_1_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff,
      twiddle_rsc_0_2_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff,
      twiddle_rsc_0_4_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff
    );
  inPlaceNTT_DIF_core_inst_p_rsc_dat <= p_rsc_dat;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d <= vec_rsc_0_0_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d <= vec_rsc_0_1_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d <= vec_rsc_0_2_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d <= vec_rsc_0_3_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d <= vec_rsc_0_4_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d <= vec_rsc_0_5_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d <= vec_rsc_0_6_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d <= vec_rsc_0_7_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d <= vec_rsc_0_8_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d <= vec_rsc_0_9_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d <= vec_rsc_0_10_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d <= vec_rsc_0_11_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d <= vec_rsc_0_12_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d <= vec_rsc_0_13_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d <= vec_rsc_0_14_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d <= vec_rsc_0_15_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_16_i_q_d <= vec_rsc_0_16_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_17_i_q_d <= vec_rsc_0_17_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_18_i_q_d <= vec_rsc_0_18_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_19_i_q_d <= vec_rsc_0_19_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_20_i_q_d <= vec_rsc_0_20_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_21_i_q_d <= vec_rsc_0_21_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_22_i_q_d <= vec_rsc_0_22_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_23_i_q_d <= vec_rsc_0_23_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_24_i_q_d <= vec_rsc_0_24_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_25_i_q_d <= vec_rsc_0_25_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_26_i_q_d <= vec_rsc_0_26_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_27_i_q_d <= vec_rsc_0_27_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_28_i_q_d <= vec_rsc_0_28_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_29_i_q_d <= vec_rsc_0_29_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_30_i_q_d <= vec_rsc_0_30_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_31_i_q_d <= vec_rsc_0_31_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d <= twiddle_rsc_0_0_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d <= twiddle_rsc_0_1_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d <= twiddle_rsc_0_2_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d <= twiddle_rsc_0_3_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d <= twiddle_rsc_0_4_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d <= twiddle_rsc_0_5_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d <= twiddle_rsc_0_6_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d <= twiddle_rsc_0_7_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d <= twiddle_rsc_0_8_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d <= twiddle_rsc_0_9_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d <= twiddle_rsc_0_10_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d <= twiddle_rsc_0_11_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d <= twiddle_rsc_0_12_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d <= twiddle_rsc_0_13_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d <= twiddle_rsc_0_14_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d <= twiddle_rsc_0_15_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_16_i_q_d <= twiddle_rsc_0_16_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_17_i_q_d <= twiddle_rsc_0_17_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_18_i_q_d <= twiddle_rsc_0_18_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_19_i_q_d <= twiddle_rsc_0_19_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_20_i_q_d <= twiddle_rsc_0_20_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_21_i_q_d <= twiddle_rsc_0_21_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_22_i_q_d <= twiddle_rsc_0_22_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_23_i_q_d <= twiddle_rsc_0_23_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_24_i_q_d <= twiddle_rsc_0_24_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_25_i_q_d <= twiddle_rsc_0_25_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_26_i_q_d <= twiddle_rsc_0_26_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_27_i_q_d <= twiddle_rsc_0_27_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_28_i_q_d <= twiddle_rsc_0_28_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_29_i_q_d <= twiddle_rsc_0_29_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_30_i_q_d <= twiddle_rsc_0_30_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_31_i_q_d <= twiddle_rsc_0_31_i_q_d;
  vec_rsc_0_0_i_d_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff;
  vec_rsc_0_0_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff;
  vec_rsc_0_0_i_wadr_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff;
  twiddle_rsc_0_0_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d_pff;
  twiddle_rsc_0_1_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff;
  twiddle_rsc_0_2_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff;
  twiddle_rsc_0_4_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff;

END v13;



