
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_out_dreg_pkg_v2 IS

COMPONENT mgc_out_dreg_v2
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_out_dreg_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_out_dreg_v2 IS
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END mgc_out_dreg_v2;

ARCHITECTURE beh OF mgc_out_dreg_v2 IS
BEGIN

  z <= d;

END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_rem IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END mgc_rem;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_rem IS
BEGIN
  z <= std_logic_vector(unsigned(a) rem unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) rem   signed(b));
END beh;

--------> ../td_ccore_solutions/modulo_dev_d3e65941ee7586d7daaa2e36d0d005555a5b_0/rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Thu Aug 26 01:37:25 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    modulo_dev_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_dev_core IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_dev_core;

ARCHITECTURE v1 OF modulo_dev_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL base_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat : STD_LOGIC;
  SIGNAL result_rem_12_cmp_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_a : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_b : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_result_acc_tmp : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_dcpl_1 : STD_LOGIC;
  SIGNAL and_dcpl_2 : STD_LOGIC;
  SIGNAL and_dcpl_3 : STD_LOGIC;
  SIGNAL and_dcpl_4 : STD_LOGIC;
  SIGNAL and_dcpl_6 : STD_LOGIC;
  SIGNAL and_dcpl_8 : STD_LOGIC;
  SIGNAL and_dcpl_9 : STD_LOGIC;
  SIGNAL and_dcpl_11 : STD_LOGIC;
  SIGNAL and_dcpl_13 : STD_LOGIC;
  SIGNAL and_dcpl_18 : STD_LOGIC;
  SIGNAL and_dcpl_26 : STD_LOGIC;
  SIGNAL and_dcpl_27 : STD_LOGIC;
  SIGNAL and_dcpl_28 : STD_LOGIC;
  SIGNAL and_dcpl_29 : STD_LOGIC;
  SIGNAL and_dcpl_30 : STD_LOGIC;
  SIGNAL and_dcpl_31 : STD_LOGIC;
  SIGNAL and_dcpl_32 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_34 : STD_LOGIC;
  SIGNAL and_dcpl_35 : STD_LOGIC;
  SIGNAL and_dcpl_36 : STD_LOGIC;
  SIGNAL and_dcpl_37 : STD_LOGIC;
  SIGNAL and_dcpl_38 : STD_LOGIC;
  SIGNAL and_dcpl_39 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_41 : STD_LOGIC;
  SIGNAL and_dcpl_42 : STD_LOGIC;
  SIGNAL and_dcpl_43 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_47 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL and_dcpl_51 : STD_LOGIC;
  SIGNAL and_dcpl_52 : STD_LOGIC;
  SIGNAL and_dcpl_53 : STD_LOGIC;
  SIGNAL and_dcpl_54 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_56 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_59 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_dcpl_68 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_73 : STD_LOGIC;
  SIGNAL and_dcpl_74 : STD_LOGIC;
  SIGNAL and_dcpl_75 : STD_LOGIC;
  SIGNAL and_dcpl_76 : STD_LOGIC;
  SIGNAL and_dcpl_77 : STD_LOGIC;
  SIGNAL and_dcpl_78 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL and_dcpl_80 : STD_LOGIC;
  SIGNAL and_dcpl_81 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_86 : STD_LOGIC;
  SIGNAL and_dcpl_88 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_96 : STD_LOGIC;
  SIGNAL and_dcpl_98 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_100 : STD_LOGIC;
  SIGNAL and_dcpl_101 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_105 : STD_LOGIC;
  SIGNAL and_dcpl_106 : STD_LOGIC;
  SIGNAL and_dcpl_107 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_113 : STD_LOGIC;
  SIGNAL and_dcpl_114 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_116 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_118 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL and_dcpl_120 : STD_LOGIC;
  SIGNAL and_dcpl_122 : STD_LOGIC;
  SIGNAL and_dcpl_125 : STD_LOGIC;
  SIGNAL and_dcpl_127 : STD_LOGIC;
  SIGNAL and_dcpl_128 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL and_dcpl_130 : STD_LOGIC;
  SIGNAL and_dcpl_131 : STD_LOGIC;
  SIGNAL and_dcpl_132 : STD_LOGIC;
  SIGNAL and_dcpl_133 : STD_LOGIC;
  SIGNAL and_dcpl_134 : STD_LOGIC;
  SIGNAL and_dcpl_135 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_137 : STD_LOGIC;
  SIGNAL and_dcpl_139 : STD_LOGIC;
  SIGNAL and_dcpl_140 : STD_LOGIC;
  SIGNAL and_dcpl_142 : STD_LOGIC;
  SIGNAL and_dcpl_143 : STD_LOGIC;
  SIGNAL and_dcpl_145 : STD_LOGIC;
  SIGNAL and_dcpl_147 : STD_LOGIC;
  SIGNAL and_dcpl_149 : STD_LOGIC;
  SIGNAL and_dcpl_150 : STD_LOGIC;
  SIGNAL and_dcpl_151 : STD_LOGIC;
  SIGNAL and_dcpl_152 : STD_LOGIC;
  SIGNAL and_dcpl_153 : STD_LOGIC;
  SIGNAL and_dcpl_154 : STD_LOGIC;
  SIGNAL and_dcpl_155 : STD_LOGIC;
  SIGNAL and_dcpl_156 : STD_LOGIC;
  SIGNAL and_dcpl_157 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_159 : STD_LOGIC;
  SIGNAL and_dcpl_160 : STD_LOGIC;
  SIGNAL and_dcpl_161 : STD_LOGIC;
  SIGNAL and_dcpl_162 : STD_LOGIC;
  SIGNAL and_dcpl_163 : STD_LOGIC;
  SIGNAL and_dcpl_165 : STD_LOGIC;
  SIGNAL and_dcpl_166 : STD_LOGIC;
  SIGNAL and_dcpl_168 : STD_LOGIC;
  SIGNAL and_dcpl_170 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_176 : STD_LOGIC;
  SIGNAL and_dcpl_177 : STD_LOGIC;
  SIGNAL and_dcpl_178 : STD_LOGIC;
  SIGNAL and_dcpl_179 : STD_LOGIC;
  SIGNAL and_dcpl_180 : STD_LOGIC;
  SIGNAL and_dcpl_181 : STD_LOGIC;
  SIGNAL and_dcpl_182 : STD_LOGIC;
  SIGNAL and_dcpl_183 : STD_LOGIC;
  SIGNAL and_dcpl_184 : STD_LOGIC;
  SIGNAL and_dcpl_185 : STD_LOGIC;
  SIGNAL and_dcpl_186 : STD_LOGIC;
  SIGNAL and_dcpl_187 : STD_LOGIC;
  SIGNAL and_dcpl_188 : STD_LOGIC;
  SIGNAL and_dcpl_189 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_194 : STD_LOGIC;
  SIGNAL and_dcpl_196 : STD_LOGIC;
  SIGNAL and_dcpl_197 : STD_LOGIC;
  SIGNAL and_dcpl_199 : STD_LOGIC;
  SIGNAL and_dcpl_201 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_203 : STD_LOGIC;
  SIGNAL and_dcpl_204 : STD_LOGIC;
  SIGNAL and_dcpl_205 : STD_LOGIC;
  SIGNAL and_dcpl_206 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL and_dcpl_208 : STD_LOGIC;
  SIGNAL and_dcpl_209 : STD_LOGIC;
  SIGNAL and_dcpl_211 : STD_LOGIC;
  SIGNAL and_dcpl_212 : STD_LOGIC;
  SIGNAL and_dcpl_214 : STD_LOGIC;
  SIGNAL and_dcpl_218 : STD_LOGIC;
  SIGNAL and_dcpl_221 : STD_LOGIC;
  SIGNAL and_dcpl_228 : STD_LOGIC;
  SIGNAL and_dcpl_232 : STD_LOGIC;
  SIGNAL and_dcpl_233 : STD_LOGIC;
  SIGNAL and_dcpl_234 : STD_LOGIC;
  SIGNAL and_dcpl_235 : STD_LOGIC;
  SIGNAL and_dcpl_237 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_240 : STD_LOGIC;
  SIGNAL and_dcpl_244 : STD_LOGIC;
  SIGNAL and_dcpl_249 : STD_LOGIC;
  SIGNAL and_dcpl_254 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL and_dcpl_261 : STD_LOGIC;
  SIGNAL and_dcpl_262 : STD_LOGIC;
  SIGNAL and_dcpl_263 : STD_LOGIC;
  SIGNAL or_tmp_2 : STD_LOGIC;
  SIGNAL and_dcpl_269 : STD_LOGIC;
  SIGNAL mux_tmp_1 : STD_LOGIC;
  SIGNAL and_dcpl_275 : STD_LOGIC;
  SIGNAL mux_tmp_3 : STD_LOGIC;
  SIGNAL mux_tmp_4 : STD_LOGIC;
  SIGNAL and_dcpl_281 : STD_LOGIC;
  SIGNAL mux_tmp_6 : STD_LOGIC;
  SIGNAL mux_tmp_7 : STD_LOGIC;
  SIGNAL mux_tmp_8 : STD_LOGIC;
  SIGNAL and_dcpl_287 : STD_LOGIC;
  SIGNAL mux_tmp_10 : STD_LOGIC;
  SIGNAL mux_tmp_11 : STD_LOGIC;
  SIGNAL mux_tmp_12 : STD_LOGIC;
  SIGNAL mux_tmp_13 : STD_LOGIC;
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL mux_tmp_15 : STD_LOGIC;
  SIGNAL mux_tmp_16 : STD_LOGIC;
  SIGNAL mux_tmp_17 : STD_LOGIC;
  SIGNAL mux_tmp_18 : STD_LOGIC;
  SIGNAL mux_tmp_19 : STD_LOGIC;
  SIGNAL and_dcpl_299 : STD_LOGIC;
  SIGNAL mux_tmp_21 : STD_LOGIC;
  SIGNAL mux_tmp_22 : STD_LOGIC;
  SIGNAL mux_tmp_23 : STD_LOGIC;
  SIGNAL mux_tmp_24 : STD_LOGIC;
  SIGNAL mux_tmp_25 : STD_LOGIC;
  SIGNAL mux_tmp_26 : STD_LOGIC;
  SIGNAL and_dcpl_305 : STD_LOGIC;
  SIGNAL mux_tmp_28 : STD_LOGIC;
  SIGNAL mux_tmp_29 : STD_LOGIC;
  SIGNAL mux_tmp_30 : STD_LOGIC;
  SIGNAL mux_tmp_31 : STD_LOGIC;
  SIGNAL mux_tmp_32 : STD_LOGIC;
  SIGNAL mux_tmp_33 : STD_LOGIC;
  SIGNAL mux_tmp_34 : STD_LOGIC;
  SIGNAL and_dcpl_311 : STD_LOGIC;
  SIGNAL and_tmp_6 : STD_LOGIC;
  SIGNAL mux_tmp_36 : STD_LOGIC;
  SIGNAL mux_tmp_37 : STD_LOGIC;
  SIGNAL and_dcpl_318 : STD_LOGIC;
  SIGNAL and_dcpl_319 : STD_LOGIC;
  SIGNAL or_tmp_102 : STD_LOGIC;
  SIGNAL and_dcpl_322 : STD_LOGIC;
  SIGNAL mux_tmp_39 : STD_LOGIC;
  SIGNAL and_dcpl_325 : STD_LOGIC;
  SIGNAL mux_tmp_41 : STD_LOGIC;
  SIGNAL mux_tmp_42 : STD_LOGIC;
  SIGNAL and_dcpl_329 : STD_LOGIC;
  SIGNAL mux_tmp_44 : STD_LOGIC;
  SIGNAL mux_tmp_45 : STD_LOGIC;
  SIGNAL mux_tmp_46 : STD_LOGIC;
  SIGNAL and_dcpl_333 : STD_LOGIC;
  SIGNAL mux_tmp_48 : STD_LOGIC;
  SIGNAL mux_tmp_49 : STD_LOGIC;
  SIGNAL mux_tmp_50 : STD_LOGIC;
  SIGNAL mux_tmp_51 : STD_LOGIC;
  SIGNAL and_dcpl_337 : STD_LOGIC;
  SIGNAL mux_tmp_53 : STD_LOGIC;
  SIGNAL mux_tmp_54 : STD_LOGIC;
  SIGNAL mux_tmp_55 : STD_LOGIC;
  SIGNAL mux_tmp_56 : STD_LOGIC;
  SIGNAL mux_tmp_57 : STD_LOGIC;
  SIGNAL and_dcpl_341 : STD_LOGIC;
  SIGNAL mux_tmp_59 : STD_LOGIC;
  SIGNAL mux_tmp_60 : STD_LOGIC;
  SIGNAL mux_tmp_61 : STD_LOGIC;
  SIGNAL mux_tmp_62 : STD_LOGIC;
  SIGNAL mux_tmp_63 : STD_LOGIC;
  SIGNAL mux_tmp_64 : STD_LOGIC;
  SIGNAL and_dcpl_344 : STD_LOGIC;
  SIGNAL mux_tmp_66 : STD_LOGIC;
  SIGNAL mux_tmp_67 : STD_LOGIC;
  SIGNAL mux_tmp_68 : STD_LOGIC;
  SIGNAL mux_tmp_69 : STD_LOGIC;
  SIGNAL mux_tmp_70 : STD_LOGIC;
  SIGNAL mux_tmp_71 : STD_LOGIC;
  SIGNAL mux_tmp_72 : STD_LOGIC;
  SIGNAL and_dcpl_347 : STD_LOGIC;
  SIGNAL and_tmp_13 : STD_LOGIC;
  SIGNAL mux_tmp_74 : STD_LOGIC;
  SIGNAL mux_tmp_75 : STD_LOGIC;
  SIGNAL and_dcpl_352 : STD_LOGIC;
  SIGNAL and_dcpl_353 : STD_LOGIC;
  SIGNAL or_tmp_202 : STD_LOGIC;
  SIGNAL and_dcpl_357 : STD_LOGIC;
  SIGNAL mux_tmp_77 : STD_LOGIC;
  SIGNAL and_dcpl_361 : STD_LOGIC;
  SIGNAL mux_tmp_79 : STD_LOGIC;
  SIGNAL mux_tmp_80 : STD_LOGIC;
  SIGNAL and_dcpl_364 : STD_LOGIC;
  SIGNAL mux_tmp_82 : STD_LOGIC;
  SIGNAL mux_tmp_83 : STD_LOGIC;
  SIGNAL mux_tmp_84 : STD_LOGIC;
  SIGNAL and_dcpl_367 : STD_LOGIC;
  SIGNAL mux_tmp_86 : STD_LOGIC;
  SIGNAL mux_tmp_87 : STD_LOGIC;
  SIGNAL mux_tmp_88 : STD_LOGIC;
  SIGNAL mux_tmp_89 : STD_LOGIC;
  SIGNAL and_dcpl_370 : STD_LOGIC;
  SIGNAL mux_tmp_91 : STD_LOGIC;
  SIGNAL mux_tmp_92 : STD_LOGIC;
  SIGNAL mux_tmp_93 : STD_LOGIC;
  SIGNAL mux_tmp_94 : STD_LOGIC;
  SIGNAL mux_tmp_95 : STD_LOGIC;
  SIGNAL and_dcpl_373 : STD_LOGIC;
  SIGNAL mux_tmp_97 : STD_LOGIC;
  SIGNAL mux_tmp_98 : STD_LOGIC;
  SIGNAL mux_tmp_99 : STD_LOGIC;
  SIGNAL mux_tmp_100 : STD_LOGIC;
  SIGNAL mux_tmp_101 : STD_LOGIC;
  SIGNAL mux_tmp_102 : STD_LOGIC;
  SIGNAL and_dcpl_377 : STD_LOGIC;
  SIGNAL mux_tmp_104 : STD_LOGIC;
  SIGNAL mux_tmp_105 : STD_LOGIC;
  SIGNAL mux_tmp_106 : STD_LOGIC;
  SIGNAL mux_tmp_107 : STD_LOGIC;
  SIGNAL mux_tmp_108 : STD_LOGIC;
  SIGNAL mux_tmp_109 : STD_LOGIC;
  SIGNAL mux_tmp_110 : STD_LOGIC;
  SIGNAL and_dcpl_381 : STD_LOGIC;
  SIGNAL and_tmp_20 : STD_LOGIC;
  SIGNAL mux_tmp_112 : STD_LOGIC;
  SIGNAL mux_tmp_113 : STD_LOGIC;
  SIGNAL and_dcpl_386 : STD_LOGIC;
  SIGNAL and_dcpl_387 : STD_LOGIC;
  SIGNAL or_tmp_302 : STD_LOGIC;
  SIGNAL and_dcpl_390 : STD_LOGIC;
  SIGNAL mux_tmp_115 : STD_LOGIC;
  SIGNAL and_dcpl_393 : STD_LOGIC;
  SIGNAL mux_tmp_117 : STD_LOGIC;
  SIGNAL mux_tmp_118 : STD_LOGIC;
  SIGNAL and_dcpl_396 : STD_LOGIC;
  SIGNAL mux_tmp_120 : STD_LOGIC;
  SIGNAL mux_tmp_121 : STD_LOGIC;
  SIGNAL mux_tmp_122 : STD_LOGIC;
  SIGNAL and_dcpl_399 : STD_LOGIC;
  SIGNAL mux_tmp_124 : STD_LOGIC;
  SIGNAL mux_tmp_125 : STD_LOGIC;
  SIGNAL mux_tmp_126 : STD_LOGIC;
  SIGNAL mux_tmp_127 : STD_LOGIC;
  SIGNAL and_dcpl_402 : STD_LOGIC;
  SIGNAL mux_tmp_129 : STD_LOGIC;
  SIGNAL mux_tmp_130 : STD_LOGIC;
  SIGNAL mux_tmp_131 : STD_LOGIC;
  SIGNAL mux_tmp_132 : STD_LOGIC;
  SIGNAL mux_tmp_133 : STD_LOGIC;
  SIGNAL and_dcpl_405 : STD_LOGIC;
  SIGNAL mux_tmp_135 : STD_LOGIC;
  SIGNAL mux_tmp_136 : STD_LOGIC;
  SIGNAL mux_tmp_137 : STD_LOGIC;
  SIGNAL mux_tmp_138 : STD_LOGIC;
  SIGNAL mux_tmp_139 : STD_LOGIC;
  SIGNAL mux_tmp_140 : STD_LOGIC;
  SIGNAL and_dcpl_408 : STD_LOGIC;
  SIGNAL mux_tmp_142 : STD_LOGIC;
  SIGNAL mux_tmp_143 : STD_LOGIC;
  SIGNAL mux_tmp_144 : STD_LOGIC;
  SIGNAL mux_tmp_145 : STD_LOGIC;
  SIGNAL mux_tmp_146 : STD_LOGIC;
  SIGNAL mux_tmp_147 : STD_LOGIC;
  SIGNAL mux_tmp_148 : STD_LOGIC;
  SIGNAL and_dcpl_411 : STD_LOGIC;
  SIGNAL and_tmp_27 : STD_LOGIC;
  SIGNAL mux_tmp_150 : STD_LOGIC;
  SIGNAL mux_tmp_151 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL and_dcpl_418 : STD_LOGIC;
  SIGNAL or_tmp_402 : STD_LOGIC;
  SIGNAL and_dcpl_422 : STD_LOGIC;
  SIGNAL mux_tmp_153 : STD_LOGIC;
  SIGNAL and_dcpl_426 : STD_LOGIC;
  SIGNAL mux_tmp_155 : STD_LOGIC;
  SIGNAL mux_tmp_156 : STD_LOGIC;
  SIGNAL and_dcpl_430 : STD_LOGIC;
  SIGNAL mux_tmp_158 : STD_LOGIC;
  SIGNAL mux_tmp_159 : STD_LOGIC;
  SIGNAL mux_tmp_160 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL mux_tmp_162 : STD_LOGIC;
  SIGNAL mux_tmp_163 : STD_LOGIC;
  SIGNAL mux_tmp_164 : STD_LOGIC;
  SIGNAL mux_tmp_165 : STD_LOGIC;
  SIGNAL and_dcpl_437 : STD_LOGIC;
  SIGNAL mux_tmp_167 : STD_LOGIC;
  SIGNAL mux_tmp_168 : STD_LOGIC;
  SIGNAL mux_tmp_169 : STD_LOGIC;
  SIGNAL mux_tmp_170 : STD_LOGIC;
  SIGNAL mux_tmp_171 : STD_LOGIC;
  SIGNAL and_dcpl_441 : STD_LOGIC;
  SIGNAL mux_tmp_173 : STD_LOGIC;
  SIGNAL mux_tmp_174 : STD_LOGIC;
  SIGNAL mux_tmp_175 : STD_LOGIC;
  SIGNAL mux_tmp_176 : STD_LOGIC;
  SIGNAL mux_tmp_177 : STD_LOGIC;
  SIGNAL mux_tmp_178 : STD_LOGIC;
  SIGNAL and_dcpl_444 : STD_LOGIC;
  SIGNAL mux_tmp_180 : STD_LOGIC;
  SIGNAL mux_tmp_181 : STD_LOGIC;
  SIGNAL mux_tmp_182 : STD_LOGIC;
  SIGNAL mux_tmp_183 : STD_LOGIC;
  SIGNAL mux_tmp_184 : STD_LOGIC;
  SIGNAL mux_tmp_185 : STD_LOGIC;
  SIGNAL mux_tmp_186 : STD_LOGIC;
  SIGNAL and_dcpl_447 : STD_LOGIC;
  SIGNAL and_tmp_34 : STD_LOGIC;
  SIGNAL mux_tmp_188 : STD_LOGIC;
  SIGNAL mux_tmp_189 : STD_LOGIC;
  SIGNAL and_dcpl_452 : STD_LOGIC;
  SIGNAL or_tmp_502 : STD_LOGIC;
  SIGNAL and_dcpl_455 : STD_LOGIC;
  SIGNAL mux_tmp_191 : STD_LOGIC;
  SIGNAL and_dcpl_458 : STD_LOGIC;
  SIGNAL mux_tmp_193 : STD_LOGIC;
  SIGNAL mux_tmp_194 : STD_LOGIC;
  SIGNAL and_dcpl_462 : STD_LOGIC;
  SIGNAL mux_tmp_196 : STD_LOGIC;
  SIGNAL mux_tmp_197 : STD_LOGIC;
  SIGNAL mux_tmp_198 : STD_LOGIC;
  SIGNAL and_dcpl_464 : STD_LOGIC;
  SIGNAL mux_tmp_200 : STD_LOGIC;
  SIGNAL mux_tmp_201 : STD_LOGIC;
  SIGNAL mux_tmp_202 : STD_LOGIC;
  SIGNAL mux_tmp_203 : STD_LOGIC;
  SIGNAL and_dcpl_468 : STD_LOGIC;
  SIGNAL mux_tmp_205 : STD_LOGIC;
  SIGNAL mux_tmp_206 : STD_LOGIC;
  SIGNAL mux_tmp_207 : STD_LOGIC;
  SIGNAL mux_tmp_208 : STD_LOGIC;
  SIGNAL mux_tmp_209 : STD_LOGIC;
  SIGNAL and_dcpl_472 : STD_LOGIC;
  SIGNAL mux_tmp_211 : STD_LOGIC;
  SIGNAL mux_tmp_212 : STD_LOGIC;
  SIGNAL mux_tmp_213 : STD_LOGIC;
  SIGNAL mux_tmp_214 : STD_LOGIC;
  SIGNAL mux_tmp_215 : STD_LOGIC;
  SIGNAL mux_tmp_216 : STD_LOGIC;
  SIGNAL and_dcpl_474 : STD_LOGIC;
  SIGNAL mux_tmp_218 : STD_LOGIC;
  SIGNAL mux_tmp_219 : STD_LOGIC;
  SIGNAL mux_tmp_220 : STD_LOGIC;
  SIGNAL mux_tmp_221 : STD_LOGIC;
  SIGNAL mux_tmp_222 : STD_LOGIC;
  SIGNAL mux_tmp_223 : STD_LOGIC;
  SIGNAL mux_tmp_224 : STD_LOGIC;
  SIGNAL and_dcpl_476 : STD_LOGIC;
  SIGNAL and_tmp_41 : STD_LOGIC;
  SIGNAL mux_tmp_226 : STD_LOGIC;
  SIGNAL mux_tmp_227 : STD_LOGIC;
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL or_tmp_602 : STD_LOGIC;
  SIGNAL and_dcpl_484 : STD_LOGIC;
  SIGNAL mux_tmp_229 : STD_LOGIC;
  SIGNAL and_dcpl_488 : STD_LOGIC;
  SIGNAL mux_tmp_231 : STD_LOGIC;
  SIGNAL mux_tmp_232 : STD_LOGIC;
  SIGNAL and_dcpl_491 : STD_LOGIC;
  SIGNAL mux_tmp_234 : STD_LOGIC;
  SIGNAL mux_tmp_235 : STD_LOGIC;
  SIGNAL mux_tmp_236 : STD_LOGIC;
  SIGNAL and_dcpl_493 : STD_LOGIC;
  SIGNAL mux_tmp_238 : STD_LOGIC;
  SIGNAL mux_tmp_239 : STD_LOGIC;
  SIGNAL mux_tmp_240 : STD_LOGIC;
  SIGNAL mux_tmp_241 : STD_LOGIC;
  SIGNAL and_dcpl_496 : STD_LOGIC;
  SIGNAL mux_tmp_243 : STD_LOGIC;
  SIGNAL mux_tmp_244 : STD_LOGIC;
  SIGNAL mux_tmp_245 : STD_LOGIC;
  SIGNAL mux_tmp_246 : STD_LOGIC;
  SIGNAL mux_tmp_247 : STD_LOGIC;
  SIGNAL and_dcpl_499 : STD_LOGIC;
  SIGNAL mux_tmp_249 : STD_LOGIC;
  SIGNAL mux_tmp_250 : STD_LOGIC;
  SIGNAL mux_tmp_251 : STD_LOGIC;
  SIGNAL mux_tmp_252 : STD_LOGIC;
  SIGNAL mux_tmp_253 : STD_LOGIC;
  SIGNAL mux_tmp_254 : STD_LOGIC;
  SIGNAL and_dcpl_501 : STD_LOGIC;
  SIGNAL mux_tmp_256 : STD_LOGIC;
  SIGNAL mux_tmp_257 : STD_LOGIC;
  SIGNAL mux_tmp_258 : STD_LOGIC;
  SIGNAL mux_tmp_259 : STD_LOGIC;
  SIGNAL mux_tmp_260 : STD_LOGIC;
  SIGNAL mux_tmp_261 : STD_LOGIC;
  SIGNAL mux_tmp_262 : STD_LOGIC;
  SIGNAL and_dcpl_503 : STD_LOGIC;
  SIGNAL and_tmp_48 : STD_LOGIC;
  SIGNAL mux_tmp_264 : STD_LOGIC;
  SIGNAL mux_tmp_265 : STD_LOGIC;
  SIGNAL and_dcpl_507 : STD_LOGIC;
  SIGNAL or_tmp_702 : STD_LOGIC;
  SIGNAL and_dcpl_510 : STD_LOGIC;
  SIGNAL mux_tmp_267 : STD_LOGIC;
  SIGNAL and_dcpl_513 : STD_LOGIC;
  SIGNAL mux_tmp_269 : STD_LOGIC;
  SIGNAL mux_tmp_270 : STD_LOGIC;
  SIGNAL and_dcpl_516 : STD_LOGIC;
  SIGNAL mux_tmp_272 : STD_LOGIC;
  SIGNAL mux_tmp_273 : STD_LOGIC;
  SIGNAL mux_tmp_274 : STD_LOGIC;
  SIGNAL and_dcpl_518 : STD_LOGIC;
  SIGNAL mux_tmp_276 : STD_LOGIC;
  SIGNAL mux_tmp_277 : STD_LOGIC;
  SIGNAL mux_tmp_278 : STD_LOGIC;
  SIGNAL mux_tmp_279 : STD_LOGIC;
  SIGNAL and_dcpl_521 : STD_LOGIC;
  SIGNAL mux_tmp_281 : STD_LOGIC;
  SIGNAL mux_tmp_282 : STD_LOGIC;
  SIGNAL mux_tmp_283 : STD_LOGIC;
  SIGNAL mux_tmp_284 : STD_LOGIC;
  SIGNAL mux_tmp_285 : STD_LOGIC;
  SIGNAL and_dcpl_524 : STD_LOGIC;
  SIGNAL mux_tmp_287 : STD_LOGIC;
  SIGNAL mux_tmp_288 : STD_LOGIC;
  SIGNAL mux_tmp_289 : STD_LOGIC;
  SIGNAL mux_tmp_290 : STD_LOGIC;
  SIGNAL mux_tmp_291 : STD_LOGIC;
  SIGNAL mux_tmp_292 : STD_LOGIC;
  SIGNAL and_dcpl_526 : STD_LOGIC;
  SIGNAL mux_tmp_294 : STD_LOGIC;
  SIGNAL mux_tmp_295 : STD_LOGIC;
  SIGNAL mux_tmp_296 : STD_LOGIC;
  SIGNAL mux_tmp_297 : STD_LOGIC;
  SIGNAL mux_tmp_298 : STD_LOGIC;
  SIGNAL mux_tmp_299 : STD_LOGIC;
  SIGNAL mux_tmp_300 : STD_LOGIC;
  SIGNAL and_dcpl_528 : STD_LOGIC;
  SIGNAL and_tmp_55 : STD_LOGIC;
  SIGNAL mux_tmp_302 : STD_LOGIC;
  SIGNAL mux_tmp_303 : STD_LOGIC;
  SIGNAL and_dcpl_532 : STD_LOGIC;
  SIGNAL and_dcpl_533 : STD_LOGIC;
  SIGNAL not_tmp_645 : STD_LOGIC;
  SIGNAL or_tmp_801 : STD_LOGIC;
  SIGNAL and_dcpl_536 : STD_LOGIC;
  SIGNAL mux_tmp_305 : STD_LOGIC;
  SIGNAL and_dcpl_539 : STD_LOGIC;
  SIGNAL mux_tmp_307 : STD_LOGIC;
  SIGNAL mux_tmp_308 : STD_LOGIC;
  SIGNAL and_dcpl_542 : STD_LOGIC;
  SIGNAL mux_tmp_310 : STD_LOGIC;
  SIGNAL mux_tmp_311 : STD_LOGIC;
  SIGNAL mux_tmp_312 : STD_LOGIC;
  SIGNAL and_dcpl_546 : STD_LOGIC;
  SIGNAL mux_tmp_314 : STD_LOGIC;
  SIGNAL mux_tmp_315 : STD_LOGIC;
  SIGNAL mux_tmp_316 : STD_LOGIC;
  SIGNAL mux_tmp_317 : STD_LOGIC;
  SIGNAL and_dcpl_549 : STD_LOGIC;
  SIGNAL mux_tmp_319 : STD_LOGIC;
  SIGNAL mux_tmp_320 : STD_LOGIC;
  SIGNAL mux_tmp_321 : STD_LOGIC;
  SIGNAL mux_tmp_322 : STD_LOGIC;
  SIGNAL mux_tmp_323 : STD_LOGIC;
  SIGNAL and_dcpl_552 : STD_LOGIC;
  SIGNAL mux_tmp_325 : STD_LOGIC;
  SIGNAL mux_tmp_326 : STD_LOGIC;
  SIGNAL mux_tmp_327 : STD_LOGIC;
  SIGNAL mux_tmp_328 : STD_LOGIC;
  SIGNAL mux_tmp_329 : STD_LOGIC;
  SIGNAL mux_tmp_330 : STD_LOGIC;
  SIGNAL and_dcpl_556 : STD_LOGIC;
  SIGNAL mux_tmp_332 : STD_LOGIC;
  SIGNAL mux_tmp_333 : STD_LOGIC;
  SIGNAL mux_tmp_334 : STD_LOGIC;
  SIGNAL mux_tmp_335 : STD_LOGIC;
  SIGNAL mux_tmp_336 : STD_LOGIC;
  SIGNAL mux_tmp_337 : STD_LOGIC;
  SIGNAL mux_tmp_338 : STD_LOGIC;
  SIGNAL and_dcpl_560 : STD_LOGIC;
  SIGNAL or_tmp_897 : STD_LOGIC;
  SIGNAL mux_tmp_340 : STD_LOGIC;
  SIGNAL mux_tmp_341 : STD_LOGIC;
  SIGNAL mux_tmp_342 : STD_LOGIC;
  SIGNAL mux_tmp_343 : STD_LOGIC;
  SIGNAL mux_tmp_344 : STD_LOGIC;
  SIGNAL mux_tmp_345 : STD_LOGIC;
  SIGNAL mux_tmp_346 : STD_LOGIC;
  SIGNAL mux_tmp_347 : STD_LOGIC;
  SIGNAL mux_tmp_348 : STD_LOGIC;
  SIGNAL and_dcpl_566 : STD_LOGIC;
  SIGNAL or_tmp_909 : STD_LOGIC;
  SIGNAL and_dcpl_568 : STD_LOGIC;
  SIGNAL mux_tmp_350 : STD_LOGIC;
  SIGNAL and_dcpl_570 : STD_LOGIC;
  SIGNAL mux_tmp_352 : STD_LOGIC;
  SIGNAL mux_tmp_353 : STD_LOGIC;
  SIGNAL and_dcpl_572 : STD_LOGIC;
  SIGNAL mux_tmp_355 : STD_LOGIC;
  SIGNAL mux_tmp_356 : STD_LOGIC;
  SIGNAL mux_tmp_357 : STD_LOGIC;
  SIGNAL and_dcpl_576 : STD_LOGIC;
  SIGNAL mux_tmp_359 : STD_LOGIC;
  SIGNAL mux_tmp_360 : STD_LOGIC;
  SIGNAL mux_tmp_361 : STD_LOGIC;
  SIGNAL mux_tmp_362 : STD_LOGIC;
  SIGNAL and_dcpl_578 : STD_LOGIC;
  SIGNAL mux_tmp_364 : STD_LOGIC;
  SIGNAL mux_tmp_365 : STD_LOGIC;
  SIGNAL mux_tmp_366 : STD_LOGIC;
  SIGNAL mux_tmp_367 : STD_LOGIC;
  SIGNAL mux_tmp_368 : STD_LOGIC;
  SIGNAL and_dcpl_580 : STD_LOGIC;
  SIGNAL mux_tmp_370 : STD_LOGIC;
  SIGNAL mux_tmp_371 : STD_LOGIC;
  SIGNAL mux_tmp_372 : STD_LOGIC;
  SIGNAL mux_tmp_373 : STD_LOGIC;
  SIGNAL mux_tmp_374 : STD_LOGIC;
  SIGNAL mux_tmp_375 : STD_LOGIC;
  SIGNAL and_dcpl_583 : STD_LOGIC;
  SIGNAL mux_tmp_377 : STD_LOGIC;
  SIGNAL mux_tmp_378 : STD_LOGIC;
  SIGNAL mux_tmp_379 : STD_LOGIC;
  SIGNAL mux_tmp_380 : STD_LOGIC;
  SIGNAL mux_tmp_381 : STD_LOGIC;
  SIGNAL mux_tmp_382 : STD_LOGIC;
  SIGNAL mux_tmp_383 : STD_LOGIC;
  SIGNAL and_dcpl_586 : STD_LOGIC;
  SIGNAL or_tmp_1005 : STD_LOGIC;
  SIGNAL mux_tmp_385 : STD_LOGIC;
  SIGNAL mux_tmp_386 : STD_LOGIC;
  SIGNAL mux_tmp_387 : STD_LOGIC;
  SIGNAL mux_tmp_388 : STD_LOGIC;
  SIGNAL mux_tmp_389 : STD_LOGIC;
  SIGNAL mux_tmp_390 : STD_LOGIC;
  SIGNAL mux_tmp_391 : STD_LOGIC;
  SIGNAL mux_tmp_392 : STD_LOGIC;
  SIGNAL mux_tmp_393 : STD_LOGIC;
  SIGNAL and_dcpl_590 : STD_LOGIC;
  SIGNAL or_tmp_1017 : STD_LOGIC;
  SIGNAL and_dcpl_592 : STD_LOGIC;
  SIGNAL mux_tmp_395 : STD_LOGIC;
  SIGNAL and_dcpl_594 : STD_LOGIC;
  SIGNAL mux_tmp_397 : STD_LOGIC;
  SIGNAL mux_tmp_398 : STD_LOGIC;
  SIGNAL and_dcpl_596 : STD_LOGIC;
  SIGNAL mux_tmp_400 : STD_LOGIC;
  SIGNAL mux_tmp_401 : STD_LOGIC;
  SIGNAL mux_tmp_402 : STD_LOGIC;
  SIGNAL and_dcpl_599 : STD_LOGIC;
  SIGNAL mux_tmp_404 : STD_LOGIC;
  SIGNAL mux_tmp_405 : STD_LOGIC;
  SIGNAL mux_tmp_406 : STD_LOGIC;
  SIGNAL mux_tmp_407 : STD_LOGIC;
  SIGNAL and_dcpl_601 : STD_LOGIC;
  SIGNAL mux_tmp_409 : STD_LOGIC;
  SIGNAL mux_tmp_410 : STD_LOGIC;
  SIGNAL mux_tmp_411 : STD_LOGIC;
  SIGNAL mux_tmp_412 : STD_LOGIC;
  SIGNAL mux_tmp_413 : STD_LOGIC;
  SIGNAL and_dcpl_603 : STD_LOGIC;
  SIGNAL mux_tmp_415 : STD_LOGIC;
  SIGNAL mux_tmp_416 : STD_LOGIC;
  SIGNAL mux_tmp_417 : STD_LOGIC;
  SIGNAL mux_tmp_418 : STD_LOGIC;
  SIGNAL mux_tmp_419 : STD_LOGIC;
  SIGNAL mux_tmp_420 : STD_LOGIC;
  SIGNAL and_dcpl_607 : STD_LOGIC;
  SIGNAL mux_tmp_422 : STD_LOGIC;
  SIGNAL mux_tmp_423 : STD_LOGIC;
  SIGNAL mux_tmp_424 : STD_LOGIC;
  SIGNAL mux_tmp_425 : STD_LOGIC;
  SIGNAL mux_tmp_426 : STD_LOGIC;
  SIGNAL mux_tmp_427 : STD_LOGIC;
  SIGNAL mux_tmp_428 : STD_LOGIC;
  SIGNAL and_dcpl_611 : STD_LOGIC;
  SIGNAL or_tmp_1113 : STD_LOGIC;
  SIGNAL mux_tmp_430 : STD_LOGIC;
  SIGNAL mux_tmp_431 : STD_LOGIC;
  SIGNAL mux_tmp_432 : STD_LOGIC;
  SIGNAL mux_tmp_433 : STD_LOGIC;
  SIGNAL mux_tmp_434 : STD_LOGIC;
  SIGNAL mux_tmp_435 : STD_LOGIC;
  SIGNAL mux_tmp_436 : STD_LOGIC;
  SIGNAL mux_tmp_437 : STD_LOGIC;
  SIGNAL mux_tmp_438 : STD_LOGIC;
  SIGNAL main_stage_0_11 : STD_LOGIC;
  SIGNAL asn_itm_10 : STD_LOGIC;
  SIGNAL result_rem_11cyc_st_9 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_8 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_7 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_6 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_5 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_4 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_3 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_2 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_11 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL asn_itm_11 : STD_LOGIC;
  SIGNAL main_stage_0_12 : STD_LOGIC;
  SIGNAL main_stage_0_3 : STD_LOGIC;
  SIGNAL asn_itm_2 : STD_LOGIC;
  SIGNAL main_stage_0_4 : STD_LOGIC;
  SIGNAL asn_itm_3 : STD_LOGIC;
  SIGNAL main_stage_0_5 : STD_LOGIC;
  SIGNAL asn_itm_4 : STD_LOGIC;
  SIGNAL main_stage_0_6 : STD_LOGIC;
  SIGNAL asn_itm_5 : STD_LOGIC;
  SIGNAL main_stage_0_7 : STD_LOGIC;
  SIGNAL asn_itm_6 : STD_LOGIC;
  SIGNAL main_stage_0_8 : STD_LOGIC;
  SIGNAL asn_itm_7 : STD_LOGIC;
  SIGNAL main_stage_0_9 : STD_LOGIC;
  SIGNAL asn_itm_8 : STD_LOGIC;
  SIGNAL main_stage_0_10 : STD_LOGIC;
  SIGNAL asn_itm_9 : STD_LOGIC;
  SIGNAL main_stage_0_2 : STD_LOGIC;
  SIGNAL asn_itm_1 : STD_LOGIC;
  SIGNAL result_and_1_cse : STD_LOGIC;
  SIGNAL result_and_3_cse : STD_LOGIC;
  SIGNAL result_and_5_cse : STD_LOGIC;
  SIGNAL result_and_7_cse : STD_LOGIC;
  SIGNAL result_and_9_cse : STD_LOGIC;
  SIGNAL result_and_11_cse : STD_LOGIC;
  SIGNAL result_and_13_cse : STD_LOGIC;
  SIGNAL result_and_15_cse : STD_LOGIC;
  SIGNAL result_and_17_cse : STD_LOGIC;
  SIGNAL result_and_19_cse : STD_LOGIC;
  SIGNAL result_and_21_cse : STD_LOGIC;
  SIGNAL or_3_cse : STD_LOGIC;
  SIGNAL or_8_cse : STD_LOGIC;
  SIGNAL or_15_cse : STD_LOGIC;
  SIGNAL or_24_cse : STD_LOGIC;
  SIGNAL or_35_cse : STD_LOGIC;
  SIGNAL or_48_cse : STD_LOGIC;
  SIGNAL or_63_cse : STD_LOGIC;
  SIGNAL or_107_cse : STD_LOGIC;
  SIGNAL or_112_cse : STD_LOGIC;
  SIGNAL or_119_cse : STD_LOGIC;
  SIGNAL or_128_cse : STD_LOGIC;
  SIGNAL or_139_cse : STD_LOGIC;
  SIGNAL or_152_cse : STD_LOGIC;
  SIGNAL or_167_cse : STD_LOGIC;
  SIGNAL or_209_cse : STD_LOGIC;
  SIGNAL or_214_cse : STD_LOGIC;
  SIGNAL or_221_cse : STD_LOGIC;
  SIGNAL or_230_cse : STD_LOGIC;
  SIGNAL or_241_cse : STD_LOGIC;
  SIGNAL or_254_cse : STD_LOGIC;
  SIGNAL or_269_cse : STD_LOGIC;
  SIGNAL or_311_cse : STD_LOGIC;
  SIGNAL or_316_cse : STD_LOGIC;
  SIGNAL or_323_cse : STD_LOGIC;
  SIGNAL or_332_cse : STD_LOGIC;
  SIGNAL or_343_cse : STD_LOGIC;
  SIGNAL or_356_cse : STD_LOGIC;
  SIGNAL or_371_cse : STD_LOGIC;
  SIGNAL nand_144_cse : STD_LOGIC;
  SIGNAL or_413_cse : STD_LOGIC;
  SIGNAL or_418_cse : STD_LOGIC;
  SIGNAL or_425_cse : STD_LOGIC;
  SIGNAL or_434_cse : STD_LOGIC;
  SIGNAL or_445_cse : STD_LOGIC;
  SIGNAL or_458_cse : STD_LOGIC;
  SIGNAL or_473_cse : STD_LOGIC;
  SIGNAL nand_138_cse : STD_LOGIC;
  SIGNAL or_516_cse : STD_LOGIC;
  SIGNAL or_521_cse : STD_LOGIC;
  SIGNAL or_528_cse : STD_LOGIC;
  SIGNAL or_537_cse : STD_LOGIC;
  SIGNAL and_790_cse : STD_LOGIC;
  SIGNAL or_548_cse : STD_LOGIC;
  SIGNAL or_561_cse : STD_LOGIC;
  SIGNAL or_576_cse : STD_LOGIC;
  SIGNAL nand_146_cse : STD_LOGIC;
  SIGNAL or_617_cse : STD_LOGIC;
  SIGNAL or_622_cse : STD_LOGIC;
  SIGNAL or_629_cse : STD_LOGIC;
  SIGNAL or_638_cse : STD_LOGIC;
  SIGNAL or_649_cse : STD_LOGIC;
  SIGNAL or_662_cse : STD_LOGIC;
  SIGNAL or_677_cse : STD_LOGIC;
  SIGNAL or_718_cse : STD_LOGIC;
  SIGNAL nand_112_cse : STD_LOGIC;
  SIGNAL nand_108_cse : STD_LOGIC;
  SIGNAL nand_103_cse : STD_LOGIC;
  SIGNAL nand_97_cse : STD_LOGIC;
  SIGNAL or_763_cse : STD_LOGIC;
  SIGNAL nand_83_cse : STD_LOGIC;
  SIGNAL or_818_cse : STD_LOGIC;
  SIGNAL or_823_cse : STD_LOGIC;
  SIGNAL or_830_cse : STD_LOGIC;
  SIGNAL or_839_cse : STD_LOGIC;
  SIGNAL nand_58_cse : STD_LOGIC;
  SIGNAL or_850_cse : STD_LOGIC;
  SIGNAL nand_55_cse : STD_LOGIC;
  SIGNAL or_863_cse : STD_LOGIC;
  SIGNAL nand_51_cse : STD_LOGIC;
  SIGNAL or_878_cse : STD_LOGIC;
  SIGNAL and_749_cse : STD_LOGIC;
  SIGNAL or_928_cse : STD_LOGIC;
  SIGNAL and_747_cse : STD_LOGIC;
  SIGNAL or_933_cse : STD_LOGIC;
  SIGNAL and_744_cse : STD_LOGIC;
  SIGNAL or_940_cse : STD_LOGIC;
  SIGNAL and_740_cse : STD_LOGIC;
  SIGNAL or_949_cse : STD_LOGIC;
  SIGNAL or_960_cse : STD_LOGIC;
  SIGNAL and_731_cse : STD_LOGIC;
  SIGNAL or_973_cse : STD_LOGIC;
  SIGNAL and_725_cse : STD_LOGIC;
  SIGNAL nand_42_cse : STD_LOGIC;
  SIGNAL or_988_cse : STD_LOGIC;
  SIGNAL or_1037_cse : STD_LOGIC;
  SIGNAL or_1042_cse : STD_LOGIC;
  SIGNAL or_1049_cse : STD_LOGIC;
  SIGNAL or_1058_cse : STD_LOGIC;
  SIGNAL or_1069_cse : STD_LOGIC;
  SIGNAL or_1082_cse : STD_LOGIC;
  SIGNAL or_1097_cse : STD_LOGIC;
  SIGNAL base_buf_sva_mut_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_1_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_1_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_2_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_2_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_3_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_3_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_4_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_4_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_5_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_5_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_6_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_6_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_7_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_7_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_8_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_8_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_9_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_9_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_buf_sva_mut_10_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_mut_10_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_11cyc_st_10 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL return_rsci_d_mx0c0 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c1 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c2 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c3 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c4 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c5 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c6 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c7 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c8 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c9 : STD_LOGIC;
  SIGNAL return_rsci_d_mx0c10 : STD_LOGIC;
  SIGNAL result_acc_imod_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL result_acc_idiv_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL m_and_cse : STD_LOGIC;
  SIGNAL m_and_1_cse : STD_LOGIC;
  SIGNAL m_and_2_cse : STD_LOGIC;
  SIGNAL m_and_3_cse : STD_LOGIC;
  SIGNAL m_and_4_cse : STD_LOGIC;
  SIGNAL m_and_5_cse : STD_LOGIC;
  SIGNAL m_and_6_cse : STD_LOGIC;
  SIGNAL m_and_7_cse : STD_LOGIC;
  SIGNAL m_and_8_cse : STD_LOGIC;
  SIGNAL m_and_9_cse : STD_LOGIC;
  SIGNAL m_and_10_cse : STD_LOGIC;
  SIGNAL m_and_11_cse : STD_LOGIC;
  SIGNAL m_and_12_cse : STD_LOGIC;
  SIGNAL m_and_13_cse : STD_LOGIC;
  SIGNAL m_and_14_cse : STD_LOGIC;
  SIGNAL m_and_15_cse : STD_LOGIC;
  SIGNAL m_and_16_cse : STD_LOGIC;
  SIGNAL m_and_17_cse : STD_LOGIC;
  SIGNAL m_and_18_cse : STD_LOGIC;
  SIGNAL m_and_19_cse : STD_LOGIC;
  SIGNAL m_and_20_cse : STD_LOGIC;
  SIGNAL m_and_21_cse : STD_LOGIC;
  SIGNAL m_and_22_cse : STD_LOGIC;
  SIGNAL m_and_23_cse : STD_LOGIC;
  SIGNAL m_and_24_cse : STD_LOGIC;
  SIGNAL m_and_25_cse : STD_LOGIC;
  SIGNAL m_and_26_cse : STD_LOGIC;
  SIGNAL m_and_27_cse : STD_LOGIC;
  SIGNAL m_and_28_cse : STD_LOGIC;
  SIGNAL m_and_29_cse : STD_LOGIC;
  SIGNAL m_and_30_cse : STD_LOGIC;
  SIGNAL m_and_31_cse : STD_LOGIC;
  SIGNAL m_and_32_cse : STD_LOGIC;
  SIGNAL m_and_33_cse : STD_LOGIC;
  SIGNAL m_and_34_cse : STD_LOGIC;
  SIGNAL m_and_35_cse : STD_LOGIC;
  SIGNAL m_and_36_cse : STD_LOGIC;
  SIGNAL m_and_37_cse : STD_LOGIC;
  SIGNAL m_and_38_cse : STD_LOGIC;
  SIGNAL m_and_39_cse : STD_LOGIC;
  SIGNAL m_and_40_cse : STD_LOGIC;
  SIGNAL m_and_41_cse : STD_LOGIC;
  SIGNAL m_and_42_cse : STD_LOGIC;
  SIGNAL m_and_43_cse : STD_LOGIC;
  SIGNAL m_and_44_cse : STD_LOGIC;
  SIGNAL m_and_45_cse : STD_LOGIC;
  SIGNAL m_and_46_cse : STD_LOGIC;
  SIGNAL m_and_47_cse : STD_LOGIC;
  SIGNAL m_and_48_cse : STD_LOGIC;
  SIGNAL m_and_49_cse : STD_LOGIC;
  SIGNAL m_and_50_cse : STD_LOGIC;
  SIGNAL m_and_51_cse : STD_LOGIC;
  SIGNAL m_and_52_cse : STD_LOGIC;
  SIGNAL m_and_53_cse : STD_LOGIC;
  SIGNAL m_and_54_cse : STD_LOGIC;
  SIGNAL m_and_55_cse : STD_LOGIC;
  SIGNAL m_and_56_cse : STD_LOGIC;
  SIGNAL m_and_57_cse : STD_LOGIC;
  SIGNAL m_and_58_cse : STD_LOGIC;
  SIGNAL m_and_59_cse : STD_LOGIC;
  SIGNAL m_and_60_cse : STD_LOGIC;
  SIGNAL m_and_61_cse : STD_LOGIC;
  SIGNAL m_and_62_cse : STD_LOGIC;
  SIGNAL m_and_63_cse : STD_LOGIC;
  SIGNAL m_and_64_cse : STD_LOGIC;
  SIGNAL m_and_65_cse : STD_LOGIC;
  SIGNAL m_and_66_cse : STD_LOGIC;
  SIGNAL m_and_67_cse : STD_LOGIC;
  SIGNAL m_and_68_cse : STD_LOGIC;
  SIGNAL m_and_69_cse : STD_LOGIC;
  SIGNAL m_and_70_cse : STD_LOGIC;
  SIGNAL m_and_71_cse : STD_LOGIC;
  SIGNAL m_and_72_cse : STD_LOGIC;
  SIGNAL m_and_73_cse : STD_LOGIC;
  SIGNAL m_and_74_cse : STD_LOGIC;
  SIGNAL m_and_75_cse : STD_LOGIC;
  SIGNAL m_and_76_cse : STD_LOGIC;
  SIGNAL m_and_77_cse : STD_LOGIC;
  SIGNAL m_and_78_cse : STD_LOGIC;
  SIGNAL m_and_79_cse : STD_LOGIC;
  SIGNAL m_and_80_cse : STD_LOGIC;
  SIGNAL m_and_81_cse : STD_LOGIC;
  SIGNAL m_and_82_cse : STD_LOGIC;
  SIGNAL m_and_83_cse : STD_LOGIC;
  SIGNAL m_and_84_cse : STD_LOGIC;
  SIGNAL m_and_85_cse : STD_LOGIC;
  SIGNAL m_and_86_cse : STD_LOGIC;
  SIGNAL m_and_87_cse : STD_LOGIC;
  SIGNAL m_and_88_cse : STD_LOGIC;
  SIGNAL m_and_89_cse : STD_LOGIC;
  SIGNAL m_and_90_cse : STD_LOGIC;
  SIGNAL m_and_91_cse : STD_LOGIC;
  SIGNAL m_and_92_cse : STD_LOGIC;
  SIGNAL m_and_93_cse : STD_LOGIC;
  SIGNAL m_and_94_cse : STD_LOGIC;
  SIGNAL m_and_95_cse : STD_LOGIC;
  SIGNAL m_and_96_cse : STD_LOGIC;
  SIGNAL m_and_97_cse : STD_LOGIC;
  SIGNAL m_and_98_cse : STD_LOGIC;

  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL nor_691_nl : STD_LOGIC;
  SIGNAL nor_690_nl : STD_LOGIC;
  SIGNAL or_10_nl : STD_LOGIC;
  SIGNAL mux_2_nl : STD_LOGIC;
  SIGNAL nor_689_nl : STD_LOGIC;
  SIGNAL nor_687_nl : STD_LOGIC;
  SIGNAL or_17_nl : STD_LOGIC;
  SIGNAL nor_688_nl : STD_LOGIC;
  SIGNAL mux_5_nl : STD_LOGIC;
  SIGNAL nor_686_nl : STD_LOGIC;
  SIGNAL nor_683_nl : STD_LOGIC;
  SIGNAL or_26_nl : STD_LOGIC;
  SIGNAL nor_684_nl : STD_LOGIC;
  SIGNAL nor_685_nl : STD_LOGIC;
  SIGNAL mux_9_nl : STD_LOGIC;
  SIGNAL nor_682_nl : STD_LOGIC;
  SIGNAL nor_678_nl : STD_LOGIC;
  SIGNAL or_37_nl : STD_LOGIC;
  SIGNAL nor_679_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL mux_14_nl : STD_LOGIC;
  SIGNAL nor_677_nl : STD_LOGIC;
  SIGNAL nor_672_nl : STD_LOGIC;
  SIGNAL or_50_nl : STD_LOGIC;
  SIGNAL nor_673_nl : STD_LOGIC;
  SIGNAL nor_674_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL nor_676_nl : STD_LOGIC;
  SIGNAL mux_20_nl : STD_LOGIC;
  SIGNAL nor_671_nl : STD_LOGIC;
  SIGNAL nor_665_nl : STD_LOGIC;
  SIGNAL or_65_nl : STD_LOGIC;
  SIGNAL nor_666_nl : STD_LOGIC;
  SIGNAL nor_667_nl : STD_LOGIC;
  SIGNAL nor_668_nl : STD_LOGIC;
  SIGNAL nor_669_nl : STD_LOGIC;
  SIGNAL nor_670_nl : STD_LOGIC;
  SIGNAL mux_27_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL nor_656_nl : STD_LOGIC;
  SIGNAL or_82_nl : STD_LOGIC;
  SIGNAL or_80_nl : STD_LOGIC;
  SIGNAL nor_657_nl : STD_LOGIC;
  SIGNAL nor_658_nl : STD_LOGIC;
  SIGNAL nor_659_nl : STD_LOGIC;
  SIGNAL nor_660_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL nor_662_nl : STD_LOGIC;
  SIGNAL mux_35_nl : STD_LOGIC;
  SIGNAL nor_663_nl : STD_LOGIC;
  SIGNAL nor_654_nl : STD_LOGIC;
  SIGNAL nor_655_nl : STD_LOGIC;
  SIGNAL mux_38_nl : STD_LOGIC;
  SIGNAL nor_653_nl : STD_LOGIC;
  SIGNAL nor_652_nl : STD_LOGIC;
  SIGNAL or_114_nl : STD_LOGIC;
  SIGNAL mux_40_nl : STD_LOGIC;
  SIGNAL nor_651_nl : STD_LOGIC;
  SIGNAL nor_649_nl : STD_LOGIC;
  SIGNAL or_121_nl : STD_LOGIC;
  SIGNAL nor_650_nl : STD_LOGIC;
  SIGNAL mux_43_nl : STD_LOGIC;
  SIGNAL nor_648_nl : STD_LOGIC;
  SIGNAL nor_645_nl : STD_LOGIC;
  SIGNAL or_130_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL nor_647_nl : STD_LOGIC;
  SIGNAL mux_47_nl : STD_LOGIC;
  SIGNAL nor_644_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL or_141_nl : STD_LOGIC;
  SIGNAL nor_641_nl : STD_LOGIC;
  SIGNAL nor_642_nl : STD_LOGIC;
  SIGNAL nor_643_nl : STD_LOGIC;
  SIGNAL mux_52_nl : STD_LOGIC;
  SIGNAL nor_639_nl : STD_LOGIC;
  SIGNAL nor_634_nl : STD_LOGIC;
  SIGNAL or_154_nl : STD_LOGIC;
  SIGNAL nor_635_nl : STD_LOGIC;
  SIGNAL nor_636_nl : STD_LOGIC;
  SIGNAL nor_637_nl : STD_LOGIC;
  SIGNAL nor_638_nl : STD_LOGIC;
  SIGNAL mux_58_nl : STD_LOGIC;
  SIGNAL nor_633_nl : STD_LOGIC;
  SIGNAL nor_627_nl : STD_LOGIC;
  SIGNAL or_169_nl : STD_LOGIC;
  SIGNAL nor_628_nl : STD_LOGIC;
  SIGNAL nor_629_nl : STD_LOGIC;
  SIGNAL nor_630_nl : STD_LOGIC;
  SIGNAL nor_631_nl : STD_LOGIC;
  SIGNAL nor_632_nl : STD_LOGIC;
  SIGNAL mux_65_nl : STD_LOGIC;
  SIGNAL nor_626_nl : STD_LOGIC;
  SIGNAL nor_618_nl : STD_LOGIC;
  SIGNAL or_186_nl : STD_LOGIC;
  SIGNAL or_184_nl : STD_LOGIC;
  SIGNAL nor_619_nl : STD_LOGIC;
  SIGNAL nor_620_nl : STD_LOGIC;
  SIGNAL nor_621_nl : STD_LOGIC;
  SIGNAL nor_622_nl : STD_LOGIC;
  SIGNAL nor_623_nl : STD_LOGIC;
  SIGNAL nor_624_nl : STD_LOGIC;
  SIGNAL mux_73_nl : STD_LOGIC;
  SIGNAL nor_625_nl : STD_LOGIC;
  SIGNAL nor_617_nl : STD_LOGIC;
  SIGNAL and_797_nl : STD_LOGIC;
  SIGNAL or_195_nl : STD_LOGIC;
  SIGNAL mux_76_nl : STD_LOGIC;
  SIGNAL nor_616_nl : STD_LOGIC;
  SIGNAL nor_615_nl : STD_LOGIC;
  SIGNAL or_216_nl : STD_LOGIC;
  SIGNAL mux_78_nl : STD_LOGIC;
  SIGNAL nor_614_nl : STD_LOGIC;
  SIGNAL nor_612_nl : STD_LOGIC;
  SIGNAL or_223_nl : STD_LOGIC;
  SIGNAL nor_613_nl : STD_LOGIC;
  SIGNAL mux_81_nl : STD_LOGIC;
  SIGNAL nor_611_nl : STD_LOGIC;
  SIGNAL nor_608_nl : STD_LOGIC;
  SIGNAL or_232_nl : STD_LOGIC;
  SIGNAL nor_609_nl : STD_LOGIC;
  SIGNAL nor_610_nl : STD_LOGIC;
  SIGNAL mux_85_nl : STD_LOGIC;
  SIGNAL nor_607_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL or_243_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL nor_605_nl : STD_LOGIC;
  SIGNAL nor_606_nl : STD_LOGIC;
  SIGNAL mux_90_nl : STD_LOGIC;
  SIGNAL nor_602_nl : STD_LOGIC;
  SIGNAL nor_597_nl : STD_LOGIC;
  SIGNAL or_256_nl : STD_LOGIC;
  SIGNAL nor_598_nl : STD_LOGIC;
  SIGNAL nor_599_nl : STD_LOGIC;
  SIGNAL nor_600_nl : STD_LOGIC;
  SIGNAL nor_601_nl : STD_LOGIC;
  SIGNAL mux_96_nl : STD_LOGIC;
  SIGNAL nor_596_nl : STD_LOGIC;
  SIGNAL nor_590_nl : STD_LOGIC;
  SIGNAL or_271_nl : STD_LOGIC;
  SIGNAL nor_591_nl : STD_LOGIC;
  SIGNAL nor_592_nl : STD_LOGIC;
  SIGNAL nor_593_nl : STD_LOGIC;
  SIGNAL nor_594_nl : STD_LOGIC;
  SIGNAL nor_595_nl : STD_LOGIC;
  SIGNAL mux_103_nl : STD_LOGIC;
  SIGNAL nor_589_nl : STD_LOGIC;
  SIGNAL nor_581_nl : STD_LOGIC;
  SIGNAL or_288_nl : STD_LOGIC;
  SIGNAL or_286_nl : STD_LOGIC;
  SIGNAL nor_582_nl : STD_LOGIC;
  SIGNAL nor_583_nl : STD_LOGIC;
  SIGNAL nor_584_nl : STD_LOGIC;
  SIGNAL nor_585_nl : STD_LOGIC;
  SIGNAL nor_586_nl : STD_LOGIC;
  SIGNAL nor_587_nl : STD_LOGIC;
  SIGNAL mux_111_nl : STD_LOGIC;
  SIGNAL nor_588_nl : STD_LOGIC;
  SIGNAL nor_579_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL mux_114_nl : STD_LOGIC;
  SIGNAL nor_578_nl : STD_LOGIC;
  SIGNAL nor_577_nl : STD_LOGIC;
  SIGNAL or_318_nl : STD_LOGIC;
  SIGNAL mux_116_nl : STD_LOGIC;
  SIGNAL nor_576_nl : STD_LOGIC;
  SIGNAL nor_574_nl : STD_LOGIC;
  SIGNAL or_325_nl : STD_LOGIC;
  SIGNAL nor_575_nl : STD_LOGIC;
  SIGNAL mux_119_nl : STD_LOGIC;
  SIGNAL nor_573_nl : STD_LOGIC;
  SIGNAL nor_570_nl : STD_LOGIC;
  SIGNAL or_334_nl : STD_LOGIC;
  SIGNAL nor_571_nl : STD_LOGIC;
  SIGNAL nor_572_nl : STD_LOGIC;
  SIGNAL mux_123_nl : STD_LOGIC;
  SIGNAL nor_569_nl : STD_LOGIC;
  SIGNAL nor_565_nl : STD_LOGIC;
  SIGNAL or_345_nl : STD_LOGIC;
  SIGNAL nor_566_nl : STD_LOGIC;
  SIGNAL nor_567_nl : STD_LOGIC;
  SIGNAL nor_568_nl : STD_LOGIC;
  SIGNAL mux_128_nl : STD_LOGIC;
  SIGNAL nor_564_nl : STD_LOGIC;
  SIGNAL nor_559_nl : STD_LOGIC;
  SIGNAL or_358_nl : STD_LOGIC;
  SIGNAL nor_560_nl : STD_LOGIC;
  SIGNAL nor_561_nl : STD_LOGIC;
  SIGNAL nor_562_nl : STD_LOGIC;
  SIGNAL nor_563_nl : STD_LOGIC;
  SIGNAL mux_134_nl : STD_LOGIC;
  SIGNAL nor_558_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL or_373_nl : STD_LOGIC;
  SIGNAL nor_553_nl : STD_LOGIC;
  SIGNAL nor_554_nl : STD_LOGIC;
  SIGNAL nor_555_nl : STD_LOGIC;
  SIGNAL nor_556_nl : STD_LOGIC;
  SIGNAL nor_557_nl : STD_LOGIC;
  SIGNAL mux_141_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL nor_543_nl : STD_LOGIC;
  SIGNAL or_390_nl : STD_LOGIC;
  SIGNAL or_388_nl : STD_LOGIC;
  SIGNAL nor_544_nl : STD_LOGIC;
  SIGNAL nor_545_nl : STD_LOGIC;
  SIGNAL nor_546_nl : STD_LOGIC;
  SIGNAL nor_547_nl : STD_LOGIC;
  SIGNAL nor_548_nl : STD_LOGIC;
  SIGNAL nor_549_nl : STD_LOGIC;
  SIGNAL mux_149_nl : STD_LOGIC;
  SIGNAL nor_550_nl : STD_LOGIC;
  SIGNAL nor_542_nl : STD_LOGIC;
  SIGNAL and_796_nl : STD_LOGIC;
  SIGNAL or_399_nl : STD_LOGIC;
  SIGNAL mux_152_nl : STD_LOGIC;
  SIGNAL and_795_nl : STD_LOGIC;
  SIGNAL nor_541_nl : STD_LOGIC;
  SIGNAL or_420_nl : STD_LOGIC;
  SIGNAL mux_154_nl : STD_LOGIC;
  SIGNAL and_794_nl : STD_LOGIC;
  SIGNAL nor_539_nl : STD_LOGIC;
  SIGNAL or_427_nl : STD_LOGIC;
  SIGNAL nor_540_nl : STD_LOGIC;
  SIGNAL mux_157_nl : STD_LOGIC;
  SIGNAL and_793_nl : STD_LOGIC;
  SIGNAL nor_536_nl : STD_LOGIC;
  SIGNAL or_436_nl : STD_LOGIC;
  SIGNAL nor_537_nl : STD_LOGIC;
  SIGNAL nor_538_nl : STD_LOGIC;
  SIGNAL mux_161_nl : STD_LOGIC;
  SIGNAL and_792_nl : STD_LOGIC;
  SIGNAL nor_532_nl : STD_LOGIC;
  SIGNAL or_447_nl : STD_LOGIC;
  SIGNAL nor_533_nl : STD_LOGIC;
  SIGNAL nor_534_nl : STD_LOGIC;
  SIGNAL nor_535_nl : STD_LOGIC;
  SIGNAL mux_166_nl : STD_LOGIC;
  SIGNAL and_791_nl : STD_LOGIC;
  SIGNAL nor_527_nl : STD_LOGIC;
  SIGNAL or_460_nl : STD_LOGIC;
  SIGNAL nor_528_nl : STD_LOGIC;
  SIGNAL nor_529_nl : STD_LOGIC;
  SIGNAL nor_530_nl : STD_LOGIC;
  SIGNAL nor_531_nl : STD_LOGIC;
  SIGNAL mux_172_nl : STD_LOGIC;
  SIGNAL and_789_nl : STD_LOGIC;
  SIGNAL nor_522_nl : STD_LOGIC;
  SIGNAL or_475_nl : STD_LOGIC;
  SIGNAL and_788_nl : STD_LOGIC;
  SIGNAL nor_523_nl : STD_LOGIC;
  SIGNAL nor_524_nl : STD_LOGIC;
  SIGNAL nor_525_nl : STD_LOGIC;
  SIGNAL nor_526_nl : STD_LOGIC;
  SIGNAL mux_179_nl : STD_LOGIC;
  SIGNAL and_787_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL or_492_nl : STD_LOGIC;
  SIGNAL or_490_nl : STD_LOGIC;
  SIGNAL nor_517_nl : STD_LOGIC;
  SIGNAL and_785_nl : STD_LOGIC;
  SIGNAL nor_518_nl : STD_LOGIC;
  SIGNAL nor_519_nl : STD_LOGIC;
  SIGNAL nor_520_nl : STD_LOGIC;
  SIGNAL nor_521_nl : STD_LOGIC;
  SIGNAL mux_187_nl : STD_LOGIC;
  SIGNAL and_786_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL or_501_nl : STD_LOGIC;
  SIGNAL mux_190_nl : STD_LOGIC;
  SIGNAL and_784_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL or_523_nl : STD_LOGIC;
  SIGNAL mux_192_nl : STD_LOGIC;
  SIGNAL and_783_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL or_530_nl : STD_LOGIC;
  SIGNAL nor_512_nl : STD_LOGIC;
  SIGNAL mux_195_nl : STD_LOGIC;
  SIGNAL and_782_nl : STD_LOGIC;
  SIGNAL nor_508_nl : STD_LOGIC;
  SIGNAL or_539_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL mux_199_nl : STD_LOGIC;
  SIGNAL and_781_nl : STD_LOGIC;
  SIGNAL nor_504_nl : STD_LOGIC;
  SIGNAL or_550_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL nor_506_nl : STD_LOGIC;
  SIGNAL nor_507_nl : STD_LOGIC;
  SIGNAL mux_204_nl : STD_LOGIC;
  SIGNAL and_780_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL or_563_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL nor_501_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL nor_503_nl : STD_LOGIC;
  SIGNAL mux_210_nl : STD_LOGIC;
  SIGNAL and_778_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL or_578_nl : STD_LOGIC;
  SIGNAL and_777_nl : STD_LOGIC;
  SIGNAL nor_495_nl : STD_LOGIC;
  SIGNAL nor_496_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL mux_217_nl : STD_LOGIC;
  SIGNAL and_776_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL or_595_nl : STD_LOGIC;
  SIGNAL or_593_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL and_774_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL nor_491_nl : STD_LOGIC;
  SIGNAL nor_492_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL mux_225_nl : STD_LOGIC;
  SIGNAL and_775_nl : STD_LOGIC;
  SIGNAL nor_487_nl : STD_LOGIC;
  SIGNAL and_773_nl : STD_LOGIC;
  SIGNAL or_604_nl : STD_LOGIC;
  SIGNAL mux_228_nl : STD_LOGIC;
  SIGNAL and_772_nl : STD_LOGIC;
  SIGNAL nor_486_nl : STD_LOGIC;
  SIGNAL or_624_nl : STD_LOGIC;
  SIGNAL mux_230_nl : STD_LOGIC;
  SIGNAL and_771_nl : STD_LOGIC;
  SIGNAL nor_484_nl : STD_LOGIC;
  SIGNAL or_631_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL mux_233_nl : STD_LOGIC;
  SIGNAL and_770_nl : STD_LOGIC;
  SIGNAL nor_481_nl : STD_LOGIC;
  SIGNAL or_640_nl : STD_LOGIC;
  SIGNAL nor_482_nl : STD_LOGIC;
  SIGNAL nor_483_nl : STD_LOGIC;
  SIGNAL mux_237_nl : STD_LOGIC;
  SIGNAL and_769_nl : STD_LOGIC;
  SIGNAL nor_477_nl : STD_LOGIC;
  SIGNAL or_651_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL nor_479_nl : STD_LOGIC;
  SIGNAL nor_480_nl : STD_LOGIC;
  SIGNAL mux_242_nl : STD_LOGIC;
  SIGNAL and_768_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL or_664_nl : STD_LOGIC;
  SIGNAL nor_473_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL nor_476_nl : STD_LOGIC;
  SIGNAL mux_248_nl : STD_LOGIC;
  SIGNAL and_766_nl : STD_LOGIC;
  SIGNAL nor_467_nl : STD_LOGIC;
  SIGNAL or_679_nl : STD_LOGIC;
  SIGNAL and_765_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL nor_471_nl : STD_LOGIC;
  SIGNAL mux_255_nl : STD_LOGIC;
  SIGNAL and_764_nl : STD_LOGIC;
  SIGNAL nor_461_nl : STD_LOGIC;
  SIGNAL or_696_nl : STD_LOGIC;
  SIGNAL or_694_nl : STD_LOGIC;
  SIGNAL nor_462_nl : STD_LOGIC;
  SIGNAL and_762_nl : STD_LOGIC;
  SIGNAL nor_463_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL nor_465_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL mux_263_nl : STD_LOGIC;
  SIGNAL and_763_nl : STD_LOGIC;
  SIGNAL nor_459_nl : STD_LOGIC;
  SIGNAL nor_460_nl : STD_LOGIC;
  SIGNAL or_705_nl : STD_LOGIC;
  SIGNAL mux_266_nl : STD_LOGIC;
  SIGNAL and_761_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL nand_153_nl : STD_LOGIC;
  SIGNAL mux_268_nl : STD_LOGIC;
  SIGNAL and_760_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL nand_152_nl : STD_LOGIC;
  SIGNAL nor_457_nl : STD_LOGIC;
  SIGNAL mux_271_nl : STD_LOGIC;
  SIGNAL and_759_nl : STD_LOGIC;
  SIGNAL nor_453_nl : STD_LOGIC;
  SIGNAL nand_151_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL mux_275_nl : STD_LOGIC;
  SIGNAL and_758_nl : STD_LOGIC;
  SIGNAL nor_449_nl : STD_LOGIC;
  SIGNAL nand_96_nl : STD_LOGIC;
  SIGNAL nor_450_nl : STD_LOGIC;
  SIGNAL nor_451_nl : STD_LOGIC;
  SIGNAL nor_452_nl : STD_LOGIC;
  SIGNAL mux_280_nl : STD_LOGIC;
  SIGNAL and_757_nl : STD_LOGIC;
  SIGNAL nor_444_nl : STD_LOGIC;
  SIGNAL nand_150_nl : STD_LOGIC;
  SIGNAL nor_445_nl : STD_LOGIC;
  SIGNAL nor_446_nl : STD_LOGIC;
  SIGNAL nor_447_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL mux_286_nl : STD_LOGIC;
  SIGNAL and_755_nl : STD_LOGIC;
  SIGNAL nor_439_nl : STD_LOGIC;
  SIGNAL nand_149_nl : STD_LOGIC;
  SIGNAL and_754_nl : STD_LOGIC;
  SIGNAL nor_440_nl : STD_LOGIC;
  SIGNAL nor_441_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL nor_443_nl : STD_LOGIC;
  SIGNAL mux_293_nl : STD_LOGIC;
  SIGNAL and_753_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL nand_72_nl : STD_LOGIC;
  SIGNAL nand_73_nl : STD_LOGIC;
  SIGNAL nor_434_nl : STD_LOGIC;
  SIGNAL and_751_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL nor_436_nl : STD_LOGIC;
  SIGNAL nor_437_nl : STD_LOGIC;
  SIGNAL nor_438_nl : STD_LOGIC;
  SIGNAL mux_301_nl : STD_LOGIC;
  SIGNAL and_752_nl : STD_LOGIC;
  SIGNAL nor_432_nl : STD_LOGIC;
  SIGNAL and_750_nl : STD_LOGIC;
  SIGNAL mux_304_nl : STD_LOGIC;
  SIGNAL nor_431_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL or_825_nl : STD_LOGIC;
  SIGNAL mux_306_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL nor_428_nl : STD_LOGIC;
  SIGNAL or_832_nl : STD_LOGIC;
  SIGNAL and_748_nl : STD_LOGIC;
  SIGNAL mux_309_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL nor_426_nl : STD_LOGIC;
  SIGNAL or_841_nl : STD_LOGIC;
  SIGNAL and_745_nl : STD_LOGIC;
  SIGNAL and_746_nl : STD_LOGIC;
  SIGNAL mux_313_nl : STD_LOGIC;
  SIGNAL nor_425_nl : STD_LOGIC;
  SIGNAL nor_424_nl : STD_LOGIC;
  SIGNAL or_852_nl : STD_LOGIC;
  SIGNAL and_741_nl : STD_LOGIC;
  SIGNAL and_742_nl : STD_LOGIC;
  SIGNAL and_743_nl : STD_LOGIC;
  SIGNAL mux_318_nl : STD_LOGIC;
  SIGNAL nor_423_nl : STD_LOGIC;
  SIGNAL nor_422_nl : STD_LOGIC;
  SIGNAL or_865_nl : STD_LOGIC;
  SIGNAL and_736_nl : STD_LOGIC;
  SIGNAL and_737_nl : STD_LOGIC;
  SIGNAL and_738_nl : STD_LOGIC;
  SIGNAL and_739_nl : STD_LOGIC;
  SIGNAL mux_324_nl : STD_LOGIC;
  SIGNAL nor_421_nl : STD_LOGIC;
  SIGNAL nor_419_nl : STD_LOGIC;
  SIGNAL or_880_nl : STD_LOGIC;
  SIGNAL nor_420_nl : STD_LOGIC;
  SIGNAL and_732_nl : STD_LOGIC;
  SIGNAL and_733_nl : STD_LOGIC;
  SIGNAL and_734_nl : STD_LOGIC;
  SIGNAL and_735_nl : STD_LOGIC;
  SIGNAL mux_331_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL nor_415_nl : STD_LOGIC;
  SIGNAL or_897_nl : STD_LOGIC;
  SIGNAL or_895_nl : STD_LOGIC;
  SIGNAL and_726_nl : STD_LOGIC;
  SIGNAL nor_416_nl : STD_LOGIC;
  SIGNAL and_727_nl : STD_LOGIC;
  SIGNAL and_728_nl : STD_LOGIC;
  SIGNAL and_729_nl : STD_LOGIC;
  SIGNAL and_730_nl : STD_LOGIC;
  SIGNAL mux_339_nl : STD_LOGIC;
  SIGNAL nor_417_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL or_914_nl : STD_LOGIC;
  SIGNAL nor_408_nl : STD_LOGIC;
  SIGNAL or_913_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL or_912_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL or_911_nl : STD_LOGIC;
  SIGNAL nor_411_nl : STD_LOGIC;
  SIGNAL or_910_nl : STD_LOGIC;
  SIGNAL nor_412_nl : STD_LOGIC;
  SIGNAL or_909_nl : STD_LOGIC;
  SIGNAL nor_413_nl : STD_LOGIC;
  SIGNAL or_908_nl : STD_LOGIC;
  SIGNAL and_724_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL mux_349_nl : STD_LOGIC;
  SIGNAL nor_406_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL or_935_nl : STD_LOGIC;
  SIGNAL mux_351_nl : STD_LOGIC;
  SIGNAL nor_404_nl : STD_LOGIC;
  SIGNAL nor_403_nl : STD_LOGIC;
  SIGNAL or_942_nl : STD_LOGIC;
  SIGNAL and_722_nl : STD_LOGIC;
  SIGNAL mux_354_nl : STD_LOGIC;
  SIGNAL nor_402_nl : STD_LOGIC;
  SIGNAL nor_401_nl : STD_LOGIC;
  SIGNAL or_951_nl : STD_LOGIC;
  SIGNAL and_719_nl : STD_LOGIC;
  SIGNAL and_720_nl : STD_LOGIC;
  SIGNAL mux_358_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL nor_399_nl : STD_LOGIC;
  SIGNAL or_962_nl : STD_LOGIC;
  SIGNAL and_715_nl : STD_LOGIC;
  SIGNAL and_716_nl : STD_LOGIC;
  SIGNAL and_717_nl : STD_LOGIC;
  SIGNAL mux_363_nl : STD_LOGIC;
  SIGNAL nor_398_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL or_975_nl : STD_LOGIC;
  SIGNAL and_710_nl : STD_LOGIC;
  SIGNAL and_711_nl : STD_LOGIC;
  SIGNAL and_712_nl : STD_LOGIC;
  SIGNAL and_713_nl : STD_LOGIC;
  SIGNAL mux_369_nl : STD_LOGIC;
  SIGNAL nor_396_nl : STD_LOGIC;
  SIGNAL nor_394_nl : STD_LOGIC;
  SIGNAL or_990_nl : STD_LOGIC;
  SIGNAL nor_395_nl : STD_LOGIC;
  SIGNAL and_706_nl : STD_LOGIC;
  SIGNAL and_707_nl : STD_LOGIC;
  SIGNAL and_708_nl : STD_LOGIC;
  SIGNAL and_709_nl : STD_LOGIC;
  SIGNAL mux_376_nl : STD_LOGIC;
  SIGNAL nor_393_nl : STD_LOGIC;
  SIGNAL nor_390_nl : STD_LOGIC;
  SIGNAL or_1007_nl : STD_LOGIC;
  SIGNAL or_1005_nl : STD_LOGIC;
  SIGNAL and_700_nl : STD_LOGIC;
  SIGNAL nor_391_nl : STD_LOGIC;
  SIGNAL and_701_nl : STD_LOGIC;
  SIGNAL and_702_nl : STD_LOGIC;
  SIGNAL and_703_nl : STD_LOGIC;
  SIGNAL and_704_nl : STD_LOGIC;
  SIGNAL mux_384_nl : STD_LOGIC;
  SIGNAL nor_392_nl : STD_LOGIC;
  SIGNAL nor_383_nl : STD_LOGIC;
  SIGNAL or_1024_nl : STD_LOGIC;
  SIGNAL nor_384_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL nor_385_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL or_1021_nl : STD_LOGIC;
  SIGNAL nor_387_nl : STD_LOGIC;
  SIGNAL or_1020_nl : STD_LOGIC;
  SIGNAL nor_388_nl : STD_LOGIC;
  SIGNAL or_1019_nl : STD_LOGIC;
  SIGNAL nor_389_nl : STD_LOGIC;
  SIGNAL or_1018_nl : STD_LOGIC;
  SIGNAL and_697_nl : STD_LOGIC;
  SIGNAL and_698_nl : STD_LOGIC;
  SIGNAL or_1016_nl : STD_LOGIC;
  SIGNAL mux_394_nl : STD_LOGIC;
  SIGNAL nor_382_nl : STD_LOGIC;
  SIGNAL nor_381_nl : STD_LOGIC;
  SIGNAL or_1044_nl : STD_LOGIC;
  SIGNAL mux_396_nl : STD_LOGIC;
  SIGNAL nor_380_nl : STD_LOGIC;
  SIGNAL nor_379_nl : STD_LOGIC;
  SIGNAL or_1051_nl : STD_LOGIC;
  SIGNAL and_695_nl : STD_LOGIC;
  SIGNAL mux_399_nl : STD_LOGIC;
  SIGNAL nor_378_nl : STD_LOGIC;
  SIGNAL nor_377_nl : STD_LOGIC;
  SIGNAL or_1060_nl : STD_LOGIC;
  SIGNAL and_692_nl : STD_LOGIC;
  SIGNAL and_693_nl : STD_LOGIC;
  SIGNAL mux_403_nl : STD_LOGIC;
  SIGNAL nor_376_nl : STD_LOGIC;
  SIGNAL nor_375_nl : STD_LOGIC;
  SIGNAL or_1071_nl : STD_LOGIC;
  SIGNAL and_688_nl : STD_LOGIC;
  SIGNAL and_689_nl : STD_LOGIC;
  SIGNAL and_690_nl : STD_LOGIC;
  SIGNAL mux_408_nl : STD_LOGIC;
  SIGNAL nor_374_nl : STD_LOGIC;
  SIGNAL nor_373_nl : STD_LOGIC;
  SIGNAL or_1084_nl : STD_LOGIC;
  SIGNAL and_683_nl : STD_LOGIC;
  SIGNAL and_684_nl : STD_LOGIC;
  SIGNAL and_685_nl : STD_LOGIC;
  SIGNAL and_686_nl : STD_LOGIC;
  SIGNAL mux_414_nl : STD_LOGIC;
  SIGNAL nor_372_nl : STD_LOGIC;
  SIGNAL nor_370_nl : STD_LOGIC;
  SIGNAL or_1099_nl : STD_LOGIC;
  SIGNAL nor_371_nl : STD_LOGIC;
  SIGNAL and_679_nl : STD_LOGIC;
  SIGNAL and_680_nl : STD_LOGIC;
  SIGNAL and_681_nl : STD_LOGIC;
  SIGNAL and_682_nl : STD_LOGIC;
  SIGNAL mux_421_nl : STD_LOGIC;
  SIGNAL nor_369_nl : STD_LOGIC;
  SIGNAL nor_366_nl : STD_LOGIC;
  SIGNAL or_1116_nl : STD_LOGIC;
  SIGNAL or_1114_nl : STD_LOGIC;
  SIGNAL and_673_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL and_674_nl : STD_LOGIC;
  SIGNAL and_675_nl : STD_LOGIC;
  SIGNAL and_676_nl : STD_LOGIC;
  SIGNAL and_677_nl : STD_LOGIC;
  SIGNAL mux_429_nl : STD_LOGIC;
  SIGNAL nor_368_nl : STD_LOGIC;
  SIGNAL nor_358_nl : STD_LOGIC;
  SIGNAL or_1133_nl : STD_LOGIC;
  SIGNAL nor_359_nl : STD_LOGIC;
  SIGNAL or_1132_nl : STD_LOGIC;
  SIGNAL nor_360_nl : STD_LOGIC;
  SIGNAL or_1131_nl : STD_LOGIC;
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL or_1130_nl : STD_LOGIC;
  SIGNAL nor_362_nl : STD_LOGIC;
  SIGNAL or_1129_nl : STD_LOGIC;
  SIGNAL nor_363_nl : STD_LOGIC;
  SIGNAL or_1128_nl : STD_LOGIC;
  SIGNAL nor_364_nl : STD_LOGIC;
  SIGNAL or_1127_nl : STD_LOGIC;
  SIGNAL and_671_nl : STD_LOGIC;
  SIGNAL nor_365_nl : STD_LOGIC;
  SIGNAL base_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL m_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL return_rsci_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL ccs_ccore_start_rsci_dat : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat_1 : STD_LOGIC_VECTOR (0 DOWNTO 0);

  SIGNAL result_rem_12_cmp_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_1_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_1_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_2_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_2_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_3_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_3_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_4_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_4_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_5_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_5_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_6_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_6_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_7_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_7_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_8_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_8_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_9_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_9_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL result_rem_12_cmp_10_a_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_b_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL result_rem_12_cmp_10_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_v_64_10_2(input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(9 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_11_2(input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  base_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 1,
      width => 64
      )
    PORT MAP(
      dat => base_rsci_dat,
      idat => base_rsci_idat_1
    );
  base_rsci_dat <= base_rsc_dat;
  base_rsci_idat <= base_rsci_idat_1;

  m_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => m_rsci_dat,
      idat => m_rsci_idat_1
    );
  m_rsci_dat <= m_rsc_dat;
  m_rsci_idat <= m_rsci_idat_1;

  return_rsci : work.mgc_out_dreg_pkg_v2.mgc_out_dreg_v2
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      d => return_rsci_d_1,
      z => return_rsci_z
    );
  return_rsci_d_1 <= return_rsci_d;
  return_rsc_z <= return_rsci_z;

  ccs_ccore_start_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 8,
      width => 1
      )
    PORT MAP(
      dat => ccs_ccore_start_rsci_dat,
      idat => ccs_ccore_start_rsci_idat_1
    );
  ccs_ccore_start_rsci_dat(0) <= ccs_ccore_start_rsc_dat;
  ccs_ccore_start_rsci_idat <= ccs_ccore_start_rsci_idat_1(0);

  result_rem_12_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_a_1,
      b => result_rem_12_cmp_b_1,
      z => result_rem_12_cmp_z_1
    );
  result_rem_12_cmp_a_1 <= result_rem_12_cmp_a;
  result_rem_12_cmp_b_1 <= result_rem_12_cmp_b;
  result_rem_12_cmp_z <= result_rem_12_cmp_z_1;

  result_rem_12_cmp_1 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_1_a_1,
      b => result_rem_12_cmp_1_b_1,
      z => result_rem_12_cmp_1_z_1
    );
  result_rem_12_cmp_1_a_1 <= result_rem_12_cmp_1_a;
  result_rem_12_cmp_1_b_1 <= result_rem_12_cmp_1_b;
  result_rem_12_cmp_1_z <= result_rem_12_cmp_1_z_1;

  result_rem_12_cmp_2 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_2_a_1,
      b => result_rem_12_cmp_2_b_1,
      z => result_rem_12_cmp_2_z_1
    );
  result_rem_12_cmp_2_a_1 <= result_rem_12_cmp_2_a;
  result_rem_12_cmp_2_b_1 <= result_rem_12_cmp_2_b;
  result_rem_12_cmp_2_z <= result_rem_12_cmp_2_z_1;

  result_rem_12_cmp_3 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_3_a_1,
      b => result_rem_12_cmp_3_b_1,
      z => result_rem_12_cmp_3_z_1
    );
  result_rem_12_cmp_3_a_1 <= result_rem_12_cmp_3_a;
  result_rem_12_cmp_3_b_1 <= result_rem_12_cmp_3_b;
  result_rem_12_cmp_3_z <= result_rem_12_cmp_3_z_1;

  result_rem_12_cmp_4 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_4_a_1,
      b => result_rem_12_cmp_4_b_1,
      z => result_rem_12_cmp_4_z_1
    );
  result_rem_12_cmp_4_a_1 <= result_rem_12_cmp_4_a;
  result_rem_12_cmp_4_b_1 <= result_rem_12_cmp_4_b;
  result_rem_12_cmp_4_z <= result_rem_12_cmp_4_z_1;

  result_rem_12_cmp_5 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_5_a_1,
      b => result_rem_12_cmp_5_b_1,
      z => result_rem_12_cmp_5_z_1
    );
  result_rem_12_cmp_5_a_1 <= result_rem_12_cmp_5_a;
  result_rem_12_cmp_5_b_1 <= result_rem_12_cmp_5_b;
  result_rem_12_cmp_5_z <= result_rem_12_cmp_5_z_1;

  result_rem_12_cmp_6 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_6_a_1,
      b => result_rem_12_cmp_6_b_1,
      z => result_rem_12_cmp_6_z_1
    );
  result_rem_12_cmp_6_a_1 <= result_rem_12_cmp_6_a;
  result_rem_12_cmp_6_b_1 <= result_rem_12_cmp_6_b;
  result_rem_12_cmp_6_z <= result_rem_12_cmp_6_z_1;

  result_rem_12_cmp_7 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_7_a_1,
      b => result_rem_12_cmp_7_b_1,
      z => result_rem_12_cmp_7_z_1
    );
  result_rem_12_cmp_7_a_1 <= result_rem_12_cmp_7_a;
  result_rem_12_cmp_7_b_1 <= result_rem_12_cmp_7_b;
  result_rem_12_cmp_7_z <= result_rem_12_cmp_7_z_1;

  result_rem_12_cmp_8 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_8_a_1,
      b => result_rem_12_cmp_8_b_1,
      z => result_rem_12_cmp_8_z_1
    );
  result_rem_12_cmp_8_a_1 <= result_rem_12_cmp_8_a;
  result_rem_12_cmp_8_b_1 <= result_rem_12_cmp_8_b;
  result_rem_12_cmp_8_z <= result_rem_12_cmp_8_z_1;

  result_rem_12_cmp_9 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_9_a_1,
      b => result_rem_12_cmp_9_b_1,
      z => result_rem_12_cmp_9_z_1
    );
  result_rem_12_cmp_9_a_1 <= result_rem_12_cmp_9_a;
  result_rem_12_cmp_9_b_1 <= result_rem_12_cmp_9_b;
  result_rem_12_cmp_9_z <= result_rem_12_cmp_9_z_1;

  result_rem_12_cmp_10 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 64,
      width_b => 64,
      signd => 0
      )
    PORT MAP(
      a => result_rem_12_cmp_10_a_1,
      b => result_rem_12_cmp_10_b_1,
      z => result_rem_12_cmp_10_z_1
    );
  result_rem_12_cmp_10_a_1 <= result_rem_12_cmp_10_a;
  result_rem_12_cmp_10_b_1 <= result_rem_12_cmp_10_b;
  result_rem_12_cmp_10_z <= result_rem_12_cmp_10_z_1;

  result_and_1_cse <= ccs_ccore_en AND (and_dcpl_263 OR and_dcpl_269 OR and_dcpl_275
      OR and_dcpl_281 OR and_dcpl_287 OR and_dcpl_293 OR and_dcpl_299 OR and_dcpl_305
      OR and_dcpl_311 OR mux_tmp_37);
  result_and_3_cse <= ccs_ccore_en AND (and_dcpl_319 OR and_dcpl_322 OR and_dcpl_325
      OR and_dcpl_329 OR and_dcpl_333 OR and_dcpl_337 OR and_dcpl_341 OR and_dcpl_344
      OR and_dcpl_347 OR mux_tmp_75);
  result_and_5_cse <= ccs_ccore_en AND (and_dcpl_353 OR and_dcpl_357 OR and_dcpl_361
      OR and_dcpl_364 OR and_dcpl_367 OR and_dcpl_370 OR and_dcpl_373 OR and_dcpl_377
      OR and_dcpl_381 OR mux_tmp_113);
  result_and_7_cse <= ccs_ccore_en AND (and_dcpl_387 OR and_dcpl_390 OR and_dcpl_393
      OR and_dcpl_396 OR and_dcpl_399 OR and_dcpl_402 OR and_dcpl_405 OR and_dcpl_408
      OR and_dcpl_411 OR mux_tmp_151);
  result_and_9_cse <= ccs_ccore_en AND (and_dcpl_418 OR and_dcpl_422 OR and_dcpl_426
      OR and_dcpl_430 OR and_dcpl_433 OR and_dcpl_437 OR and_dcpl_441 OR and_dcpl_444
      OR and_dcpl_447 OR mux_tmp_189);
  result_and_11_cse <= ccs_ccore_en AND (and_dcpl_452 OR and_dcpl_455 OR and_dcpl_458
      OR and_dcpl_462 OR and_dcpl_464 OR and_dcpl_468 OR and_dcpl_472 OR and_dcpl_474
      OR and_dcpl_476 OR mux_tmp_227);
  result_and_13_cse <= ccs_ccore_en AND (and_dcpl_480 OR and_dcpl_484 OR and_dcpl_488
      OR and_dcpl_491 OR and_dcpl_493 OR and_dcpl_496 OR and_dcpl_499 OR and_dcpl_501
      OR and_dcpl_503 OR mux_tmp_265);
  result_and_15_cse <= ccs_ccore_en AND (and_dcpl_507 OR and_dcpl_510 OR and_dcpl_513
      OR and_dcpl_516 OR and_dcpl_518 OR and_dcpl_521 OR and_dcpl_524 OR and_dcpl_526
      OR and_dcpl_528 OR mux_tmp_303);
  result_and_17_cse <= ccs_ccore_en AND (and_dcpl_533 OR and_dcpl_536 OR and_dcpl_539
      OR and_dcpl_542 OR and_dcpl_546 OR and_dcpl_549 OR and_dcpl_552 OR and_dcpl_556
      OR and_dcpl_560 OR mux_tmp_348);
  result_and_19_cse <= ccs_ccore_en AND (and_dcpl_566 OR and_dcpl_568 OR and_dcpl_570
      OR and_dcpl_572 OR and_dcpl_576 OR and_dcpl_578 OR and_dcpl_580 OR and_dcpl_583
      OR and_dcpl_586 OR mux_tmp_393);
  result_and_21_cse <= ccs_ccore_en AND (and_dcpl_590 OR and_dcpl_592 OR and_dcpl_594
      OR and_dcpl_596 OR and_dcpl_599 OR and_dcpl_601 OR and_dcpl_603 OR and_dcpl_607
      OR and_dcpl_611 OR mux_tmp_438);
  m_and_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_2;
  m_and_1_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_6;
  m_and_2_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_9;
  m_and_3_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_11;
  m_and_4_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_2;
  m_and_5_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_6;
  m_and_6_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_9;
  m_and_7_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_11;
  m_and_8_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (NOT (result_rem_11cyc_st_9(0)));
  m_and_9_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (result_rem_11cyc_st_9(0));
  m_and_10_cse <= ccs_ccore_en AND and_dcpl_4 AND (result_rem_11cyc_st_9(3)) AND
      (result_rem_11cyc_st_9(1)) AND (NOT (result_rem_11cyc_st_9(0)));
  m_and_11_cse <= ccs_ccore_en AND and_dcpl_30;
  m_and_12_cse <= ccs_ccore_en AND and_dcpl_32;
  m_and_13_cse <= ccs_ccore_en AND and_dcpl_35;
  m_and_14_cse <= ccs_ccore_en AND and_dcpl_37;
  m_and_15_cse <= ccs_ccore_en AND and_dcpl_39;
  m_and_16_cse <= ccs_ccore_en AND and_dcpl_40;
  m_and_17_cse <= ccs_ccore_en AND and_dcpl_41;
  m_and_18_cse <= ccs_ccore_en AND and_dcpl_42;
  m_and_19_cse <= ccs_ccore_en AND and_dcpl_45;
  m_and_20_cse <= ccs_ccore_en AND and_dcpl_47;
  m_and_21_cse <= ccs_ccore_en AND and_dcpl_50;
  m_and_22_cse <= ccs_ccore_en AND and_dcpl_55;
  m_and_23_cse <= ccs_ccore_en AND and_dcpl_58;
  m_and_24_cse <= ccs_ccore_en AND and_dcpl_60;
  m_and_25_cse <= ccs_ccore_en AND and_dcpl_62;
  m_and_26_cse <= ccs_ccore_en AND and_dcpl_65;
  m_and_27_cse <= ccs_ccore_en AND and_dcpl_68;
  m_and_28_cse <= ccs_ccore_en AND and_dcpl_70;
  m_and_29_cse <= ccs_ccore_en AND and_dcpl_72;
  m_and_30_cse <= ccs_ccore_en AND and_dcpl_74;
  m_and_31_cse <= ccs_ccore_en AND and_dcpl_75;
  m_and_32_cse <= ccs_ccore_en AND and_dcpl_76;
  m_and_33_cse <= ccs_ccore_en AND and_dcpl_81;
  m_and_34_cse <= ccs_ccore_en AND and_dcpl_84;
  m_and_35_cse <= ccs_ccore_en AND and_dcpl_86;
  m_and_36_cse <= ccs_ccore_en AND and_dcpl_88;
  m_and_37_cse <= ccs_ccore_en AND and_dcpl_91;
  m_and_38_cse <= ccs_ccore_en AND and_dcpl_94;
  m_and_39_cse <= ccs_ccore_en AND and_dcpl_96;
  m_and_40_cse <= ccs_ccore_en AND and_dcpl_98;
  m_and_41_cse <= ccs_ccore_en AND and_dcpl_100;
  m_and_42_cse <= ccs_ccore_en AND and_dcpl_101;
  m_and_43_cse <= ccs_ccore_en AND and_dcpl_102;
  m_and_44_cse <= ccs_ccore_en AND and_dcpl_107;
  m_and_45_cse <= ccs_ccore_en AND and_dcpl_110;
  m_and_46_cse <= ccs_ccore_en AND and_dcpl_112;
  m_and_47_cse <= ccs_ccore_en AND and_dcpl_114;
  m_and_48_cse <= ccs_ccore_en AND and_dcpl_116;
  m_and_49_cse <= ccs_ccore_en AND and_dcpl_117;
  m_and_50_cse <= ccs_ccore_en AND and_dcpl_118;
  m_and_51_cse <= ccs_ccore_en AND and_dcpl_119;
  m_and_52_cse <= ccs_ccore_en AND and_dcpl_122;
  m_and_53_cse <= ccs_ccore_en AND and_dcpl_125;
  m_and_54_cse <= ccs_ccore_en AND and_dcpl_127;
  m_and_55_cse <= ccs_ccore_en AND and_dcpl_132;
  m_and_56_cse <= ccs_ccore_en AND and_dcpl_135;
  m_and_57_cse <= ccs_ccore_en AND and_dcpl_137;
  m_and_58_cse <= ccs_ccore_en AND and_dcpl_139;
  m_and_59_cse <= ccs_ccore_en AND and_dcpl_142;
  m_and_60_cse <= ccs_ccore_en AND and_dcpl_145;
  m_and_61_cse <= ccs_ccore_en AND and_dcpl_147;
  m_and_62_cse <= ccs_ccore_en AND and_dcpl_149;
  m_and_63_cse <= ccs_ccore_en AND and_dcpl_151;
  m_and_64_cse <= ccs_ccore_en AND and_dcpl_152;
  m_and_65_cse <= ccs_ccore_en AND and_dcpl_153;
  m_and_66_cse <= ccs_ccore_en AND and_dcpl_158;
  m_and_67_cse <= ccs_ccore_en AND and_dcpl_160;
  m_and_68_cse <= ccs_ccore_en AND and_dcpl_163;
  m_and_69_cse <= ccs_ccore_en AND and_dcpl_165;
  m_and_70_cse <= ccs_ccore_en AND and_dcpl_168;
  m_and_71_cse <= ccs_ccore_en AND and_dcpl_170;
  m_and_72_cse <= ccs_ccore_en AND and_dcpl_173;
  m_and_73_cse <= ccs_ccore_en AND and_dcpl_175;
  m_and_74_cse <= ccs_ccore_en AND and_dcpl_177;
  m_and_75_cse <= ccs_ccore_en AND and_dcpl_178;
  m_and_76_cse <= ccs_ccore_en AND and_dcpl_179;
  m_and_77_cse <= ccs_ccore_en AND and_dcpl_184;
  m_and_78_cse <= ccs_ccore_en AND and_dcpl_186;
  m_and_79_cse <= ccs_ccore_en AND and_dcpl_189;
  m_and_80_cse <= ccs_ccore_en AND and_dcpl_191;
  m_and_81_cse <= ccs_ccore_en AND and_dcpl_194;
  m_and_82_cse <= ccs_ccore_en AND and_dcpl_196;
  m_and_83_cse <= ccs_ccore_en AND and_dcpl_199;
  m_and_84_cse <= ccs_ccore_en AND and_dcpl_201;
  m_and_85_cse <= ccs_ccore_en AND and_dcpl_203;
  m_and_86_cse <= ccs_ccore_en AND and_dcpl_204;
  m_and_87_cse <= ccs_ccore_en AND and_dcpl_205;
  m_and_88_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_207;
  m_and_89_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_212;
  m_and_90_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_214;
  m_and_91_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_211 AND (result_rem_11cyc(1));
  m_and_92_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_218 AND (NOT (result_rem_11cyc(1)));
  m_and_93_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_221 AND (NOT (result_rem_11cyc(1)));
  m_and_94_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_218 AND (result_rem_11cyc(1));
  m_and_95_cse <= ccs_ccore_en AND and_dcpl_209 AND and_dcpl_221 AND (result_rem_11cyc(1));
  m_and_96_cse <= ccs_ccore_en AND and_dcpl_228 AND and_dcpl_207;
  m_and_97_cse <= ccs_ccore_en AND and_dcpl_228 AND and_dcpl_212;
  m_and_98_cse <= ccs_ccore_en AND and_dcpl_228 AND and_dcpl_214;
  result_result_acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(CONV_SIGNED(CONV_SIGNED(result_acc_imod_1(3),
      1),2)), 2), 4) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(result_acc_imod_1(2 DOWNTO
      0)), 3), 4), 4));
  result_acc_imod_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(result_acc_idiv_1(2
      DOWNTO 0)), 3), 4) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED((NOT (result_acc_idiv_1(3)))
      & STD_LOGIC_VECTOR'( "00")), 3), 4) + CONV_SIGNED(CONV_SIGNED(SIGNED(STD_LOGIC_VECTOR'(
      "10") & (result_acc_idiv_1(3))), 3), 4), 4));
  result_acc_idiv_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(result_rem_11cyc)
      + UNSIGNED'( "0001"), 4));
  and_dcpl_1 <= NOT((result_rem_11cyc_st_9(3)) OR (result_rem_11cyc_st_9(1)));
  and_dcpl_2 <= and_dcpl_1 AND (NOT (result_rem_11cyc_st_9(0)));
  and_dcpl_3 <= main_stage_0_10 AND asn_itm_9;
  and_dcpl_4 <= and_dcpl_3 AND (NOT (result_rem_11cyc_st_9(2)));
  and_dcpl_6 <= and_dcpl_1 AND (result_rem_11cyc_st_9(0));
  and_dcpl_8 <= (NOT (result_rem_11cyc_st_9(3))) AND (result_rem_11cyc_st_9(1));
  and_dcpl_9 <= and_dcpl_8 AND (NOT (result_rem_11cyc_st_9(0)));
  and_dcpl_11 <= and_dcpl_8 AND (result_rem_11cyc_st_9(0));
  and_dcpl_13 <= and_dcpl_3 AND (result_rem_11cyc_st_9(2));
  and_dcpl_18 <= (result_rem_11cyc_st_9(3)) AND (NOT (result_rem_11cyc_st_9(1)));
  and_dcpl_26 <= NOT((result_rem_11cyc_st_8(3)) OR (result_rem_11cyc_st_8(1)));
  and_dcpl_27 <= and_dcpl_26 AND (NOT (result_rem_11cyc_st_8(0)));
  and_dcpl_28 <= main_stage_0_9 AND asn_itm_8;
  and_dcpl_29 <= and_dcpl_28 AND (NOT (result_rem_11cyc_st_8(2)));
  and_dcpl_30 <= and_dcpl_29 AND and_dcpl_27;
  and_dcpl_31 <= and_dcpl_26 AND (result_rem_11cyc_st_8(0));
  and_dcpl_32 <= and_dcpl_29 AND and_dcpl_31;
  and_dcpl_33 <= (NOT (result_rem_11cyc_st_8(3))) AND (result_rem_11cyc_st_8(1));
  and_dcpl_34 <= and_dcpl_33 AND (NOT (result_rem_11cyc_st_8(0)));
  and_dcpl_35 <= and_dcpl_29 AND and_dcpl_34;
  and_dcpl_36 <= and_dcpl_33 AND (result_rem_11cyc_st_8(0));
  and_dcpl_37 <= and_dcpl_29 AND and_dcpl_36;
  and_dcpl_38 <= and_dcpl_28 AND (result_rem_11cyc_st_8(2));
  and_dcpl_39 <= and_dcpl_38 AND and_dcpl_27;
  and_dcpl_40 <= and_dcpl_38 AND and_dcpl_31;
  and_dcpl_41 <= and_dcpl_38 AND and_dcpl_34;
  and_dcpl_42 <= and_dcpl_38 AND and_dcpl_36;
  and_dcpl_43 <= (result_rem_11cyc_st_8(3)) AND (NOT (result_rem_11cyc_st_8(1)));
  and_dcpl_45 <= and_dcpl_29 AND and_dcpl_43 AND (NOT (result_rem_11cyc_st_8(0)));
  and_dcpl_47 <= and_dcpl_29 AND and_dcpl_43 AND (result_rem_11cyc_st_8(0));
  and_dcpl_50 <= and_dcpl_29 AND (result_rem_11cyc_st_8(3)) AND (result_rem_11cyc_st_8(1))
      AND (NOT (result_rem_11cyc_st_8(0)));
  and_dcpl_51 <= NOT((result_rem_11cyc_st_7(2)) OR (result_rem_11cyc_st_7(0)));
  and_dcpl_52 <= and_dcpl_51 AND (NOT (result_rem_11cyc_st_7(1)));
  and_dcpl_53 <= main_stage_0_8 AND asn_itm_7;
  and_dcpl_54 <= and_dcpl_53 AND (NOT (result_rem_11cyc_st_7(3)));
  and_dcpl_55 <= and_dcpl_54 AND and_dcpl_52;
  and_dcpl_56 <= (NOT (result_rem_11cyc_st_7(2))) AND (result_rem_11cyc_st_7(0));
  and_dcpl_57 <= and_dcpl_56 AND (NOT (result_rem_11cyc_st_7(1)));
  and_dcpl_58 <= and_dcpl_54 AND and_dcpl_57;
  and_dcpl_59 <= and_dcpl_51 AND (result_rem_11cyc_st_7(1));
  and_dcpl_60 <= and_dcpl_54 AND and_dcpl_59;
  and_dcpl_62 <= and_dcpl_54 AND and_dcpl_56 AND (result_rem_11cyc_st_7(1));
  and_dcpl_63 <= (result_rem_11cyc_st_7(2)) AND (NOT (result_rem_11cyc_st_7(0)));
  and_dcpl_65 <= and_dcpl_54 AND and_dcpl_63 AND (NOT (result_rem_11cyc_st_7(1)));
  and_dcpl_66 <= (result_rem_11cyc_st_7(2)) AND (result_rem_11cyc_st_7(0));
  and_dcpl_68 <= and_dcpl_54 AND and_dcpl_66 AND (NOT (result_rem_11cyc_st_7(1)));
  and_dcpl_70 <= and_dcpl_54 AND and_dcpl_63 AND (result_rem_11cyc_st_7(1));
  and_dcpl_72 <= and_dcpl_54 AND and_dcpl_66 AND (result_rem_11cyc_st_7(1));
  and_dcpl_73 <= and_dcpl_53 AND (result_rem_11cyc_st_7(3));
  and_dcpl_74 <= and_dcpl_73 AND and_dcpl_52;
  and_dcpl_75 <= and_dcpl_73 AND and_dcpl_57;
  and_dcpl_76 <= and_dcpl_73 AND and_dcpl_59;
  and_dcpl_77 <= NOT((result_rem_11cyc_st_6(2)) OR (result_rem_11cyc_st_6(0)));
  and_dcpl_78 <= and_dcpl_77 AND (NOT (result_rem_11cyc_st_6(1)));
  and_dcpl_79 <= main_stage_0_7 AND asn_itm_6;
  and_dcpl_80 <= and_dcpl_79 AND (NOT (result_rem_11cyc_st_6(3)));
  and_dcpl_81 <= and_dcpl_80 AND and_dcpl_78;
  and_dcpl_82 <= (NOT (result_rem_11cyc_st_6(2))) AND (result_rem_11cyc_st_6(0));
  and_dcpl_83 <= and_dcpl_82 AND (NOT (result_rem_11cyc_st_6(1)));
  and_dcpl_84 <= and_dcpl_80 AND and_dcpl_83;
  and_dcpl_85 <= and_dcpl_77 AND (result_rem_11cyc_st_6(1));
  and_dcpl_86 <= and_dcpl_80 AND and_dcpl_85;
  and_dcpl_88 <= and_dcpl_80 AND and_dcpl_82 AND (result_rem_11cyc_st_6(1));
  and_dcpl_89 <= (result_rem_11cyc_st_6(2)) AND (NOT (result_rem_11cyc_st_6(0)));
  and_dcpl_91 <= and_dcpl_80 AND and_dcpl_89 AND (NOT (result_rem_11cyc_st_6(1)));
  and_dcpl_92 <= (result_rem_11cyc_st_6(2)) AND (result_rem_11cyc_st_6(0));
  and_dcpl_94 <= and_dcpl_80 AND and_dcpl_92 AND (NOT (result_rem_11cyc_st_6(1)));
  and_dcpl_96 <= and_dcpl_80 AND and_dcpl_89 AND (result_rem_11cyc_st_6(1));
  and_dcpl_98 <= and_dcpl_80 AND and_dcpl_92 AND (result_rem_11cyc_st_6(1));
  and_dcpl_99 <= and_dcpl_79 AND (result_rem_11cyc_st_6(3));
  and_dcpl_100 <= and_dcpl_99 AND and_dcpl_78;
  and_dcpl_101 <= and_dcpl_99 AND and_dcpl_83;
  and_dcpl_102 <= and_dcpl_99 AND and_dcpl_85;
  and_dcpl_103 <= NOT((result_rem_11cyc_st_5(3)) OR (result_rem_11cyc_st_5(0)));
  and_dcpl_104 <= and_dcpl_103 AND (NOT (result_rem_11cyc_st_5(1)));
  and_dcpl_105 <= main_stage_0_6 AND asn_itm_5;
  and_dcpl_106 <= and_dcpl_105 AND (NOT (result_rem_11cyc_st_5(2)));
  and_dcpl_107 <= and_dcpl_106 AND and_dcpl_104;
  and_dcpl_108 <= (NOT (result_rem_11cyc_st_5(3))) AND (result_rem_11cyc_st_5(0));
  and_dcpl_109 <= and_dcpl_108 AND (NOT (result_rem_11cyc_st_5(1)));
  and_dcpl_110 <= and_dcpl_106 AND and_dcpl_109;
  and_dcpl_111 <= and_dcpl_103 AND (result_rem_11cyc_st_5(1));
  and_dcpl_112 <= and_dcpl_106 AND and_dcpl_111;
  and_dcpl_113 <= and_dcpl_108 AND (result_rem_11cyc_st_5(1));
  and_dcpl_114 <= and_dcpl_106 AND and_dcpl_113;
  and_dcpl_115 <= and_dcpl_105 AND (result_rem_11cyc_st_5(2));
  and_dcpl_116 <= and_dcpl_115 AND and_dcpl_104;
  and_dcpl_117 <= and_dcpl_115 AND and_dcpl_109;
  and_dcpl_118 <= and_dcpl_115 AND and_dcpl_111;
  and_dcpl_119 <= and_dcpl_115 AND and_dcpl_113;
  and_dcpl_120 <= (result_rem_11cyc_st_5(3)) AND (NOT (result_rem_11cyc_st_5(0)));
  and_dcpl_122 <= and_dcpl_106 AND and_dcpl_120 AND (NOT (result_rem_11cyc_st_5(1)));
  and_dcpl_125 <= and_dcpl_106 AND (result_rem_11cyc_st_5(3)) AND (result_rem_11cyc_st_5(0))
      AND (NOT (result_rem_11cyc_st_5(1)));
  and_dcpl_127 <= and_dcpl_106 AND and_dcpl_120 AND (result_rem_11cyc_st_5(1));
  and_dcpl_128 <= NOT((result_rem_11cyc_st_4(2)) OR (result_rem_11cyc_st_4(0)));
  and_dcpl_129 <= and_dcpl_128 AND (NOT (result_rem_11cyc_st_4(1)));
  and_dcpl_130 <= main_stage_0_5 AND asn_itm_4;
  and_dcpl_131 <= and_dcpl_130 AND (NOT (result_rem_11cyc_st_4(3)));
  and_dcpl_132 <= and_dcpl_131 AND and_dcpl_129;
  and_dcpl_133 <= (NOT (result_rem_11cyc_st_4(2))) AND (result_rem_11cyc_st_4(0));
  and_dcpl_134 <= and_dcpl_133 AND (NOT (result_rem_11cyc_st_4(1)));
  and_dcpl_135 <= and_dcpl_131 AND and_dcpl_134;
  and_dcpl_136 <= and_dcpl_128 AND (result_rem_11cyc_st_4(1));
  and_dcpl_137 <= and_dcpl_131 AND and_dcpl_136;
  and_dcpl_139 <= and_dcpl_131 AND and_dcpl_133 AND (result_rem_11cyc_st_4(1));
  and_dcpl_140 <= (result_rem_11cyc_st_4(2)) AND (NOT (result_rem_11cyc_st_4(0)));
  and_dcpl_142 <= and_dcpl_131 AND and_dcpl_140 AND (NOT (result_rem_11cyc_st_4(1)));
  and_dcpl_143 <= (result_rem_11cyc_st_4(2)) AND (result_rem_11cyc_st_4(0));
  and_dcpl_145 <= and_dcpl_131 AND and_dcpl_143 AND (NOT (result_rem_11cyc_st_4(1)));
  and_dcpl_147 <= and_dcpl_131 AND and_dcpl_140 AND (result_rem_11cyc_st_4(1));
  and_dcpl_149 <= and_dcpl_131 AND and_dcpl_143 AND (result_rem_11cyc_st_4(1));
  and_dcpl_150 <= and_dcpl_130 AND (result_rem_11cyc_st_4(3));
  and_dcpl_151 <= and_dcpl_150 AND and_dcpl_129;
  and_dcpl_152 <= and_dcpl_150 AND and_dcpl_134;
  and_dcpl_153 <= and_dcpl_150 AND and_dcpl_136;
  and_dcpl_154 <= NOT(CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_155 <= and_dcpl_154 AND (NOT (result_rem_11cyc_st_3(0)));
  and_dcpl_156 <= main_stage_0_4 AND asn_itm_3;
  and_dcpl_157 <= and_dcpl_156 AND (NOT (result_rem_11cyc_st_3(3)));
  and_dcpl_158 <= and_dcpl_157 AND and_dcpl_155;
  and_dcpl_159 <= and_dcpl_154 AND (result_rem_11cyc_st_3(0));
  and_dcpl_160 <= and_dcpl_157 AND and_dcpl_159;
  and_dcpl_161 <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_162 <= and_dcpl_161 AND (NOT (result_rem_11cyc_st_3(0)));
  and_dcpl_163 <= and_dcpl_157 AND and_dcpl_162;
  and_dcpl_165 <= and_dcpl_157 AND and_dcpl_161 AND (result_rem_11cyc_st_3(0));
  and_dcpl_166 <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_168 <= and_dcpl_157 AND and_dcpl_166 AND (NOT (result_rem_11cyc_st_3(0)));
  and_dcpl_170 <= and_dcpl_157 AND and_dcpl_166 AND (result_rem_11cyc_st_3(0));
  and_dcpl_171 <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_173 <= and_dcpl_157 AND and_dcpl_171 AND (NOT (result_rem_11cyc_st_3(0)));
  and_dcpl_175 <= and_dcpl_157 AND and_dcpl_171 AND (result_rem_11cyc_st_3(0));
  and_dcpl_176 <= and_dcpl_156 AND (result_rem_11cyc_st_3(3));
  and_dcpl_177 <= and_dcpl_176 AND and_dcpl_155;
  and_dcpl_178 <= and_dcpl_176 AND and_dcpl_159;
  and_dcpl_179 <= and_dcpl_176 AND and_dcpl_162;
  and_dcpl_180 <= NOT(CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_181 <= and_dcpl_180 AND (NOT (result_rem_11cyc_st_2(0)));
  and_dcpl_182 <= main_stage_0_3 AND asn_itm_2;
  and_dcpl_183 <= and_dcpl_182 AND (NOT (result_rem_11cyc_st_2(3)));
  and_dcpl_184 <= and_dcpl_183 AND and_dcpl_181;
  and_dcpl_185 <= and_dcpl_180 AND (result_rem_11cyc_st_2(0));
  and_dcpl_186 <= and_dcpl_183 AND and_dcpl_185;
  and_dcpl_187 <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_188 <= and_dcpl_187 AND (NOT (result_rem_11cyc_st_2(0)));
  and_dcpl_189 <= and_dcpl_183 AND and_dcpl_188;
  and_dcpl_191 <= and_dcpl_183 AND and_dcpl_187 AND (result_rem_11cyc_st_2(0));
  and_dcpl_192 <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_194 <= and_dcpl_183 AND and_dcpl_192 AND (NOT (result_rem_11cyc_st_2(0)));
  and_dcpl_196 <= and_dcpl_183 AND and_dcpl_192 AND (result_rem_11cyc_st_2(0));
  and_dcpl_197 <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_199 <= and_dcpl_183 AND and_dcpl_197 AND (NOT (result_rem_11cyc_st_2(0)));
  and_dcpl_201 <= and_dcpl_183 AND and_dcpl_197 AND (result_rem_11cyc_st_2(0));
  and_dcpl_202 <= and_dcpl_182 AND (result_rem_11cyc_st_2(3));
  and_dcpl_203 <= and_dcpl_202 AND and_dcpl_181;
  and_dcpl_204 <= and_dcpl_202 AND and_dcpl_185;
  and_dcpl_205 <= and_dcpl_202 AND and_dcpl_188;
  and_dcpl_206 <= NOT((result_rem_11cyc(2)) OR (result_rem_11cyc(0)));
  and_dcpl_207 <= and_dcpl_206 AND (NOT (result_rem_11cyc(1)));
  and_dcpl_208 <= main_stage_0_2 AND asn_itm_1;
  and_dcpl_209 <= and_dcpl_208 AND (NOT (result_rem_11cyc(3)));
  and_dcpl_211 <= (NOT (result_rem_11cyc(2))) AND (result_rem_11cyc(0));
  and_dcpl_212 <= and_dcpl_211 AND (NOT (result_rem_11cyc(1)));
  and_dcpl_214 <= and_dcpl_206 AND (result_rem_11cyc(1));
  and_dcpl_218 <= (result_rem_11cyc(2)) AND (NOT (result_rem_11cyc(0)));
  and_dcpl_221 <= (result_rem_11cyc(2)) AND (result_rem_11cyc(0));
  and_dcpl_228 <= and_dcpl_208 AND (result_rem_11cyc(3));
  and_dcpl_232 <= NOT(CONV_SL_1_1(result_rem_11cyc_st_11(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_233 <= and_dcpl_232 AND (NOT (result_rem_11cyc_st_11(0)));
  and_dcpl_234 <= main_stage_0_12 AND asn_itm_11;
  and_dcpl_235 <= and_dcpl_234 AND (NOT (result_rem_11cyc_st_11(3)));
  and_dcpl_237 <= and_dcpl_232 AND (result_rem_11cyc_st_11(0));
  and_dcpl_239 <= CONV_SL_1_1(result_rem_11cyc_st_11(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_240 <= and_dcpl_239 AND (NOT (result_rem_11cyc_st_11(0)));
  and_dcpl_244 <= CONV_SL_1_1(result_rem_11cyc_st_11(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_249 <= CONV_SL_1_1(result_rem_11cyc_st_11(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_254 <= and_dcpl_234 AND (result_rem_11cyc_st_11(3));
  and_dcpl_260 <= NOT(CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_261 <= ccs_ccore_start_rsci_idat AND (NOT (result_result_acc_tmp(2)));
  and_dcpl_262 <= and_dcpl_261 AND (NOT (result_result_acc_tmp(3)));
  and_dcpl_263 <= and_dcpl_262 AND and_dcpl_260;
  or_tmp_2 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0000")) OR (NOT and_dcpl_208);
  or_3_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0000"));
  nor_691_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_2));
  mux_nl <= MUX_s_1_2_2(nor_691_nl, or_tmp_2, or_3_cse);
  and_dcpl_269 <= mux_nl AND and_dcpl_184;
  or_8_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0000"));
  nor_690_nl <= NOT(and_dcpl_208 OR and_dcpl_184);
  or_10_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_182);
  mux_tmp_1 <= MUX_s_1_2_2(nor_690_nl, or_10_nl, or_8_cse);
  nor_689_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_1));
  mux_2_nl <= MUX_s_1_2_2(nor_689_nl, mux_tmp_1, or_3_cse);
  and_dcpl_275 <= mux_2_nl AND and_dcpl_158;
  or_15_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0000"));
  nor_687_nl <= NOT(and_dcpl_182 OR and_dcpl_158);
  or_17_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_156);
  mux_tmp_3 <= MUX_s_1_2_2(nor_687_nl, or_17_nl, or_15_cse);
  nor_688_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_3));
  mux_tmp_4 <= MUX_s_1_2_2(nor_688_nl, mux_tmp_3, or_8_cse);
  nor_686_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_4));
  mux_5_nl <= MUX_s_1_2_2(nor_686_nl, mux_tmp_4, or_3_cse);
  and_dcpl_281 <= mux_5_nl AND and_dcpl_132;
  or_24_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0000"));
  nor_683_nl <= NOT(and_dcpl_156 OR and_dcpl_132);
  or_26_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_130);
  mux_tmp_6 <= MUX_s_1_2_2(nor_683_nl, or_26_nl, or_24_cse);
  nor_684_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_6));
  mux_tmp_7 <= MUX_s_1_2_2(nor_684_nl, mux_tmp_6, or_15_cse);
  nor_685_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_7));
  mux_tmp_8 <= MUX_s_1_2_2(nor_685_nl, mux_tmp_7, or_8_cse);
  nor_682_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_8));
  mux_9_nl <= MUX_s_1_2_2(nor_682_nl, mux_tmp_8, or_3_cse);
  and_dcpl_287 <= mux_9_nl AND and_dcpl_107;
  or_35_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0000"));
  nor_678_nl <= NOT(and_dcpl_130 OR and_dcpl_107);
  or_37_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_105);
  mux_tmp_10 <= MUX_s_1_2_2(nor_678_nl, or_37_nl, or_35_cse);
  nor_679_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_10));
  mux_tmp_11 <= MUX_s_1_2_2(nor_679_nl, mux_tmp_10, or_24_cse);
  nor_680_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_11));
  mux_tmp_12 <= MUX_s_1_2_2(nor_680_nl, mux_tmp_11, or_15_cse);
  nor_681_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_12));
  mux_tmp_13 <= MUX_s_1_2_2(nor_681_nl, mux_tmp_12, or_8_cse);
  nor_677_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_13));
  mux_14_nl <= MUX_s_1_2_2(nor_677_nl, mux_tmp_13, or_3_cse);
  and_dcpl_293 <= mux_14_nl AND and_dcpl_81;
  or_48_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0000"));
  nor_672_nl <= NOT(and_dcpl_105 OR and_dcpl_81);
  or_50_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_79);
  mux_tmp_15 <= MUX_s_1_2_2(nor_672_nl, or_50_nl, or_48_cse);
  nor_673_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_15));
  mux_tmp_16 <= MUX_s_1_2_2(nor_673_nl, mux_tmp_15, or_35_cse);
  nor_674_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_16));
  mux_tmp_17 <= MUX_s_1_2_2(nor_674_nl, mux_tmp_16, or_24_cse);
  nor_675_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_17));
  mux_tmp_18 <= MUX_s_1_2_2(nor_675_nl, mux_tmp_17, or_15_cse);
  nor_676_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_18));
  mux_tmp_19 <= MUX_s_1_2_2(nor_676_nl, mux_tmp_18, or_8_cse);
  nor_671_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_19));
  mux_20_nl <= MUX_s_1_2_2(nor_671_nl, mux_tmp_19, or_3_cse);
  and_dcpl_299 <= mux_20_nl AND and_dcpl_55;
  or_63_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0000"));
  nor_665_nl <= NOT(and_dcpl_79 OR and_dcpl_55);
  or_65_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_53);
  mux_tmp_21 <= MUX_s_1_2_2(nor_665_nl, or_65_nl, or_63_cse);
  nor_666_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_21));
  mux_tmp_22 <= MUX_s_1_2_2(nor_666_nl, mux_tmp_21, or_48_cse);
  nor_667_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_22));
  mux_tmp_23 <= MUX_s_1_2_2(nor_667_nl, mux_tmp_22, or_35_cse);
  nor_668_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_23));
  mux_tmp_24 <= MUX_s_1_2_2(nor_668_nl, mux_tmp_23, or_24_cse);
  nor_669_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_24));
  mux_tmp_25 <= MUX_s_1_2_2(nor_669_nl, mux_tmp_24, or_15_cse);
  nor_670_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_25));
  mux_tmp_26 <= MUX_s_1_2_2(nor_670_nl, mux_tmp_25, or_8_cse);
  nor_664_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_26));
  mux_27_nl <= MUX_s_1_2_2(nor_664_nl, mux_tmp_26, or_3_cse);
  and_dcpl_305 <= mux_27_nl AND and_dcpl_30;
  nor_656_nl <= NOT(and_dcpl_53 OR and_dcpl_30);
  or_82_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0000")) OR (NOT
      and_dcpl_28);
  or_80_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0000"));
  mux_tmp_28 <= MUX_s_1_2_2(nor_656_nl, or_82_nl, or_80_nl);
  nor_657_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_28));
  mux_tmp_29 <= MUX_s_1_2_2(nor_657_nl, mux_tmp_28, or_63_cse);
  nor_658_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_29));
  mux_tmp_30 <= MUX_s_1_2_2(nor_658_nl, mux_tmp_29, or_48_cse);
  nor_659_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_30));
  mux_tmp_31 <= MUX_s_1_2_2(nor_659_nl, mux_tmp_30, or_35_cse);
  nor_660_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_31));
  mux_tmp_32 <= MUX_s_1_2_2(nor_660_nl, mux_tmp_31, or_24_cse);
  nor_661_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_32));
  mux_tmp_33 <= MUX_s_1_2_2(nor_661_nl, mux_tmp_32, or_15_cse);
  nor_662_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_33));
  mux_tmp_34 <= MUX_s_1_2_2(nor_662_nl, mux_tmp_33, or_8_cse);
  nor_663_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_34));
  mux_35_nl <= MUX_s_1_2_2(nor_663_nl, mux_tmp_34, or_3_cse);
  and_dcpl_311 <= mux_35_nl AND and_dcpl_4 AND and_dcpl_2;
  and_tmp_6 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0000")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0000")));
  nor_654_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_6));
  mux_tmp_36 <= MUX_s_1_2_2(nor_654_nl, and_tmp_6, or_8_cse);
  nor_655_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_36));
  mux_tmp_37 <= MUX_s_1_2_2(nor_655_nl, mux_tmp_36, or_3_cse);
  and_dcpl_318 <= CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_319 <= and_dcpl_262 AND and_dcpl_318;
  or_tmp_102 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_208);
  or_107_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0001"));
  nor_653_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_102));
  mux_38_nl <= MUX_s_1_2_2(nor_653_nl, or_tmp_102, or_107_cse);
  and_dcpl_322 <= mux_38_nl AND and_dcpl_186;
  or_112_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0001"));
  nor_652_nl <= NOT(and_dcpl_208 OR and_dcpl_186);
  or_114_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_182);
  mux_tmp_39 <= MUX_s_1_2_2(nor_652_nl, or_114_nl, or_112_cse);
  nor_651_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_39));
  mux_40_nl <= MUX_s_1_2_2(nor_651_nl, mux_tmp_39, or_107_cse);
  and_dcpl_325 <= mux_40_nl AND and_dcpl_160;
  or_119_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0001"));
  nor_649_nl <= NOT(and_dcpl_182 OR and_dcpl_160);
  or_121_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_156);
  mux_tmp_41 <= MUX_s_1_2_2(nor_649_nl, or_121_nl, or_119_cse);
  nor_650_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_41));
  mux_tmp_42 <= MUX_s_1_2_2(nor_650_nl, mux_tmp_41, or_112_cse);
  nor_648_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_42));
  mux_43_nl <= MUX_s_1_2_2(nor_648_nl, mux_tmp_42, or_107_cse);
  and_dcpl_329 <= mux_43_nl AND and_dcpl_135;
  or_128_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0001"));
  nor_645_nl <= NOT(and_dcpl_156 OR and_dcpl_135);
  or_130_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_130);
  mux_tmp_44 <= MUX_s_1_2_2(nor_645_nl, or_130_nl, or_128_cse);
  nor_646_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_44));
  mux_tmp_45 <= MUX_s_1_2_2(nor_646_nl, mux_tmp_44, or_119_cse);
  nor_647_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_45));
  mux_tmp_46 <= MUX_s_1_2_2(nor_647_nl, mux_tmp_45, or_112_cse);
  nor_644_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_46));
  mux_47_nl <= MUX_s_1_2_2(nor_644_nl, mux_tmp_46, or_107_cse);
  and_dcpl_333 <= mux_47_nl AND and_dcpl_110;
  or_139_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0001"));
  nor_640_nl <= NOT(and_dcpl_130 OR and_dcpl_110);
  or_141_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_105);
  mux_tmp_48 <= MUX_s_1_2_2(nor_640_nl, or_141_nl, or_139_cse);
  nor_641_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_48));
  mux_tmp_49 <= MUX_s_1_2_2(nor_641_nl, mux_tmp_48, or_128_cse);
  nor_642_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_49));
  mux_tmp_50 <= MUX_s_1_2_2(nor_642_nl, mux_tmp_49, or_119_cse);
  nor_643_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_50));
  mux_tmp_51 <= MUX_s_1_2_2(nor_643_nl, mux_tmp_50, or_112_cse);
  nor_639_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_51));
  mux_52_nl <= MUX_s_1_2_2(nor_639_nl, mux_tmp_51, or_107_cse);
  and_dcpl_337 <= mux_52_nl AND and_dcpl_84;
  or_152_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0001"));
  nor_634_nl <= NOT(and_dcpl_105 OR and_dcpl_84);
  or_154_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_79);
  mux_tmp_53 <= MUX_s_1_2_2(nor_634_nl, or_154_nl, or_152_cse);
  nor_635_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_53));
  mux_tmp_54 <= MUX_s_1_2_2(nor_635_nl, mux_tmp_53, or_139_cse);
  nor_636_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_54));
  mux_tmp_55 <= MUX_s_1_2_2(nor_636_nl, mux_tmp_54, or_128_cse);
  nor_637_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_55));
  mux_tmp_56 <= MUX_s_1_2_2(nor_637_nl, mux_tmp_55, or_119_cse);
  nor_638_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_56));
  mux_tmp_57 <= MUX_s_1_2_2(nor_638_nl, mux_tmp_56, or_112_cse);
  nor_633_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_57));
  mux_58_nl <= MUX_s_1_2_2(nor_633_nl, mux_tmp_57, or_107_cse);
  and_dcpl_341 <= mux_58_nl AND and_dcpl_58;
  or_167_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0001"));
  nor_627_nl <= NOT(and_dcpl_79 OR and_dcpl_58);
  or_169_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_53);
  mux_tmp_59 <= MUX_s_1_2_2(nor_627_nl, or_169_nl, or_167_cse);
  nor_628_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_59));
  mux_tmp_60 <= MUX_s_1_2_2(nor_628_nl, mux_tmp_59, or_152_cse);
  nor_629_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_60));
  mux_tmp_61 <= MUX_s_1_2_2(nor_629_nl, mux_tmp_60, or_139_cse);
  nor_630_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_61));
  mux_tmp_62 <= MUX_s_1_2_2(nor_630_nl, mux_tmp_61, or_128_cse);
  nor_631_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_62));
  mux_tmp_63 <= MUX_s_1_2_2(nor_631_nl, mux_tmp_62, or_119_cse);
  nor_632_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_63));
  mux_tmp_64 <= MUX_s_1_2_2(nor_632_nl, mux_tmp_63, or_112_cse);
  nor_626_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_64));
  mux_65_nl <= MUX_s_1_2_2(nor_626_nl, mux_tmp_64, or_107_cse);
  and_dcpl_344 <= mux_65_nl AND and_dcpl_32;
  nor_618_nl <= NOT(and_dcpl_53 OR and_dcpl_32);
  or_186_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      and_dcpl_28);
  or_184_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0001"));
  mux_tmp_66 <= MUX_s_1_2_2(nor_618_nl, or_186_nl, or_184_nl);
  nor_619_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_66));
  mux_tmp_67 <= MUX_s_1_2_2(nor_619_nl, mux_tmp_66, or_167_cse);
  nor_620_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_67));
  mux_tmp_68 <= MUX_s_1_2_2(nor_620_nl, mux_tmp_67, or_152_cse);
  nor_621_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_68));
  mux_tmp_69 <= MUX_s_1_2_2(nor_621_nl, mux_tmp_68, or_139_cse);
  nor_622_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_69));
  mux_tmp_70 <= MUX_s_1_2_2(nor_622_nl, mux_tmp_69, or_128_cse);
  nor_623_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_70));
  mux_tmp_71 <= MUX_s_1_2_2(nor_623_nl, mux_tmp_70, or_119_cse);
  nor_624_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_71));
  mux_tmp_72 <= MUX_s_1_2_2(nor_624_nl, mux_tmp_71, or_112_cse);
  nor_625_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_72));
  mux_73_nl <= MUX_s_1_2_2(nor_625_nl, mux_tmp_72, or_107_cse);
  and_dcpl_347 <= mux_73_nl AND and_dcpl_4 AND and_dcpl_6;
  and_tmp_13 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0001")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0001")));
  nor_617_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_13));
  mux_tmp_74 <= MUX_s_1_2_2(nor_617_nl, and_tmp_13, or_112_cse);
  nand_146_cse <= NOT((result_result_acc_tmp(0)) AND ccs_ccore_start_rsci_idat);
  and_797_nl <= nand_146_cse AND mux_tmp_74;
  or_195_nl <= CONV_SL_1_1(result_result_acc_tmp(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_75 <= MUX_s_1_2_2(and_797_nl, mux_tmp_74, or_195_nl);
  and_dcpl_352 <= CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_353 <= and_dcpl_262 AND and_dcpl_352;
  or_tmp_202 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_208);
  or_209_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0010"));
  nor_616_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_202));
  mux_76_nl <= MUX_s_1_2_2(nor_616_nl, or_tmp_202, or_209_cse);
  and_dcpl_357 <= mux_76_nl AND and_dcpl_189;
  or_214_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0010"));
  nor_615_nl <= NOT(and_dcpl_208 OR and_dcpl_189);
  or_216_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_182);
  mux_tmp_77 <= MUX_s_1_2_2(nor_615_nl, or_216_nl, or_214_cse);
  nor_614_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_77));
  mux_78_nl <= MUX_s_1_2_2(nor_614_nl, mux_tmp_77, or_209_cse);
  and_dcpl_361 <= mux_78_nl AND and_dcpl_163;
  or_221_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0010"));
  nor_612_nl <= NOT(and_dcpl_182 OR and_dcpl_163);
  or_223_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_156);
  mux_tmp_79 <= MUX_s_1_2_2(nor_612_nl, or_223_nl, or_221_cse);
  nor_613_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_79));
  mux_tmp_80 <= MUX_s_1_2_2(nor_613_nl, mux_tmp_79, or_214_cse);
  nor_611_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_80));
  mux_81_nl <= MUX_s_1_2_2(nor_611_nl, mux_tmp_80, or_209_cse);
  and_dcpl_364 <= mux_81_nl AND and_dcpl_137;
  or_230_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0010"));
  nor_608_nl <= NOT(and_dcpl_156 OR and_dcpl_137);
  or_232_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_130);
  mux_tmp_82 <= MUX_s_1_2_2(nor_608_nl, or_232_nl, or_230_cse);
  nor_609_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_82));
  mux_tmp_83 <= MUX_s_1_2_2(nor_609_nl, mux_tmp_82, or_221_cse);
  nor_610_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_83));
  mux_tmp_84 <= MUX_s_1_2_2(nor_610_nl, mux_tmp_83, or_214_cse);
  nor_607_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_84));
  mux_85_nl <= MUX_s_1_2_2(nor_607_nl, mux_tmp_84, or_209_cse);
  and_dcpl_367 <= mux_85_nl AND and_dcpl_112;
  or_241_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0010"));
  nor_603_nl <= NOT(and_dcpl_130 OR and_dcpl_112);
  or_243_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_105);
  mux_tmp_86 <= MUX_s_1_2_2(nor_603_nl, or_243_nl, or_241_cse);
  nor_604_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_86));
  mux_tmp_87 <= MUX_s_1_2_2(nor_604_nl, mux_tmp_86, or_230_cse);
  nor_605_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_87));
  mux_tmp_88 <= MUX_s_1_2_2(nor_605_nl, mux_tmp_87, or_221_cse);
  nor_606_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_88));
  mux_tmp_89 <= MUX_s_1_2_2(nor_606_nl, mux_tmp_88, or_214_cse);
  nor_602_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_89));
  mux_90_nl <= MUX_s_1_2_2(nor_602_nl, mux_tmp_89, or_209_cse);
  and_dcpl_370 <= mux_90_nl AND and_dcpl_86;
  or_254_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0010"));
  nor_597_nl <= NOT(and_dcpl_105 OR and_dcpl_86);
  or_256_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_79);
  mux_tmp_91 <= MUX_s_1_2_2(nor_597_nl, or_256_nl, or_254_cse);
  nor_598_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_91));
  mux_tmp_92 <= MUX_s_1_2_2(nor_598_nl, mux_tmp_91, or_241_cse);
  nor_599_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_92));
  mux_tmp_93 <= MUX_s_1_2_2(nor_599_nl, mux_tmp_92, or_230_cse);
  nor_600_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_93));
  mux_tmp_94 <= MUX_s_1_2_2(nor_600_nl, mux_tmp_93, or_221_cse);
  nor_601_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_94));
  mux_tmp_95 <= MUX_s_1_2_2(nor_601_nl, mux_tmp_94, or_214_cse);
  nor_596_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_95));
  mux_96_nl <= MUX_s_1_2_2(nor_596_nl, mux_tmp_95, or_209_cse);
  and_dcpl_373 <= mux_96_nl AND and_dcpl_60;
  or_269_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0010"));
  nor_590_nl <= NOT(and_dcpl_79 OR and_dcpl_60);
  or_271_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_53);
  mux_tmp_97 <= MUX_s_1_2_2(nor_590_nl, or_271_nl, or_269_cse);
  nor_591_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_97));
  mux_tmp_98 <= MUX_s_1_2_2(nor_591_nl, mux_tmp_97, or_254_cse);
  nor_592_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_98));
  mux_tmp_99 <= MUX_s_1_2_2(nor_592_nl, mux_tmp_98, or_241_cse);
  nor_593_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_99));
  mux_tmp_100 <= MUX_s_1_2_2(nor_593_nl, mux_tmp_99, or_230_cse);
  nor_594_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_100));
  mux_tmp_101 <= MUX_s_1_2_2(nor_594_nl, mux_tmp_100, or_221_cse);
  nor_595_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_101));
  mux_tmp_102 <= MUX_s_1_2_2(nor_595_nl, mux_tmp_101, or_214_cse);
  nor_589_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_102));
  mux_103_nl <= MUX_s_1_2_2(nor_589_nl, mux_tmp_102, or_209_cse);
  and_dcpl_377 <= mux_103_nl AND and_dcpl_35;
  nor_581_nl <= NOT(and_dcpl_53 OR and_dcpl_35);
  or_288_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      and_dcpl_28);
  or_286_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0010"));
  mux_tmp_104 <= MUX_s_1_2_2(nor_581_nl, or_288_nl, or_286_nl);
  nor_582_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_104));
  mux_tmp_105 <= MUX_s_1_2_2(nor_582_nl, mux_tmp_104, or_269_cse);
  nor_583_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_105));
  mux_tmp_106 <= MUX_s_1_2_2(nor_583_nl, mux_tmp_105, or_254_cse);
  nor_584_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_106));
  mux_tmp_107 <= MUX_s_1_2_2(nor_584_nl, mux_tmp_106, or_241_cse);
  nor_585_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_107));
  mux_tmp_108 <= MUX_s_1_2_2(nor_585_nl, mux_tmp_107, or_230_cse);
  nor_586_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_108));
  mux_tmp_109 <= MUX_s_1_2_2(nor_586_nl, mux_tmp_108, or_221_cse);
  nor_587_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_109));
  mux_tmp_110 <= MUX_s_1_2_2(nor_587_nl, mux_tmp_109, or_214_cse);
  nor_588_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_110));
  mux_111_nl <= MUX_s_1_2_2(nor_588_nl, mux_tmp_110, or_209_cse);
  and_dcpl_381 <= mux_111_nl AND and_dcpl_4 AND and_dcpl_9;
  and_tmp_20 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0010")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0010")));
  nor_579_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_20));
  mux_tmp_112 <= MUX_s_1_2_2(nor_579_nl, and_tmp_20, or_214_cse);
  nor_580_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_112));
  mux_tmp_113 <= MUX_s_1_2_2(nor_580_nl, mux_tmp_112, or_209_cse);
  and_dcpl_386 <= CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_387 <= and_dcpl_262 AND and_dcpl_386;
  or_tmp_302 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_208);
  or_311_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0011"));
  nor_578_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_302));
  mux_114_nl <= MUX_s_1_2_2(nor_578_nl, or_tmp_302, or_311_cse);
  and_dcpl_390 <= mux_114_nl AND and_dcpl_191;
  or_316_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0011"));
  nor_577_nl <= NOT(and_dcpl_208 OR and_dcpl_191);
  or_318_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_182);
  mux_tmp_115 <= MUX_s_1_2_2(nor_577_nl, or_318_nl, or_316_cse);
  nor_576_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_115));
  mux_116_nl <= MUX_s_1_2_2(nor_576_nl, mux_tmp_115, or_311_cse);
  and_dcpl_393 <= mux_116_nl AND and_dcpl_165;
  or_323_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0011"));
  nor_574_nl <= NOT(and_dcpl_182 OR and_dcpl_165);
  or_325_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_156);
  mux_tmp_117 <= MUX_s_1_2_2(nor_574_nl, or_325_nl, or_323_cse);
  nor_575_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_117));
  mux_tmp_118 <= MUX_s_1_2_2(nor_575_nl, mux_tmp_117, or_316_cse);
  nor_573_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_118));
  mux_119_nl <= MUX_s_1_2_2(nor_573_nl, mux_tmp_118, or_311_cse);
  and_dcpl_396 <= mux_119_nl AND and_dcpl_139;
  or_332_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0011"));
  nor_570_nl <= NOT(and_dcpl_156 OR and_dcpl_139);
  or_334_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_130);
  mux_tmp_120 <= MUX_s_1_2_2(nor_570_nl, or_334_nl, or_332_cse);
  nor_571_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_120));
  mux_tmp_121 <= MUX_s_1_2_2(nor_571_nl, mux_tmp_120, or_323_cse);
  nor_572_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_121));
  mux_tmp_122 <= MUX_s_1_2_2(nor_572_nl, mux_tmp_121, or_316_cse);
  nor_569_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_122));
  mux_123_nl <= MUX_s_1_2_2(nor_569_nl, mux_tmp_122, or_311_cse);
  and_dcpl_399 <= mux_123_nl AND and_dcpl_114;
  or_343_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0011"));
  nor_565_nl <= NOT(and_dcpl_130 OR and_dcpl_114);
  or_345_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_105);
  mux_tmp_124 <= MUX_s_1_2_2(nor_565_nl, or_345_nl, or_343_cse);
  nor_566_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_124));
  mux_tmp_125 <= MUX_s_1_2_2(nor_566_nl, mux_tmp_124, or_332_cse);
  nor_567_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_125));
  mux_tmp_126 <= MUX_s_1_2_2(nor_567_nl, mux_tmp_125, or_323_cse);
  nor_568_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_126));
  mux_tmp_127 <= MUX_s_1_2_2(nor_568_nl, mux_tmp_126, or_316_cse);
  nor_564_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_127));
  mux_128_nl <= MUX_s_1_2_2(nor_564_nl, mux_tmp_127, or_311_cse);
  and_dcpl_402 <= mux_128_nl AND and_dcpl_88;
  or_356_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0011"));
  nor_559_nl <= NOT(and_dcpl_105 OR and_dcpl_88);
  or_358_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_79);
  mux_tmp_129 <= MUX_s_1_2_2(nor_559_nl, or_358_nl, or_356_cse);
  nor_560_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_129));
  mux_tmp_130 <= MUX_s_1_2_2(nor_560_nl, mux_tmp_129, or_343_cse);
  nor_561_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_130));
  mux_tmp_131 <= MUX_s_1_2_2(nor_561_nl, mux_tmp_130, or_332_cse);
  nor_562_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_131));
  mux_tmp_132 <= MUX_s_1_2_2(nor_562_nl, mux_tmp_131, or_323_cse);
  nor_563_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_132));
  mux_tmp_133 <= MUX_s_1_2_2(nor_563_nl, mux_tmp_132, or_316_cse);
  nor_558_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_133));
  mux_134_nl <= MUX_s_1_2_2(nor_558_nl, mux_tmp_133, or_311_cse);
  and_dcpl_405 <= mux_134_nl AND and_dcpl_62;
  or_371_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0011"));
  nor_552_nl <= NOT(and_dcpl_79 OR and_dcpl_62);
  or_373_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_53);
  mux_tmp_135 <= MUX_s_1_2_2(nor_552_nl, or_373_nl, or_371_cse);
  nor_553_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_135));
  mux_tmp_136 <= MUX_s_1_2_2(nor_553_nl, mux_tmp_135, or_356_cse);
  nor_554_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_136));
  mux_tmp_137 <= MUX_s_1_2_2(nor_554_nl, mux_tmp_136, or_343_cse);
  nor_555_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_137));
  mux_tmp_138 <= MUX_s_1_2_2(nor_555_nl, mux_tmp_137, or_332_cse);
  nor_556_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_138));
  mux_tmp_139 <= MUX_s_1_2_2(nor_556_nl, mux_tmp_138, or_323_cse);
  nor_557_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_139));
  mux_tmp_140 <= MUX_s_1_2_2(nor_557_nl, mux_tmp_139, or_316_cse);
  nor_551_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_140));
  mux_141_nl <= MUX_s_1_2_2(nor_551_nl, mux_tmp_140, or_311_cse);
  and_dcpl_408 <= mux_141_nl AND and_dcpl_37;
  nor_543_nl <= NOT(and_dcpl_53 OR and_dcpl_37);
  or_390_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      and_dcpl_28);
  or_388_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0011"));
  mux_tmp_142 <= MUX_s_1_2_2(nor_543_nl, or_390_nl, or_388_nl);
  nor_544_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_142));
  mux_tmp_143 <= MUX_s_1_2_2(nor_544_nl, mux_tmp_142, or_371_cse);
  nor_545_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_143));
  mux_tmp_144 <= MUX_s_1_2_2(nor_545_nl, mux_tmp_143, or_356_cse);
  nor_546_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_144));
  mux_tmp_145 <= MUX_s_1_2_2(nor_546_nl, mux_tmp_144, or_343_cse);
  nor_547_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_145));
  mux_tmp_146 <= MUX_s_1_2_2(nor_547_nl, mux_tmp_145, or_332_cse);
  nor_548_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_146));
  mux_tmp_147 <= MUX_s_1_2_2(nor_548_nl, mux_tmp_146, or_323_cse);
  nor_549_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_147));
  mux_tmp_148 <= MUX_s_1_2_2(nor_549_nl, mux_tmp_147, or_316_cse);
  nor_550_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_148));
  mux_149_nl <= MUX_s_1_2_2(nor_550_nl, mux_tmp_148, or_311_cse);
  and_dcpl_411 <= mux_149_nl AND and_dcpl_4 AND and_dcpl_11;
  and_tmp_27 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0011")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0011")));
  nor_542_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_27));
  mux_tmp_150 <= MUX_s_1_2_2(nor_542_nl, and_tmp_27, or_316_cse);
  and_796_nl <= (NOT(CONV_SL_1_1(result_result_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND ccs_ccore_start_rsci_idat)) AND mux_tmp_150;
  or_399_nl <= CONV_SL_1_1(result_result_acc_tmp(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_151 <= MUX_s_1_2_2(and_796_nl, mux_tmp_150, or_399_nl);
  and_dcpl_417 <= ccs_ccore_start_rsci_idat AND CONV_SL_1_1(result_result_acc_tmp(3
      DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_418 <= and_dcpl_417 AND and_dcpl_260;
  or_tmp_402 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_208);
  nand_144_cse <= NOT((result_result_acc_tmp(2)) AND ccs_ccore_start_rsci_idat);
  or_413_cse <= (result_result_acc_tmp(1)) OR (result_result_acc_tmp(0)) OR (result_result_acc_tmp(3));
  and_795_nl <= nand_144_cse AND or_tmp_402;
  mux_152_nl <= MUX_s_1_2_2(and_795_nl, or_tmp_402, or_413_cse);
  and_dcpl_422 <= mux_152_nl AND and_dcpl_194;
  or_418_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0100"));
  nor_541_nl <= NOT(and_dcpl_208 OR and_dcpl_194);
  or_420_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_182);
  mux_tmp_153 <= MUX_s_1_2_2(nor_541_nl, or_420_nl, or_418_cse);
  and_794_nl <= nand_144_cse AND mux_tmp_153;
  mux_154_nl <= MUX_s_1_2_2(and_794_nl, mux_tmp_153, or_413_cse);
  and_dcpl_426 <= mux_154_nl AND and_dcpl_168;
  or_425_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0100"));
  nor_539_nl <= NOT(and_dcpl_182 OR and_dcpl_168);
  or_427_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_156);
  mux_tmp_155 <= MUX_s_1_2_2(nor_539_nl, or_427_nl, or_425_cse);
  nor_540_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_155));
  mux_tmp_156 <= MUX_s_1_2_2(nor_540_nl, mux_tmp_155, or_418_cse);
  and_793_nl <= nand_144_cse AND mux_tmp_156;
  mux_157_nl <= MUX_s_1_2_2(and_793_nl, mux_tmp_156, or_413_cse);
  and_dcpl_430 <= mux_157_nl AND and_dcpl_142;
  or_434_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0100"));
  nor_536_nl <= NOT(and_dcpl_156 OR and_dcpl_142);
  or_436_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_130);
  mux_tmp_158 <= MUX_s_1_2_2(nor_536_nl, or_436_nl, or_434_cse);
  nor_537_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_158));
  mux_tmp_159 <= MUX_s_1_2_2(nor_537_nl, mux_tmp_158, or_425_cse);
  nor_538_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_159));
  mux_tmp_160 <= MUX_s_1_2_2(nor_538_nl, mux_tmp_159, or_418_cse);
  and_792_nl <= nand_144_cse AND mux_tmp_160;
  mux_161_nl <= MUX_s_1_2_2(and_792_nl, mux_tmp_160, or_413_cse);
  and_dcpl_433 <= mux_161_nl AND and_dcpl_116;
  or_445_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0100"));
  nor_532_nl <= NOT(and_dcpl_130 OR and_dcpl_116);
  or_447_nl <= (result_rem_11cyc_st_5(1)) OR (result_rem_11cyc_st_5(0)) OR (result_rem_11cyc_st_5(3))
      OR (NOT and_dcpl_115);
  mux_tmp_162 <= MUX_s_1_2_2(nor_532_nl, or_447_nl, or_445_cse);
  nor_533_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_162));
  mux_tmp_163 <= MUX_s_1_2_2(nor_533_nl, mux_tmp_162, or_434_cse);
  nor_534_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_163));
  mux_tmp_164 <= MUX_s_1_2_2(nor_534_nl, mux_tmp_163, or_425_cse);
  nor_535_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_164));
  mux_tmp_165 <= MUX_s_1_2_2(nor_535_nl, mux_tmp_164, or_418_cse);
  and_791_nl <= nand_144_cse AND mux_tmp_165;
  mux_166_nl <= MUX_s_1_2_2(and_791_nl, mux_tmp_165, or_413_cse);
  and_dcpl_437 <= mux_166_nl AND and_dcpl_91;
  or_458_cse <= (result_rem_11cyc_st_5(1)) OR (result_rem_11cyc_st_5(0)) OR (result_rem_11cyc_st_5(3));
  and_790_cse <= (result_rem_11cyc_st_5(2)) AND asn_itm_5 AND main_stage_0_6;
  nor_527_nl <= NOT(and_790_cse OR and_dcpl_91);
  or_460_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_79);
  mux_tmp_167 <= MUX_s_1_2_2(nor_527_nl, or_460_nl, or_458_cse);
  nor_528_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_167));
  mux_tmp_168 <= MUX_s_1_2_2(nor_528_nl, mux_tmp_167, or_445_cse);
  nor_529_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_168));
  mux_tmp_169 <= MUX_s_1_2_2(nor_529_nl, mux_tmp_168, or_434_cse);
  nor_530_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_169));
  mux_tmp_170 <= MUX_s_1_2_2(nor_530_nl, mux_tmp_169, or_425_cse);
  nor_531_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_170));
  mux_tmp_171 <= MUX_s_1_2_2(nor_531_nl, mux_tmp_170, or_418_cse);
  and_789_nl <= nand_144_cse AND mux_tmp_171;
  mux_172_nl <= MUX_s_1_2_2(and_789_nl, mux_tmp_171, or_413_cse);
  and_dcpl_441 <= mux_172_nl AND and_dcpl_65;
  or_473_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0100"));
  nor_522_nl <= NOT(and_dcpl_79 OR and_dcpl_65);
  or_475_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0100")) OR (NOT
      and_dcpl_53);
  mux_tmp_173 <= MUX_s_1_2_2(nor_522_nl, or_475_nl, or_473_cse);
  nand_138_cse <= NOT((result_rem_11cyc_st_5(2)) AND asn_itm_5 AND main_stage_0_6);
  and_788_nl <= nand_138_cse AND mux_tmp_173;
  mux_tmp_174 <= MUX_s_1_2_2(and_788_nl, mux_tmp_173, or_458_cse);
  nor_523_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_174));
  mux_tmp_175 <= MUX_s_1_2_2(nor_523_nl, mux_tmp_174, or_445_cse);
  nor_524_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_175));
  mux_tmp_176 <= MUX_s_1_2_2(nor_524_nl, mux_tmp_175, or_434_cse);
  nor_525_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_176));
  mux_tmp_177 <= MUX_s_1_2_2(nor_525_nl, mux_tmp_176, or_425_cse);
  nor_526_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_177));
  mux_tmp_178 <= MUX_s_1_2_2(nor_526_nl, mux_tmp_177, or_418_cse);
  and_787_nl <= nand_144_cse AND mux_tmp_178;
  mux_179_nl <= MUX_s_1_2_2(and_787_nl, mux_tmp_178, or_413_cse);
  and_dcpl_444 <= mux_179_nl AND and_dcpl_39;
  nor_516_nl <= NOT(and_dcpl_53 OR and_dcpl_39);
  or_492_nl <= (result_rem_11cyc_st_8(0)) OR (result_rem_11cyc_st_8(1)) OR (result_rem_11cyc_st_8(3))
      OR (NOT and_dcpl_38);
  or_490_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0100"));
  mux_tmp_180 <= MUX_s_1_2_2(nor_516_nl, or_492_nl, or_490_nl);
  nor_517_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_180));
  mux_tmp_181 <= MUX_s_1_2_2(nor_517_nl, mux_tmp_180, or_473_cse);
  and_785_nl <= nand_138_cse AND mux_tmp_181;
  mux_tmp_182 <= MUX_s_1_2_2(and_785_nl, mux_tmp_181, or_458_cse);
  nor_518_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_182));
  mux_tmp_183 <= MUX_s_1_2_2(nor_518_nl, mux_tmp_182, or_445_cse);
  nor_519_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_183));
  mux_tmp_184 <= MUX_s_1_2_2(nor_519_nl, mux_tmp_183, or_434_cse);
  nor_520_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_184));
  mux_tmp_185 <= MUX_s_1_2_2(nor_520_nl, mux_tmp_184, or_425_cse);
  nor_521_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_185));
  mux_tmp_186 <= MUX_s_1_2_2(nor_521_nl, mux_tmp_185, or_418_cse);
  and_786_nl <= nand_144_cse AND mux_tmp_186;
  mux_187_nl <= MUX_s_1_2_2(and_786_nl, mux_tmp_186, or_413_cse);
  and_dcpl_447 <= mux_187_nl AND and_dcpl_13 AND and_dcpl_2;
  and_tmp_34 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0100")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0100")));
  nor_514_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_34));
  mux_tmp_188 <= MUX_s_1_2_2(nor_514_nl, and_tmp_34, or_418_cse);
  nor_515_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_188));
  or_501_nl <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0100"));
  mux_tmp_189 <= MUX_s_1_2_2(nor_515_nl, mux_tmp_188, or_501_nl);
  and_dcpl_452 <= and_dcpl_417 AND and_dcpl_318;
  or_tmp_502 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_208);
  or_516_cse <= (result_result_acc_tmp(1)) OR (NOT (result_result_acc_tmp(0))) OR
      (result_result_acc_tmp(3));
  and_784_nl <= nand_144_cse AND or_tmp_502;
  mux_190_nl <= MUX_s_1_2_2(and_784_nl, or_tmp_502, or_516_cse);
  and_dcpl_455 <= mux_190_nl AND and_dcpl_196;
  or_521_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0101"));
  nor_513_nl <= NOT(and_dcpl_208 OR and_dcpl_196);
  or_523_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_182);
  mux_tmp_191 <= MUX_s_1_2_2(nor_513_nl, or_523_nl, or_521_cse);
  and_783_nl <= nand_144_cse AND mux_tmp_191;
  mux_192_nl <= MUX_s_1_2_2(and_783_nl, mux_tmp_191, or_516_cse);
  and_dcpl_458 <= mux_192_nl AND and_dcpl_170;
  or_528_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0101"));
  nor_511_nl <= NOT(and_dcpl_182 OR and_dcpl_170);
  or_530_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_156);
  mux_tmp_193 <= MUX_s_1_2_2(nor_511_nl, or_530_nl, or_528_cse);
  nor_512_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_193));
  mux_tmp_194 <= MUX_s_1_2_2(nor_512_nl, mux_tmp_193, or_521_cse);
  and_782_nl <= nand_144_cse AND mux_tmp_194;
  mux_195_nl <= MUX_s_1_2_2(and_782_nl, mux_tmp_194, or_516_cse);
  and_dcpl_462 <= mux_195_nl AND and_dcpl_145;
  or_537_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0101"));
  nor_508_nl <= NOT(and_dcpl_156 OR and_dcpl_145);
  or_539_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_130);
  mux_tmp_196 <= MUX_s_1_2_2(nor_508_nl, or_539_nl, or_537_cse);
  nor_509_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_196));
  mux_tmp_197 <= MUX_s_1_2_2(nor_509_nl, mux_tmp_196, or_528_cse);
  nor_510_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_197));
  mux_tmp_198 <= MUX_s_1_2_2(nor_510_nl, mux_tmp_197, or_521_cse);
  and_781_nl <= nand_144_cse AND mux_tmp_198;
  mux_199_nl <= MUX_s_1_2_2(and_781_nl, mux_tmp_198, or_516_cse);
  and_dcpl_464 <= mux_199_nl AND and_dcpl_117;
  or_548_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0101"));
  nor_504_nl <= NOT(and_dcpl_130 OR and_dcpl_117);
  or_550_nl <= (result_rem_11cyc_st_5(1)) OR (NOT (result_rem_11cyc_st_5(0))) OR
      (result_rem_11cyc_st_5(3)) OR (NOT and_dcpl_115);
  mux_tmp_200 <= MUX_s_1_2_2(nor_504_nl, or_550_nl, or_548_cse);
  nor_505_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_200));
  mux_tmp_201 <= MUX_s_1_2_2(nor_505_nl, mux_tmp_200, or_537_cse);
  nor_506_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_201));
  mux_tmp_202 <= MUX_s_1_2_2(nor_506_nl, mux_tmp_201, or_528_cse);
  nor_507_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_202));
  mux_tmp_203 <= MUX_s_1_2_2(nor_507_nl, mux_tmp_202, or_521_cse);
  and_780_nl <= nand_144_cse AND mux_tmp_203;
  mux_204_nl <= MUX_s_1_2_2(and_780_nl, mux_tmp_203, or_516_cse);
  and_dcpl_468 <= mux_204_nl AND and_dcpl_94;
  or_561_cse <= (result_rem_11cyc_st_5(1)) OR (NOT (result_rem_11cyc_st_5(0))) OR
      (result_rem_11cyc_st_5(3));
  nor_499_nl <= NOT(and_790_cse OR and_dcpl_94);
  or_563_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_79);
  mux_tmp_205 <= MUX_s_1_2_2(nor_499_nl, or_563_nl, or_561_cse);
  nor_500_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_205));
  mux_tmp_206 <= MUX_s_1_2_2(nor_500_nl, mux_tmp_205, or_548_cse);
  nor_501_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_206));
  mux_tmp_207 <= MUX_s_1_2_2(nor_501_nl, mux_tmp_206, or_537_cse);
  nor_502_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_207));
  mux_tmp_208 <= MUX_s_1_2_2(nor_502_nl, mux_tmp_207, or_528_cse);
  nor_503_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_208));
  mux_tmp_209 <= MUX_s_1_2_2(nor_503_nl, mux_tmp_208, or_521_cse);
  and_778_nl <= nand_144_cse AND mux_tmp_209;
  mux_210_nl <= MUX_s_1_2_2(and_778_nl, mux_tmp_209, or_516_cse);
  and_dcpl_472 <= mux_210_nl AND and_dcpl_68;
  or_576_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0101"));
  nor_494_nl <= NOT(and_dcpl_79 OR and_dcpl_68);
  or_578_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      and_dcpl_53);
  mux_tmp_211 <= MUX_s_1_2_2(nor_494_nl, or_578_nl, or_576_cse);
  and_777_nl <= nand_138_cse AND mux_tmp_211;
  mux_tmp_212 <= MUX_s_1_2_2(and_777_nl, mux_tmp_211, or_561_cse);
  nor_495_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_212));
  mux_tmp_213 <= MUX_s_1_2_2(nor_495_nl, mux_tmp_212, or_548_cse);
  nor_496_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_213));
  mux_tmp_214 <= MUX_s_1_2_2(nor_496_nl, mux_tmp_213, or_537_cse);
  nor_497_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_214));
  mux_tmp_215 <= MUX_s_1_2_2(nor_497_nl, mux_tmp_214, or_528_cse);
  nor_498_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_215));
  mux_tmp_216 <= MUX_s_1_2_2(nor_498_nl, mux_tmp_215, or_521_cse);
  and_776_nl <= nand_144_cse AND mux_tmp_216;
  mux_217_nl <= MUX_s_1_2_2(and_776_nl, mux_tmp_216, or_516_cse);
  and_dcpl_474 <= mux_217_nl AND and_dcpl_40;
  nor_488_nl <= NOT(and_dcpl_53 OR and_dcpl_40);
  or_595_nl <= (NOT (result_rem_11cyc_st_8(0))) OR (result_rem_11cyc_st_8(1)) OR
      (result_rem_11cyc_st_8(3)) OR (NOT and_dcpl_38);
  or_593_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0101"));
  mux_tmp_218 <= MUX_s_1_2_2(nor_488_nl, or_595_nl, or_593_nl);
  nor_489_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_218));
  mux_tmp_219 <= MUX_s_1_2_2(nor_489_nl, mux_tmp_218, or_576_cse);
  and_774_nl <= nand_138_cse AND mux_tmp_219;
  mux_tmp_220 <= MUX_s_1_2_2(and_774_nl, mux_tmp_219, or_561_cse);
  nor_490_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_220));
  mux_tmp_221 <= MUX_s_1_2_2(nor_490_nl, mux_tmp_220, or_548_cse);
  nor_491_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_221));
  mux_tmp_222 <= MUX_s_1_2_2(nor_491_nl, mux_tmp_221, or_537_cse);
  nor_492_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_222));
  mux_tmp_223 <= MUX_s_1_2_2(nor_492_nl, mux_tmp_222, or_528_cse);
  nor_493_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_223));
  mux_tmp_224 <= MUX_s_1_2_2(nor_493_nl, mux_tmp_223, or_521_cse);
  and_775_nl <= nand_144_cse AND mux_tmp_224;
  mux_225_nl <= MUX_s_1_2_2(and_775_nl, mux_tmp_224, or_516_cse);
  and_dcpl_476 <= mux_225_nl AND and_dcpl_13 AND and_dcpl_6;
  and_tmp_41 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0101")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0101")));
  nor_487_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_41));
  mux_tmp_226 <= MUX_s_1_2_2(nor_487_nl, and_tmp_41, or_521_cse);
  and_773_nl <= nand_146_cse AND mux_tmp_226;
  or_604_nl <= CONV_SL_1_1(result_result_acc_tmp(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_227 <= MUX_s_1_2_2(and_773_nl, mux_tmp_226, or_604_nl);
  and_dcpl_480 <= and_dcpl_417 AND and_dcpl_352;
  or_tmp_602 <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_208);
  or_617_cse <= (NOT (result_result_acc_tmp(1))) OR (result_result_acc_tmp(0)) OR
      (result_result_acc_tmp(3));
  and_772_nl <= nand_144_cse AND or_tmp_602;
  mux_228_nl <= MUX_s_1_2_2(and_772_nl, or_tmp_602, or_617_cse);
  and_dcpl_484 <= mux_228_nl AND and_dcpl_199;
  or_622_cse <= CONV_SL_1_1(result_rem_11cyc/=STD_LOGIC_VECTOR'("0110"));
  nor_486_nl <= NOT(and_dcpl_208 OR and_dcpl_199);
  or_624_nl <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_182);
  mux_tmp_229 <= MUX_s_1_2_2(nor_486_nl, or_624_nl, or_622_cse);
  and_771_nl <= nand_144_cse AND mux_tmp_229;
  mux_230_nl <= MUX_s_1_2_2(and_771_nl, mux_tmp_229, or_617_cse);
  and_dcpl_488 <= mux_230_nl AND and_dcpl_173;
  or_629_cse <= CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0110"));
  nor_484_nl <= NOT(and_dcpl_182 OR and_dcpl_173);
  or_631_nl <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_156);
  mux_tmp_231 <= MUX_s_1_2_2(nor_484_nl, or_631_nl, or_629_cse);
  nor_485_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_231));
  mux_tmp_232 <= MUX_s_1_2_2(nor_485_nl, mux_tmp_231, or_622_cse);
  and_770_nl <= nand_144_cse AND mux_tmp_232;
  mux_233_nl <= MUX_s_1_2_2(and_770_nl, mux_tmp_232, or_617_cse);
  and_dcpl_491 <= mux_233_nl AND and_dcpl_147;
  or_638_cse <= CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0110"));
  nor_481_nl <= NOT(and_dcpl_156 OR and_dcpl_147);
  or_640_nl <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_130);
  mux_tmp_234 <= MUX_s_1_2_2(nor_481_nl, or_640_nl, or_638_cse);
  nor_482_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_234));
  mux_tmp_235 <= MUX_s_1_2_2(nor_482_nl, mux_tmp_234, or_629_cse);
  nor_483_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_235));
  mux_tmp_236 <= MUX_s_1_2_2(nor_483_nl, mux_tmp_235, or_622_cse);
  and_769_nl <= nand_144_cse AND mux_tmp_236;
  mux_237_nl <= MUX_s_1_2_2(and_769_nl, mux_tmp_236, or_617_cse);
  and_dcpl_493 <= mux_237_nl AND and_dcpl_118;
  or_649_cse <= CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0110"));
  nor_477_nl <= NOT(and_dcpl_130 OR and_dcpl_118);
  or_651_nl <= (NOT (result_rem_11cyc_st_5(1))) OR (result_rem_11cyc_st_5(0)) OR
      (result_rem_11cyc_st_5(3)) OR (NOT and_dcpl_115);
  mux_tmp_238 <= MUX_s_1_2_2(nor_477_nl, or_651_nl, or_649_cse);
  nor_478_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_238));
  mux_tmp_239 <= MUX_s_1_2_2(nor_478_nl, mux_tmp_238, or_638_cse);
  nor_479_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_239));
  mux_tmp_240 <= MUX_s_1_2_2(nor_479_nl, mux_tmp_239, or_629_cse);
  nor_480_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_240));
  mux_tmp_241 <= MUX_s_1_2_2(nor_480_nl, mux_tmp_240, or_622_cse);
  and_768_nl <= nand_144_cse AND mux_tmp_241;
  mux_242_nl <= MUX_s_1_2_2(and_768_nl, mux_tmp_241, or_617_cse);
  and_dcpl_496 <= mux_242_nl AND and_dcpl_96;
  or_662_cse <= (NOT (result_rem_11cyc_st_5(1))) OR (result_rem_11cyc_st_5(0)) OR
      (result_rem_11cyc_st_5(3));
  nor_472_nl <= NOT(and_790_cse OR and_dcpl_96);
  or_664_nl <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_79);
  mux_tmp_243 <= MUX_s_1_2_2(nor_472_nl, or_664_nl, or_662_cse);
  nor_473_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_243));
  mux_tmp_244 <= MUX_s_1_2_2(nor_473_nl, mux_tmp_243, or_649_cse);
  nor_474_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_244));
  mux_tmp_245 <= MUX_s_1_2_2(nor_474_nl, mux_tmp_244, or_638_cse);
  nor_475_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_245));
  mux_tmp_246 <= MUX_s_1_2_2(nor_475_nl, mux_tmp_245, or_629_cse);
  nor_476_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_246));
  mux_tmp_247 <= MUX_s_1_2_2(nor_476_nl, mux_tmp_246, or_622_cse);
  and_766_nl <= nand_144_cse AND mux_tmp_247;
  mux_248_nl <= MUX_s_1_2_2(and_766_nl, mux_tmp_247, or_617_cse);
  and_dcpl_499 <= mux_248_nl AND and_dcpl_70;
  or_677_cse <= CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0110"));
  nor_467_nl <= NOT(and_dcpl_79 OR and_dcpl_70);
  or_679_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      and_dcpl_53);
  mux_tmp_249 <= MUX_s_1_2_2(nor_467_nl, or_679_nl, or_677_cse);
  and_765_nl <= nand_138_cse AND mux_tmp_249;
  mux_tmp_250 <= MUX_s_1_2_2(and_765_nl, mux_tmp_249, or_662_cse);
  nor_468_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_250));
  mux_tmp_251 <= MUX_s_1_2_2(nor_468_nl, mux_tmp_250, or_649_cse);
  nor_469_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_251));
  mux_tmp_252 <= MUX_s_1_2_2(nor_469_nl, mux_tmp_251, or_638_cse);
  nor_470_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_252));
  mux_tmp_253 <= MUX_s_1_2_2(nor_470_nl, mux_tmp_252, or_629_cse);
  nor_471_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_253));
  mux_tmp_254 <= MUX_s_1_2_2(nor_471_nl, mux_tmp_253, or_622_cse);
  and_764_nl <= nand_144_cse AND mux_tmp_254;
  mux_255_nl <= MUX_s_1_2_2(and_764_nl, mux_tmp_254, or_617_cse);
  and_dcpl_501 <= mux_255_nl AND and_dcpl_41;
  nor_461_nl <= NOT(and_dcpl_53 OR and_dcpl_41);
  or_696_nl <= (result_rem_11cyc_st_8(0)) OR (NOT (result_rem_11cyc_st_8(1))) OR
      (result_rem_11cyc_st_8(3)) OR (NOT and_dcpl_38);
  or_694_nl <= CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0110"));
  mux_tmp_256 <= MUX_s_1_2_2(nor_461_nl, or_696_nl, or_694_nl);
  nor_462_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_256));
  mux_tmp_257 <= MUX_s_1_2_2(nor_462_nl, mux_tmp_256, or_677_cse);
  and_762_nl <= nand_138_cse AND mux_tmp_257;
  mux_tmp_258 <= MUX_s_1_2_2(and_762_nl, mux_tmp_257, or_662_cse);
  nor_463_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_258));
  mux_tmp_259 <= MUX_s_1_2_2(nor_463_nl, mux_tmp_258, or_649_cse);
  nor_464_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_259));
  mux_tmp_260 <= MUX_s_1_2_2(nor_464_nl, mux_tmp_259, or_638_cse);
  nor_465_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_260));
  mux_tmp_261 <= MUX_s_1_2_2(nor_465_nl, mux_tmp_260, or_629_cse);
  nor_466_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_261));
  mux_tmp_262 <= MUX_s_1_2_2(nor_466_nl, mux_tmp_261, or_622_cse);
  and_763_nl <= nand_144_cse AND mux_tmp_262;
  mux_263_nl <= MUX_s_1_2_2(and_763_nl, mux_tmp_262, or_617_cse);
  and_dcpl_503 <= mux_263_nl AND and_dcpl_13 AND and_dcpl_9;
  and_tmp_48 <= ((NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("0110")))
      AND ((NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("0110")));
  nor_459_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_48));
  mux_tmp_264 <= MUX_s_1_2_2(nor_459_nl, and_tmp_48, or_622_cse);
  nor_460_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_264));
  or_705_nl <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("0110"));
  mux_tmp_265 <= MUX_s_1_2_2(nor_460_nl, mux_tmp_264, or_705_nl);
  and_dcpl_507 <= and_dcpl_417 AND and_dcpl_386;
  or_tmp_702 <= NOT(CONV_SL_1_1(result_rem_11cyc=STD_LOGIC_VECTOR'("0111")) AND and_dcpl_208);
  or_718_cse <= (NOT (result_result_acc_tmp(1))) OR (NOT (result_result_acc_tmp(0)))
      OR (result_result_acc_tmp(3));
  and_761_nl <= nand_144_cse AND or_tmp_702;
  mux_266_nl <= MUX_s_1_2_2(and_761_nl, or_tmp_702, or_718_cse);
  and_dcpl_510 <= mux_266_nl AND and_dcpl_201;
  nand_112_cse <= NOT(CONV_SL_1_1(result_rem_11cyc=STD_LOGIC_VECTOR'("0111")));
  nor_458_nl <= NOT(and_dcpl_208 OR and_dcpl_201);
  nand_153_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_2=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_182);
  mux_tmp_267 <= MUX_s_1_2_2(nor_458_nl, nand_153_nl, nand_112_cse);
  and_760_nl <= nand_144_cse AND mux_tmp_267;
  mux_268_nl <= MUX_s_1_2_2(and_760_nl, mux_tmp_267, or_718_cse);
  and_dcpl_513 <= mux_268_nl AND and_dcpl_175;
  nand_108_cse <= NOT(CONV_SL_1_1(result_rem_11cyc_st_2=STD_LOGIC_VECTOR'("0111")));
  nor_456_nl <= NOT(and_dcpl_182 OR and_dcpl_175);
  nand_152_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_3=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_156);
  mux_tmp_269 <= MUX_s_1_2_2(nor_456_nl, nand_152_nl, nand_108_cse);
  nor_457_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_269));
  mux_tmp_270 <= MUX_s_1_2_2(nor_457_nl, mux_tmp_269, nand_112_cse);
  and_759_nl <= nand_144_cse AND mux_tmp_270;
  mux_271_nl <= MUX_s_1_2_2(and_759_nl, mux_tmp_270, or_718_cse);
  and_dcpl_516 <= mux_271_nl AND and_dcpl_149;
  nand_103_cse <= NOT(CONV_SL_1_1(result_rem_11cyc_st_3=STD_LOGIC_VECTOR'("0111")));
  nor_453_nl <= NOT(and_dcpl_156 OR and_dcpl_149);
  nand_151_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_4=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_130);
  mux_tmp_272 <= MUX_s_1_2_2(nor_453_nl, nand_151_nl, nand_103_cse);
  nor_454_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_272));
  mux_tmp_273 <= MUX_s_1_2_2(nor_454_nl, mux_tmp_272, nand_108_cse);
  nor_455_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_273));
  mux_tmp_274 <= MUX_s_1_2_2(nor_455_nl, mux_tmp_273, nand_112_cse);
  and_758_nl <= nand_144_cse AND mux_tmp_274;
  mux_275_nl <= MUX_s_1_2_2(and_758_nl, mux_tmp_274, or_718_cse);
  and_dcpl_518 <= mux_275_nl AND and_dcpl_119;
  nand_97_cse <= NOT(CONV_SL_1_1(result_rem_11cyc_st_4=STD_LOGIC_VECTOR'("0111")));
  nor_449_nl <= NOT(and_dcpl_130 OR and_dcpl_119);
  nand_96_nl <= NOT((result_rem_11cyc_st_5(1)) AND (result_rem_11cyc_st_5(0)) AND
      (NOT (result_rem_11cyc_st_5(3))) AND and_dcpl_115);
  mux_tmp_276 <= MUX_s_1_2_2(nor_449_nl, nand_96_nl, nand_97_cse);
  nor_450_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_276));
  mux_tmp_277 <= MUX_s_1_2_2(nor_450_nl, mux_tmp_276, nand_103_cse);
  nor_451_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_277));
  mux_tmp_278 <= MUX_s_1_2_2(nor_451_nl, mux_tmp_277, nand_108_cse);
  nor_452_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_278));
  mux_tmp_279 <= MUX_s_1_2_2(nor_452_nl, mux_tmp_278, nand_112_cse);
  and_757_nl <= nand_144_cse AND mux_tmp_279;
  mux_280_nl <= MUX_s_1_2_2(and_757_nl, mux_tmp_279, or_718_cse);
  and_dcpl_521 <= mux_280_nl AND and_dcpl_98;
  or_763_cse <= (NOT (result_rem_11cyc_st_5(1))) OR (NOT (result_rem_11cyc_st_5(0)))
      OR (result_rem_11cyc_st_5(3));
  nor_444_nl <= NOT(and_790_cse OR and_dcpl_98);
  nand_150_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_6=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_79);
  mux_tmp_281 <= MUX_s_1_2_2(nor_444_nl, nand_150_nl, or_763_cse);
  nor_445_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_281));
  mux_tmp_282 <= MUX_s_1_2_2(nor_445_nl, mux_tmp_281, nand_97_cse);
  nor_446_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_282));
  mux_tmp_283 <= MUX_s_1_2_2(nor_446_nl, mux_tmp_282, nand_103_cse);
  nor_447_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_283));
  mux_tmp_284 <= MUX_s_1_2_2(nor_447_nl, mux_tmp_283, nand_108_cse);
  nor_448_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_284));
  mux_tmp_285 <= MUX_s_1_2_2(nor_448_nl, mux_tmp_284, nand_112_cse);
  and_755_nl <= nand_144_cse AND mux_tmp_285;
  mux_286_nl <= MUX_s_1_2_2(and_755_nl, mux_tmp_285, or_718_cse);
  and_dcpl_524 <= mux_286_nl AND and_dcpl_72;
  nand_83_cse <= NOT(CONV_SL_1_1(result_rem_11cyc_st_6=STD_LOGIC_VECTOR'("0111")));
  nor_439_nl <= NOT(and_dcpl_79 OR and_dcpl_72);
  nand_149_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_7=STD_LOGIC_VECTOR'("0111"))
      AND and_dcpl_53);
  mux_tmp_287 <= MUX_s_1_2_2(nor_439_nl, nand_149_nl, nand_83_cse);
  and_754_nl <= nand_138_cse AND mux_tmp_287;
  mux_tmp_288 <= MUX_s_1_2_2(and_754_nl, mux_tmp_287, or_763_cse);
  nor_440_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_288));
  mux_tmp_289 <= MUX_s_1_2_2(nor_440_nl, mux_tmp_288, nand_97_cse);
  nor_441_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_289));
  mux_tmp_290 <= MUX_s_1_2_2(nor_441_nl, mux_tmp_289, nand_103_cse);
  nor_442_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_290));
  mux_tmp_291 <= MUX_s_1_2_2(nor_442_nl, mux_tmp_290, nand_108_cse);
  nor_443_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_291));
  mux_tmp_292 <= MUX_s_1_2_2(nor_443_nl, mux_tmp_291, nand_112_cse);
  and_753_nl <= nand_144_cse AND mux_tmp_292;
  mux_293_nl <= MUX_s_1_2_2(and_753_nl, mux_tmp_292, or_718_cse);
  and_dcpl_526 <= mux_293_nl AND and_dcpl_42;
  nor_433_nl <= NOT(and_dcpl_53 OR and_dcpl_42);
  nand_72_nl <= NOT((result_rem_11cyc_st_8(0)) AND (result_rem_11cyc_st_8(1)) AND
      (NOT (result_rem_11cyc_st_8(3))) AND and_dcpl_38);
  nand_73_nl <= NOT(CONV_SL_1_1(result_rem_11cyc_st_7=STD_LOGIC_VECTOR'("0111")));
  mux_tmp_294 <= MUX_s_1_2_2(nor_433_nl, nand_72_nl, nand_73_nl);
  nor_434_nl <= NOT(and_dcpl_79 OR (NOT mux_tmp_294));
  mux_tmp_295 <= MUX_s_1_2_2(nor_434_nl, mux_tmp_294, nand_83_cse);
  and_751_nl <= nand_138_cse AND mux_tmp_295;
  mux_tmp_296 <= MUX_s_1_2_2(and_751_nl, mux_tmp_295, or_763_cse);
  nor_435_nl <= NOT(and_dcpl_130 OR (NOT mux_tmp_296));
  mux_tmp_297 <= MUX_s_1_2_2(nor_435_nl, mux_tmp_296, nand_97_cse);
  nor_436_nl <= NOT(and_dcpl_156 OR (NOT mux_tmp_297));
  mux_tmp_298 <= MUX_s_1_2_2(nor_436_nl, mux_tmp_297, nand_103_cse);
  nor_437_nl <= NOT(and_dcpl_182 OR (NOT mux_tmp_298));
  mux_tmp_299 <= MUX_s_1_2_2(nor_437_nl, mux_tmp_298, nand_108_cse);
  nor_438_nl <= NOT(and_dcpl_208 OR (NOT mux_tmp_299));
  mux_tmp_300 <= MUX_s_1_2_2(nor_438_nl, mux_tmp_299, nand_112_cse);
  and_752_nl <= nand_144_cse AND mux_tmp_300;
  mux_301_nl <= MUX_s_1_2_2(and_752_nl, mux_tmp_300, or_718_cse);
  and_dcpl_528 <= mux_301_nl AND and_dcpl_13 AND and_dcpl_11;
  and_tmp_55 <= (NOT(main_stage_0_3 AND asn_itm_2 AND CONV_SL_1_1(result_rem_11cyc_st_2=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_4 AND asn_itm_3 AND CONV_SL_1_1(result_rem_11cyc_st_3=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_5 AND asn_itm_4 AND CONV_SL_1_1(result_rem_11cyc_st_4=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_6 AND asn_itm_5 AND CONV_SL_1_1(result_rem_11cyc_st_5=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_7 AND asn_itm_6 AND CONV_SL_1_1(result_rem_11cyc_st_6=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_8 AND asn_itm_7 AND CONV_SL_1_1(result_rem_11cyc_st_7=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_9 AND asn_itm_8 AND CONV_SL_1_1(result_rem_11cyc_st_8=STD_LOGIC_VECTOR'("0111"))))
      AND (NOT(main_stage_0_10 AND asn_itm_9 AND CONV_SL_1_1(result_rem_11cyc_st_9=STD_LOGIC_VECTOR'("0111"))));
  nor_432_nl <= NOT(and_dcpl_208 OR (NOT and_tmp_55));
  mux_tmp_302 <= MUX_s_1_2_2(nor_432_nl, and_tmp_55, nand_112_cse);
  and_750_nl <= (NOT(CONV_SL_1_1(result_result_acc_tmp(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND ccs_ccore_start_rsci_idat)) AND mux_tmp_302;
  mux_tmp_303 <= MUX_s_1_2_2(and_750_nl, mux_tmp_302, result_result_acc_tmp(3));
  and_dcpl_532 <= and_dcpl_261 AND (result_result_acc_tmp(3));
  and_dcpl_533 <= and_dcpl_532 AND and_dcpl_260;
  not_tmp_645 <= NOT((result_rem_11cyc(3)) AND asn_itm_1 AND main_stage_0_2);
  or_tmp_801 <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR not_tmp_645;
  or_818_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("1000"));
  nor_431_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_801));
  mux_304_nl <= MUX_s_1_2_2(nor_431_nl, or_tmp_801, or_818_cse);
  and_dcpl_536 <= mux_304_nl AND and_dcpl_203;
  or_823_cse <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_749_cse <= (result_rem_11cyc(3)) AND asn_itm_1 AND main_stage_0_2;
  nor_430_nl <= NOT(and_749_cse OR and_dcpl_203);
  or_825_nl <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_202);
  mux_tmp_305 <= MUX_s_1_2_2(nor_430_nl, or_825_nl, or_823_cse);
  nor_429_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_305));
  mux_306_nl <= MUX_s_1_2_2(nor_429_nl, mux_tmp_305, or_818_cse);
  and_dcpl_539 <= mux_306_nl AND and_dcpl_177;
  or_830_cse <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_747_cse <= (result_rem_11cyc_st_2(3)) AND asn_itm_2 AND main_stage_0_3;
  nor_428_nl <= NOT(and_747_cse OR and_dcpl_177);
  or_832_nl <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_176);
  mux_tmp_307 <= MUX_s_1_2_2(nor_428_nl, or_832_nl, or_830_cse);
  and_748_nl <= not_tmp_645 AND mux_tmp_307;
  mux_tmp_308 <= MUX_s_1_2_2(and_748_nl, mux_tmp_307, or_823_cse);
  nor_427_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_308));
  mux_309_nl <= MUX_s_1_2_2(nor_427_nl, mux_tmp_308, or_818_cse);
  and_dcpl_542 <= mux_309_nl AND and_dcpl_151;
  or_839_cse <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_744_cse <= (result_rem_11cyc_st_3(3)) AND asn_itm_3 AND main_stage_0_4;
  nor_426_nl <= NOT(and_744_cse OR and_dcpl_151);
  or_841_nl <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_150);
  mux_tmp_310 <= MUX_s_1_2_2(nor_426_nl, or_841_nl, or_839_cse);
  nand_58_cse <= NOT((result_rem_11cyc_st_2(3)) AND asn_itm_2 AND main_stage_0_3);
  and_745_nl <= nand_58_cse AND mux_tmp_310;
  mux_tmp_311 <= MUX_s_1_2_2(and_745_nl, mux_tmp_310, or_830_cse);
  and_746_nl <= not_tmp_645 AND mux_tmp_311;
  mux_tmp_312 <= MUX_s_1_2_2(and_746_nl, mux_tmp_311, or_823_cse);
  nor_425_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_312));
  mux_313_nl <= MUX_s_1_2_2(nor_425_nl, mux_tmp_312, or_818_cse);
  and_dcpl_546 <= mux_313_nl AND and_dcpl_122;
  or_850_cse <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_740_cse <= (result_rem_11cyc_st_4(3)) AND asn_itm_4 AND main_stage_0_5;
  nor_424_nl <= NOT(and_740_cse OR and_dcpl_122);
  or_852_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      and_dcpl_105);
  mux_tmp_314 <= MUX_s_1_2_2(nor_424_nl, or_852_nl, or_850_cse);
  nand_55_cse <= NOT((result_rem_11cyc_st_3(3)) AND asn_itm_3 AND main_stage_0_4);
  and_741_nl <= nand_55_cse AND mux_tmp_314;
  mux_tmp_315 <= MUX_s_1_2_2(and_741_nl, mux_tmp_314, or_839_cse);
  and_742_nl <= nand_58_cse AND mux_tmp_315;
  mux_tmp_316 <= MUX_s_1_2_2(and_742_nl, mux_tmp_315, or_830_cse);
  and_743_nl <= not_tmp_645 AND mux_tmp_316;
  mux_tmp_317 <= MUX_s_1_2_2(and_743_nl, mux_tmp_316, or_823_cse);
  nor_423_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_317));
  mux_318_nl <= MUX_s_1_2_2(nor_423_nl, mux_tmp_317, or_818_cse);
  and_dcpl_549 <= mux_318_nl AND and_dcpl_100;
  or_863_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1000"));
  nor_422_nl <= NOT(and_dcpl_105 OR and_dcpl_100);
  or_865_nl <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_99);
  mux_tmp_319 <= MUX_s_1_2_2(nor_422_nl, or_865_nl, or_863_cse);
  nand_51_cse <= NOT((result_rem_11cyc_st_4(3)) AND asn_itm_4 AND main_stage_0_5);
  and_736_nl <= nand_51_cse AND mux_tmp_319;
  mux_tmp_320 <= MUX_s_1_2_2(and_736_nl, mux_tmp_319, or_850_cse);
  and_737_nl <= nand_55_cse AND mux_tmp_320;
  mux_tmp_321 <= MUX_s_1_2_2(and_737_nl, mux_tmp_320, or_839_cse);
  and_738_nl <= nand_58_cse AND mux_tmp_321;
  mux_tmp_322 <= MUX_s_1_2_2(and_738_nl, mux_tmp_321, or_830_cse);
  and_739_nl <= not_tmp_645 AND mux_tmp_322;
  mux_tmp_323 <= MUX_s_1_2_2(and_739_nl, mux_tmp_322, or_823_cse);
  nor_421_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_323));
  mux_324_nl <= MUX_s_1_2_2(nor_421_nl, mux_tmp_323, or_818_cse);
  and_dcpl_552 <= mux_324_nl AND and_dcpl_74;
  or_878_cse <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  and_731_cse <= (result_rem_11cyc_st_6(3)) AND asn_itm_6 AND main_stage_0_7;
  nor_419_nl <= NOT(and_731_cse OR and_dcpl_74);
  or_880_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT and_dcpl_73);
  mux_tmp_325 <= MUX_s_1_2_2(nor_419_nl, or_880_nl, or_878_cse);
  nor_420_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_325));
  mux_tmp_326 <= MUX_s_1_2_2(nor_420_nl, mux_tmp_325, or_863_cse);
  and_732_nl <= nand_51_cse AND mux_tmp_326;
  mux_tmp_327 <= MUX_s_1_2_2(and_732_nl, mux_tmp_326, or_850_cse);
  and_733_nl <= nand_55_cse AND mux_tmp_327;
  mux_tmp_328 <= MUX_s_1_2_2(and_733_nl, mux_tmp_327, or_839_cse);
  and_734_nl <= nand_58_cse AND mux_tmp_328;
  mux_tmp_329 <= MUX_s_1_2_2(and_734_nl, mux_tmp_328, or_830_cse);
  and_735_nl <= not_tmp_645 AND mux_tmp_329;
  mux_tmp_330 <= MUX_s_1_2_2(and_735_nl, mux_tmp_329, or_823_cse);
  nor_418_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_330));
  mux_331_nl <= MUX_s_1_2_2(nor_418_nl, mux_tmp_330, or_818_cse);
  and_dcpl_556 <= mux_331_nl AND and_dcpl_45;
  and_725_cse <= (result_rem_11cyc_st_7(3)) AND asn_itm_7 AND main_stage_0_8;
  nor_415_nl <= NOT(and_725_cse OR and_dcpl_45);
  or_897_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("1000")) OR (NOT
      and_dcpl_28);
  or_895_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_332 <= MUX_s_1_2_2(nor_415_nl, or_897_nl, or_895_nl);
  nand_42_cse <= NOT((result_rem_11cyc_st_6(3)) AND asn_itm_6 AND main_stage_0_7);
  and_726_nl <= nand_42_cse AND mux_tmp_332;
  mux_tmp_333 <= MUX_s_1_2_2(and_726_nl, mux_tmp_332, or_878_cse);
  nor_416_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_333));
  mux_tmp_334 <= MUX_s_1_2_2(nor_416_nl, mux_tmp_333, or_863_cse);
  and_727_nl <= nand_51_cse AND mux_tmp_334;
  mux_tmp_335 <= MUX_s_1_2_2(and_727_nl, mux_tmp_334, or_850_cse);
  and_728_nl <= nand_55_cse AND mux_tmp_335;
  mux_tmp_336 <= MUX_s_1_2_2(and_728_nl, mux_tmp_335, or_839_cse);
  and_729_nl <= nand_58_cse AND mux_tmp_336;
  mux_tmp_337 <= MUX_s_1_2_2(and_729_nl, mux_tmp_336, or_830_cse);
  and_730_nl <= not_tmp_645 AND mux_tmp_337;
  mux_tmp_338 <= MUX_s_1_2_2(and_730_nl, mux_tmp_337, or_823_cse);
  nor_417_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_338));
  mux_339_nl <= MUX_s_1_2_2(nor_417_nl, mux_tmp_338, or_818_cse);
  and_dcpl_560 <= mux_339_nl AND and_dcpl_4 AND and_dcpl_18 AND (NOT (result_rem_11cyc_st_9(0)));
  or_tmp_897 <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("1000"));
  nor_407_nl <= NOT((result_rem_11cyc_st_8(3)) OR (NOT or_tmp_897));
  or_914_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_340 <= MUX_s_1_2_2(nor_407_nl, or_tmp_897, or_914_nl);
  nor_408_nl <= NOT((result_rem_11cyc_st_7(3)) OR (NOT mux_tmp_340));
  or_913_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_341 <= MUX_s_1_2_2(nor_408_nl, mux_tmp_340, or_913_nl);
  nor_409_nl <= NOT((result_rem_11cyc_st_6(3)) OR (NOT mux_tmp_341));
  or_912_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_342 <= MUX_s_1_2_2(nor_409_nl, mux_tmp_341, or_912_nl);
  nor_410_nl <= NOT((result_rem_11cyc_st_5(3)) OR (NOT mux_tmp_342));
  or_911_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_343 <= MUX_s_1_2_2(nor_410_nl, mux_tmp_342, or_911_nl);
  nor_411_nl <= NOT((result_rem_11cyc_st_4(3)) OR (NOT mux_tmp_343));
  or_910_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_344 <= MUX_s_1_2_2(nor_411_nl, mux_tmp_343, or_910_nl);
  nor_412_nl <= NOT((result_rem_11cyc_st_3(3)) OR (NOT mux_tmp_344));
  or_909_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_345 <= MUX_s_1_2_2(nor_412_nl, mux_tmp_344, or_909_nl);
  nor_413_nl <= NOT((result_rem_11cyc_st_2(3)) OR (NOT mux_tmp_345));
  or_908_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_346 <= MUX_s_1_2_2(nor_413_nl, mux_tmp_345, or_908_nl);
  and_724_nl <= not_tmp_645 AND mux_tmp_346;
  mux_tmp_347 <= MUX_s_1_2_2(and_724_nl, mux_tmp_346, or_823_cse);
  nor_414_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_347));
  mux_tmp_348 <= MUX_s_1_2_2(nor_414_nl, mux_tmp_347, or_818_cse);
  and_dcpl_566 <= and_dcpl_532 AND and_dcpl_318;
  or_tmp_909 <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR not_tmp_645;
  or_928_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("1001"));
  nor_406_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_909));
  mux_349_nl <= MUX_s_1_2_2(nor_406_nl, or_tmp_909, or_928_cse);
  and_dcpl_568 <= mux_349_nl AND and_dcpl_204;
  or_933_cse <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_405_nl <= NOT(and_749_cse OR and_dcpl_204);
  or_935_nl <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_202);
  mux_tmp_350 <= MUX_s_1_2_2(nor_405_nl, or_935_nl, or_933_cse);
  nor_404_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_350));
  mux_351_nl <= MUX_s_1_2_2(nor_404_nl, mux_tmp_350, or_928_cse);
  and_dcpl_570 <= mux_351_nl AND and_dcpl_178;
  or_940_cse <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_403_nl <= NOT(and_747_cse OR and_dcpl_178);
  or_942_nl <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_176);
  mux_tmp_352 <= MUX_s_1_2_2(nor_403_nl, or_942_nl, or_940_cse);
  and_722_nl <= not_tmp_645 AND mux_tmp_352;
  mux_tmp_353 <= MUX_s_1_2_2(and_722_nl, mux_tmp_352, or_933_cse);
  nor_402_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_353));
  mux_354_nl <= MUX_s_1_2_2(nor_402_nl, mux_tmp_353, or_928_cse);
  and_dcpl_572 <= mux_354_nl AND and_dcpl_152;
  or_949_cse <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_401_nl <= NOT(and_744_cse OR and_dcpl_152);
  or_951_nl <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_150);
  mux_tmp_355 <= MUX_s_1_2_2(nor_401_nl, or_951_nl, or_949_cse);
  and_719_nl <= nand_58_cse AND mux_tmp_355;
  mux_tmp_356 <= MUX_s_1_2_2(and_719_nl, mux_tmp_355, or_940_cse);
  and_720_nl <= not_tmp_645 AND mux_tmp_356;
  mux_tmp_357 <= MUX_s_1_2_2(and_720_nl, mux_tmp_356, or_933_cse);
  nor_400_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_357));
  mux_358_nl <= MUX_s_1_2_2(nor_400_nl, mux_tmp_357, or_928_cse);
  and_dcpl_576 <= mux_358_nl AND and_dcpl_125;
  or_960_cse <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_399_nl <= NOT(and_740_cse OR and_dcpl_125);
  or_962_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1001")) OR (NOT
      and_dcpl_105);
  mux_tmp_359 <= MUX_s_1_2_2(nor_399_nl, or_962_nl, or_960_cse);
  and_715_nl <= nand_55_cse AND mux_tmp_359;
  mux_tmp_360 <= MUX_s_1_2_2(and_715_nl, mux_tmp_359, or_949_cse);
  and_716_nl <= nand_58_cse AND mux_tmp_360;
  mux_tmp_361 <= MUX_s_1_2_2(and_716_nl, mux_tmp_360, or_940_cse);
  and_717_nl <= not_tmp_645 AND mux_tmp_361;
  mux_tmp_362 <= MUX_s_1_2_2(and_717_nl, mux_tmp_361, or_933_cse);
  nor_398_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_362));
  mux_363_nl <= MUX_s_1_2_2(nor_398_nl, mux_tmp_362, or_928_cse);
  and_dcpl_578 <= mux_363_nl AND and_dcpl_101;
  or_973_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1001"));
  nor_397_nl <= NOT(and_dcpl_105 OR and_dcpl_101);
  or_975_nl <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_99);
  mux_tmp_364 <= MUX_s_1_2_2(nor_397_nl, or_975_nl, or_973_cse);
  and_710_nl <= nand_51_cse AND mux_tmp_364;
  mux_tmp_365 <= MUX_s_1_2_2(and_710_nl, mux_tmp_364, or_960_cse);
  and_711_nl <= nand_55_cse AND mux_tmp_365;
  mux_tmp_366 <= MUX_s_1_2_2(and_711_nl, mux_tmp_365, or_949_cse);
  and_712_nl <= nand_58_cse AND mux_tmp_366;
  mux_tmp_367 <= MUX_s_1_2_2(and_712_nl, mux_tmp_366, or_940_cse);
  and_713_nl <= not_tmp_645 AND mux_tmp_367;
  mux_tmp_368 <= MUX_s_1_2_2(and_713_nl, mux_tmp_367, or_933_cse);
  nor_396_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_368));
  mux_369_nl <= MUX_s_1_2_2(nor_396_nl, mux_tmp_368, or_928_cse);
  and_dcpl_580 <= mux_369_nl AND and_dcpl_75;
  or_988_cse <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  nor_394_nl <= NOT(and_731_cse OR and_dcpl_75);
  or_990_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT and_dcpl_73);
  mux_tmp_370 <= MUX_s_1_2_2(nor_394_nl, or_990_nl, or_988_cse);
  nor_395_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_370));
  mux_tmp_371 <= MUX_s_1_2_2(nor_395_nl, mux_tmp_370, or_973_cse);
  and_706_nl <= nand_51_cse AND mux_tmp_371;
  mux_tmp_372 <= MUX_s_1_2_2(and_706_nl, mux_tmp_371, or_960_cse);
  and_707_nl <= nand_55_cse AND mux_tmp_372;
  mux_tmp_373 <= MUX_s_1_2_2(and_707_nl, mux_tmp_372, or_949_cse);
  and_708_nl <= nand_58_cse AND mux_tmp_373;
  mux_tmp_374 <= MUX_s_1_2_2(and_708_nl, mux_tmp_373, or_940_cse);
  and_709_nl <= not_tmp_645 AND mux_tmp_374;
  mux_tmp_375 <= MUX_s_1_2_2(and_709_nl, mux_tmp_374, or_933_cse);
  nor_393_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_375));
  mux_376_nl <= MUX_s_1_2_2(nor_393_nl, mux_tmp_375, or_928_cse);
  and_dcpl_583 <= mux_376_nl AND and_dcpl_47;
  nor_390_nl <= NOT(and_725_cse OR and_dcpl_47);
  or_1007_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("1001")) OR
      (NOT and_dcpl_28);
  or_1005_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_377 <= MUX_s_1_2_2(nor_390_nl, or_1007_nl, or_1005_nl);
  and_700_nl <= nand_42_cse AND mux_tmp_377;
  mux_tmp_378 <= MUX_s_1_2_2(and_700_nl, mux_tmp_377, or_988_cse);
  nor_391_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_378));
  mux_tmp_379 <= MUX_s_1_2_2(nor_391_nl, mux_tmp_378, or_973_cse);
  and_701_nl <= nand_51_cse AND mux_tmp_379;
  mux_tmp_380 <= MUX_s_1_2_2(and_701_nl, mux_tmp_379, or_960_cse);
  and_702_nl <= nand_55_cse AND mux_tmp_380;
  mux_tmp_381 <= MUX_s_1_2_2(and_702_nl, mux_tmp_380, or_949_cse);
  and_703_nl <= nand_58_cse AND mux_tmp_381;
  mux_tmp_382 <= MUX_s_1_2_2(and_703_nl, mux_tmp_381, or_940_cse);
  and_704_nl <= not_tmp_645 AND mux_tmp_382;
  mux_tmp_383 <= MUX_s_1_2_2(and_704_nl, mux_tmp_382, or_933_cse);
  nor_392_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_383));
  mux_384_nl <= MUX_s_1_2_2(nor_392_nl, mux_tmp_383, or_928_cse);
  and_dcpl_586 <= mux_384_nl AND and_dcpl_4 AND and_dcpl_18 AND (result_rem_11cyc_st_9(0));
  or_tmp_1005 <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("1001"));
  nor_383_nl <= NOT((result_rem_11cyc_st_8(3)) OR (NOT or_tmp_1005));
  or_1024_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_385 <= MUX_s_1_2_2(nor_383_nl, or_tmp_1005, or_1024_nl);
  nor_384_nl <= NOT((result_rem_11cyc_st_7(3)) OR (NOT mux_tmp_385));
  or_1023_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_386 <= MUX_s_1_2_2(nor_384_nl, mux_tmp_385, or_1023_nl);
  nor_385_nl <= NOT((result_rem_11cyc_st_6(3)) OR (NOT mux_tmp_386));
  or_1022_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_387 <= MUX_s_1_2_2(nor_385_nl, mux_tmp_386, or_1022_nl);
  nor_386_nl <= NOT((result_rem_11cyc_st_5(3)) OR (NOT mux_tmp_387));
  or_1021_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_388 <= MUX_s_1_2_2(nor_386_nl, mux_tmp_387, or_1021_nl);
  nor_387_nl <= NOT((result_rem_11cyc_st_4(3)) OR (NOT mux_tmp_388));
  or_1020_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_389 <= MUX_s_1_2_2(nor_387_nl, mux_tmp_388, or_1020_nl);
  nor_388_nl <= NOT((result_rem_11cyc_st_3(3)) OR (NOT mux_tmp_389));
  or_1019_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_390 <= MUX_s_1_2_2(nor_388_nl, mux_tmp_389, or_1019_nl);
  nor_389_nl <= NOT((result_rem_11cyc_st_2(3)) OR (NOT mux_tmp_390));
  or_1018_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_391 <= MUX_s_1_2_2(nor_389_nl, mux_tmp_390, or_1018_nl);
  and_697_nl <= not_tmp_645 AND mux_tmp_391;
  mux_tmp_392 <= MUX_s_1_2_2(and_697_nl, mux_tmp_391, or_933_cse);
  and_698_nl <= nand_146_cse AND mux_tmp_392;
  or_1016_nl <= CONV_SL_1_1(result_result_acc_tmp(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_393 <= MUX_s_1_2_2(and_698_nl, mux_tmp_392, or_1016_nl);
  and_dcpl_590 <= and_dcpl_532 AND and_dcpl_352;
  or_tmp_1017 <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR not_tmp_645;
  or_1037_cse <= CONV_SL_1_1(result_result_acc_tmp/=STD_LOGIC_VECTOR'("1010"));
  nor_382_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_1017));
  mux_394_nl <= MUX_s_1_2_2(nor_382_nl, or_tmp_1017, or_1037_cse);
  and_dcpl_592 <= mux_394_nl AND and_dcpl_205;
  or_1042_cse <= CONV_SL_1_1(result_rem_11cyc(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_381_nl <= NOT(and_749_cse OR and_dcpl_205);
  or_1044_nl <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_202);
  mux_tmp_395 <= MUX_s_1_2_2(nor_381_nl, or_1044_nl, or_1042_cse);
  nor_380_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_395));
  mux_396_nl <= MUX_s_1_2_2(nor_380_nl, mux_tmp_395, or_1037_cse);
  and_dcpl_594 <= mux_396_nl AND and_dcpl_179;
  or_1049_cse <= CONV_SL_1_1(result_rem_11cyc_st_2(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_379_nl <= NOT(and_747_cse OR and_dcpl_179);
  or_1051_nl <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_176);
  mux_tmp_397 <= MUX_s_1_2_2(nor_379_nl, or_1051_nl, or_1049_cse);
  and_695_nl <= not_tmp_645 AND mux_tmp_397;
  mux_tmp_398 <= MUX_s_1_2_2(and_695_nl, mux_tmp_397, or_1042_cse);
  nor_378_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_398));
  mux_399_nl <= MUX_s_1_2_2(nor_378_nl, mux_tmp_398, or_1037_cse);
  and_dcpl_596 <= mux_399_nl AND and_dcpl_153;
  or_1058_cse <= CONV_SL_1_1(result_rem_11cyc_st_3(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_377_nl <= NOT(and_744_cse OR and_dcpl_153);
  or_1060_nl <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_150);
  mux_tmp_400 <= MUX_s_1_2_2(nor_377_nl, or_1060_nl, or_1058_cse);
  and_692_nl <= nand_58_cse AND mux_tmp_400;
  mux_tmp_401 <= MUX_s_1_2_2(and_692_nl, mux_tmp_400, or_1049_cse);
  and_693_nl <= not_tmp_645 AND mux_tmp_401;
  mux_tmp_402 <= MUX_s_1_2_2(and_693_nl, mux_tmp_401, or_1042_cse);
  nor_376_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_402));
  mux_403_nl <= MUX_s_1_2_2(nor_376_nl, mux_tmp_402, or_1037_cse);
  and_dcpl_599 <= mux_403_nl AND and_dcpl_127;
  or_1069_cse <= CONV_SL_1_1(result_rem_11cyc_st_4(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_375_nl <= NOT(and_740_cse OR and_dcpl_127);
  or_1071_nl <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1010")) OR
      (NOT and_dcpl_105);
  mux_tmp_404 <= MUX_s_1_2_2(nor_375_nl, or_1071_nl, or_1069_cse);
  and_688_nl <= nand_55_cse AND mux_tmp_404;
  mux_tmp_405 <= MUX_s_1_2_2(and_688_nl, mux_tmp_404, or_1058_cse);
  and_689_nl <= nand_58_cse AND mux_tmp_405;
  mux_tmp_406 <= MUX_s_1_2_2(and_689_nl, mux_tmp_405, or_1049_cse);
  and_690_nl <= not_tmp_645 AND mux_tmp_406;
  mux_tmp_407 <= MUX_s_1_2_2(and_690_nl, mux_tmp_406, or_1042_cse);
  nor_374_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_407));
  mux_408_nl <= MUX_s_1_2_2(nor_374_nl, mux_tmp_407, or_1037_cse);
  and_dcpl_601 <= mux_408_nl AND and_dcpl_102;
  or_1082_cse <= CONV_SL_1_1(result_rem_11cyc_st_5/=STD_LOGIC_VECTOR'("1010"));
  nor_373_nl <= NOT(and_dcpl_105 OR and_dcpl_102);
  or_1084_nl <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_99);
  mux_tmp_409 <= MUX_s_1_2_2(nor_373_nl, or_1084_nl, or_1082_cse);
  and_683_nl <= nand_51_cse AND mux_tmp_409;
  mux_tmp_410 <= MUX_s_1_2_2(and_683_nl, mux_tmp_409, or_1069_cse);
  and_684_nl <= nand_55_cse AND mux_tmp_410;
  mux_tmp_411 <= MUX_s_1_2_2(and_684_nl, mux_tmp_410, or_1058_cse);
  and_685_nl <= nand_58_cse AND mux_tmp_411;
  mux_tmp_412 <= MUX_s_1_2_2(and_685_nl, mux_tmp_411, or_1049_cse);
  and_686_nl <= not_tmp_645 AND mux_tmp_412;
  mux_tmp_413 <= MUX_s_1_2_2(and_686_nl, mux_tmp_412, or_1042_cse);
  nor_372_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_413));
  mux_414_nl <= MUX_s_1_2_2(nor_372_nl, mux_tmp_413, or_1037_cse);
  and_dcpl_603 <= mux_414_nl AND and_dcpl_76;
  or_1097_cse <= CONV_SL_1_1(result_rem_11cyc_st_6(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  nor_370_nl <= NOT(and_731_cse OR and_dcpl_76);
  or_1099_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT and_dcpl_73);
  mux_tmp_415 <= MUX_s_1_2_2(nor_370_nl, or_1099_nl, or_1097_cse);
  nor_371_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_415));
  mux_tmp_416 <= MUX_s_1_2_2(nor_371_nl, mux_tmp_415, or_1082_cse);
  and_679_nl <= nand_51_cse AND mux_tmp_416;
  mux_tmp_417 <= MUX_s_1_2_2(and_679_nl, mux_tmp_416, or_1069_cse);
  and_680_nl <= nand_55_cse AND mux_tmp_417;
  mux_tmp_418 <= MUX_s_1_2_2(and_680_nl, mux_tmp_417, or_1058_cse);
  and_681_nl <= nand_58_cse AND mux_tmp_418;
  mux_tmp_419 <= MUX_s_1_2_2(and_681_nl, mux_tmp_418, or_1049_cse);
  and_682_nl <= not_tmp_645 AND mux_tmp_419;
  mux_tmp_420 <= MUX_s_1_2_2(and_682_nl, mux_tmp_419, or_1042_cse);
  nor_369_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_420));
  mux_421_nl <= MUX_s_1_2_2(nor_369_nl, mux_tmp_420, or_1037_cse);
  and_dcpl_607 <= mux_421_nl AND and_dcpl_50;
  nor_366_nl <= NOT(and_725_cse OR and_dcpl_50);
  or_1116_nl <= CONV_SL_1_1(result_rem_11cyc_st_8/=STD_LOGIC_VECTOR'("1010")) OR
      (NOT and_dcpl_28);
  or_1114_nl <= CONV_SL_1_1(result_rem_11cyc_st_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_422 <= MUX_s_1_2_2(nor_366_nl, or_1116_nl, or_1114_nl);
  and_673_nl <= nand_42_cse AND mux_tmp_422;
  mux_tmp_423 <= MUX_s_1_2_2(and_673_nl, mux_tmp_422, or_1097_cse);
  nor_367_nl <= NOT(and_dcpl_105 OR (NOT mux_tmp_423));
  mux_tmp_424 <= MUX_s_1_2_2(nor_367_nl, mux_tmp_423, or_1082_cse);
  and_674_nl <= nand_51_cse AND mux_tmp_424;
  mux_tmp_425 <= MUX_s_1_2_2(and_674_nl, mux_tmp_424, or_1069_cse);
  and_675_nl <= nand_55_cse AND mux_tmp_425;
  mux_tmp_426 <= MUX_s_1_2_2(and_675_nl, mux_tmp_425, or_1058_cse);
  and_676_nl <= nand_58_cse AND mux_tmp_426;
  mux_tmp_427 <= MUX_s_1_2_2(and_676_nl, mux_tmp_426, or_1049_cse);
  and_677_nl <= not_tmp_645 AND mux_tmp_427;
  mux_tmp_428 <= MUX_s_1_2_2(and_677_nl, mux_tmp_427, or_1042_cse);
  nor_368_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_428));
  mux_429_nl <= MUX_s_1_2_2(nor_368_nl, mux_tmp_428, or_1037_cse);
  and_dcpl_611 <= mux_429_nl AND and_dcpl_4 AND (result_rem_11cyc_st_9(3)) AND (result_rem_11cyc_st_9(1))
      AND (NOT (result_rem_11cyc_st_9(0)));
  or_tmp_1113 <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(result_rem_11cyc_st_9/=STD_LOGIC_VECTOR'("1010"));
  nor_358_nl <= NOT((result_rem_11cyc_st_8(3)) OR (NOT or_tmp_1113));
  or_1133_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(result_rem_11cyc_st_8(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_430 <= MUX_s_1_2_2(nor_358_nl, or_tmp_1113, or_1133_nl);
  nor_359_nl <= NOT((result_rem_11cyc_st_7(3)) OR (NOT mux_tmp_430));
  or_1132_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(result_rem_11cyc_st_7(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_431 <= MUX_s_1_2_2(nor_359_nl, mux_tmp_430, or_1132_nl);
  nor_360_nl <= NOT((result_rem_11cyc_st_6(3)) OR (NOT mux_tmp_431));
  or_1131_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(result_rem_11cyc_st_6(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_432 <= MUX_s_1_2_2(nor_360_nl, mux_tmp_431, or_1131_nl);
  nor_361_nl <= NOT((result_rem_11cyc_st_5(3)) OR (NOT mux_tmp_432));
  or_1130_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(result_rem_11cyc_st_5(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_433 <= MUX_s_1_2_2(nor_361_nl, mux_tmp_432, or_1130_nl);
  nor_362_nl <= NOT((result_rem_11cyc_st_4(3)) OR (NOT mux_tmp_433));
  or_1129_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(result_rem_11cyc_st_4(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_434 <= MUX_s_1_2_2(nor_362_nl, mux_tmp_433, or_1129_nl);
  nor_363_nl <= NOT((result_rem_11cyc_st_3(3)) OR (NOT mux_tmp_434));
  or_1128_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(result_rem_11cyc_st_3(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_435 <= MUX_s_1_2_2(nor_363_nl, mux_tmp_434, or_1128_nl);
  nor_364_nl <= NOT((result_rem_11cyc_st_2(3)) OR (NOT mux_tmp_435));
  or_1127_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(result_rem_11cyc_st_2(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_436 <= MUX_s_1_2_2(nor_364_nl, mux_tmp_435, or_1127_nl);
  and_671_nl <= not_tmp_645 AND mux_tmp_436;
  mux_tmp_437 <= MUX_s_1_2_2(and_671_nl, mux_tmp_436, or_1042_cse);
  nor_365_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_437));
  mux_tmp_438 <= MUX_s_1_2_2(nor_365_nl, mux_tmp_437, or_1037_cse);
  return_rsci_d_mx0c0 <= and_dcpl_235 AND and_dcpl_233;
  return_rsci_d_mx0c1 <= and_dcpl_235 AND and_dcpl_237;
  return_rsci_d_mx0c2 <= and_dcpl_235 AND and_dcpl_240;
  return_rsci_d_mx0c3 <= and_dcpl_235 AND and_dcpl_239 AND (result_rem_11cyc_st_11(0));
  return_rsci_d_mx0c4 <= and_dcpl_235 AND and_dcpl_244 AND (NOT (result_rem_11cyc_st_11(0)));
  return_rsci_d_mx0c5 <= and_dcpl_235 AND and_dcpl_244 AND (result_rem_11cyc_st_11(0));
  return_rsci_d_mx0c6 <= and_dcpl_235 AND and_dcpl_249 AND (NOT (result_rem_11cyc_st_11(0)));
  return_rsci_d_mx0c7 <= and_dcpl_235 AND and_dcpl_249 AND (result_rem_11cyc_st_11(0));
  return_rsci_d_mx0c8 <= and_dcpl_254 AND and_dcpl_233;
  return_rsci_d_mx0c9 <= and_dcpl_254 AND and_dcpl_237;
  return_rsci_d_mx0c10 <= and_dcpl_254 AND and_dcpl_240;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( (ccs_ccore_en AND (return_rsci_d_mx0c0 OR return_rsci_d_mx0c1 OR return_rsci_d_mx0c2
          OR return_rsci_d_mx0c3 OR return_rsci_d_mx0c4 OR return_rsci_d_mx0c5 OR
          return_rsci_d_mx0c6 OR return_rsci_d_mx0c7 OR return_rsci_d_mx0c8 OR return_rsci_d_mx0c9
          OR return_rsci_d_mx0c10)) = '1' ) THEN
        return_rsci_d <= MUX1HOT_v_64_11_2(result_rem_12_cmp_1_z, result_rem_12_cmp_2_z,
            result_rem_12_cmp_3_z, result_rem_12_cmp_4_z, result_rem_12_cmp_5_z,
            result_rem_12_cmp_6_z, result_rem_12_cmp_7_z, result_rem_12_cmp_8_z,
            result_rem_12_cmp_9_z, result_rem_12_cmp_10_z, result_rem_12_cmp_z, STD_LOGIC_VECTOR'(
            return_rsci_d_mx0c0 & return_rsci_d_mx0c1 & return_rsci_d_mx0c2 & return_rsci_d_mx0c3
            & return_rsci_d_mx0c4 & return_rsci_d_mx0c5 & return_rsci_d_mx0c6 & return_rsci_d_mx0c7
            & return_rsci_d_mx0c8 & return_rsci_d_mx0c9 & return_rsci_d_mx0c10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_11 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND main_stage_0_11 AND asn_itm_10) = '1' ) THEN
        result_rem_11cyc_st_11 <= result_rem_11cyc_st_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        asn_itm_11 <= '0';
        asn_itm_10 <= '0';
        asn_itm_9 <= '0';
        asn_itm_8 <= '0';
        asn_itm_7 <= '0';
        asn_itm_6 <= '0';
        asn_itm_5 <= '0';
        asn_itm_4 <= '0';
        asn_itm_3 <= '0';
        asn_itm_2 <= '0';
        asn_itm_1 <= '0';
        main_stage_0_2 <= '0';
        main_stage_0_3 <= '0';
        main_stage_0_4 <= '0';
        main_stage_0_5 <= '0';
        main_stage_0_6 <= '0';
        main_stage_0_7 <= '0';
        main_stage_0_8 <= '0';
        main_stage_0_9 <= '0';
        main_stage_0_10 <= '0';
        main_stage_0_11 <= '0';
        main_stage_0_12 <= '0';
      ELSIF ( ccs_ccore_en = '1' ) THEN
        asn_itm_11 <= asn_itm_10;
        asn_itm_10 <= asn_itm_9;
        asn_itm_9 <= asn_itm_8;
        asn_itm_8 <= asn_itm_7;
        asn_itm_7 <= asn_itm_6;
        asn_itm_6 <= asn_itm_5;
        asn_itm_5 <= asn_itm_4;
        asn_itm_4 <= asn_itm_3;
        asn_itm_3 <= asn_itm_2;
        asn_itm_2 <= asn_itm_1;
        asn_itm_1 <= ccs_ccore_start_rsci_idat;
        main_stage_0_2 <= '1';
        main_stage_0_3 <= main_stage_0_2;
        main_stage_0_4 <= main_stage_0_3;
        main_stage_0_5 <= main_stage_0_4;
        main_stage_0_6 <= main_stage_0_5;
        main_stage_0_7 <= main_stage_0_6;
        main_stage_0_8 <= main_stage_0_7;
        main_stage_0_9 <= main_stage_0_8;
        main_stage_0_10 <= main_stage_0_9;
        main_stage_0_11 <= main_stage_0_10;
        main_stage_0_12 <= main_stage_0_11;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_1_cse = '1' ) THEN
        result_rem_12_cmp_1_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_1_2,
            m_buf_sva_mut_1_3, m_buf_sva_mut_1_4, m_buf_sva_mut_1_5, m_buf_sva_mut_1_6,
            m_buf_sva_mut_1_7, m_buf_sva_mut_1_8, m_buf_sva_mut_1_9, m_buf_sva_mut_1_10,
            STD_LOGIC_VECTOR'( and_dcpl_263 & and_dcpl_269 & and_dcpl_275 & and_dcpl_281
            & and_dcpl_287 & and_dcpl_293 & and_dcpl_299 & and_dcpl_305 & and_dcpl_311
            & mux_tmp_37));
        result_rem_12_cmp_1_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_1_2,
            base_buf_sva_mut_1_3, base_buf_sva_mut_1_4, base_buf_sva_mut_1_5, base_buf_sva_mut_1_6,
            base_buf_sva_mut_1_7, base_buf_sva_mut_1_8, base_buf_sva_mut_1_9, base_buf_sva_mut_1_10,
            STD_LOGIC_VECTOR'( and_dcpl_263 & and_dcpl_269 & and_dcpl_275 & and_dcpl_281
            & and_dcpl_287 & and_dcpl_293 & and_dcpl_299 & and_dcpl_305 & and_dcpl_311
            & mux_tmp_37));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_3_cse = '1' ) THEN
        result_rem_12_cmp_2_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_2_2,
            m_buf_sva_mut_2_3, m_buf_sva_mut_2_4, m_buf_sva_mut_2_5, m_buf_sva_mut_2_6,
            m_buf_sva_mut_2_7, m_buf_sva_mut_2_8, m_buf_sva_mut_2_9, m_buf_sva_mut_2_10,
            STD_LOGIC_VECTOR'( and_dcpl_319 & and_dcpl_322 & and_dcpl_325 & and_dcpl_329
            & and_dcpl_333 & and_dcpl_337 & and_dcpl_341 & and_dcpl_344 & and_dcpl_347
            & mux_tmp_75));
        result_rem_12_cmp_2_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_2_2,
            base_buf_sva_mut_2_3, base_buf_sva_mut_2_4, base_buf_sva_mut_2_5, base_buf_sva_mut_2_6,
            base_buf_sva_mut_2_7, base_buf_sva_mut_2_8, base_buf_sva_mut_2_9, base_buf_sva_mut_2_10,
            STD_LOGIC_VECTOR'( and_dcpl_319 & and_dcpl_322 & and_dcpl_325 & and_dcpl_329
            & and_dcpl_333 & and_dcpl_337 & and_dcpl_341 & and_dcpl_344 & and_dcpl_347
            & mux_tmp_75));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_5_cse = '1' ) THEN
        result_rem_12_cmp_3_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_3_2,
            m_buf_sva_mut_3_3, m_buf_sva_mut_3_4, m_buf_sva_mut_3_5, m_buf_sva_mut_3_6,
            m_buf_sva_mut_3_7, m_buf_sva_mut_3_8, m_buf_sva_mut_3_9, m_buf_sva_mut_3_10,
            STD_LOGIC_VECTOR'( and_dcpl_353 & and_dcpl_357 & and_dcpl_361 & and_dcpl_364
            & and_dcpl_367 & and_dcpl_370 & and_dcpl_373 & and_dcpl_377 & and_dcpl_381
            & mux_tmp_113));
        result_rem_12_cmp_3_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_3_2,
            base_buf_sva_mut_3_3, base_buf_sva_mut_3_4, base_buf_sva_mut_3_5, base_buf_sva_mut_3_6,
            base_buf_sva_mut_3_7, base_buf_sva_mut_3_8, base_buf_sva_mut_3_9, base_buf_sva_mut_3_10,
            STD_LOGIC_VECTOR'( and_dcpl_353 & and_dcpl_357 & and_dcpl_361 & and_dcpl_364
            & and_dcpl_367 & and_dcpl_370 & and_dcpl_373 & and_dcpl_377 & and_dcpl_381
            & mux_tmp_113));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_7_cse = '1' ) THEN
        result_rem_12_cmp_4_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_4_2,
            m_buf_sva_mut_4_3, m_buf_sva_mut_4_4, m_buf_sva_mut_4_5, m_buf_sva_mut_4_6,
            m_buf_sva_mut_4_7, m_buf_sva_mut_4_8, m_buf_sva_mut_4_9, m_buf_sva_mut_4_10,
            STD_LOGIC_VECTOR'( and_dcpl_387 & and_dcpl_390 & and_dcpl_393 & and_dcpl_396
            & and_dcpl_399 & and_dcpl_402 & and_dcpl_405 & and_dcpl_408 & and_dcpl_411
            & mux_tmp_151));
        result_rem_12_cmp_4_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_4_2,
            base_buf_sva_mut_4_3, base_buf_sva_mut_4_4, base_buf_sva_mut_4_5, base_buf_sva_mut_4_6,
            base_buf_sva_mut_4_7, base_buf_sva_mut_4_8, base_buf_sva_mut_4_9, base_buf_sva_mut_4_10,
            STD_LOGIC_VECTOR'( and_dcpl_387 & and_dcpl_390 & and_dcpl_393 & and_dcpl_396
            & and_dcpl_399 & and_dcpl_402 & and_dcpl_405 & and_dcpl_408 & and_dcpl_411
            & mux_tmp_151));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_9_cse = '1' ) THEN
        result_rem_12_cmp_5_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_5_2,
            m_buf_sva_mut_5_3, m_buf_sva_mut_5_4, m_buf_sva_mut_5_5, m_buf_sva_mut_5_6,
            m_buf_sva_mut_5_7, m_buf_sva_mut_5_8, m_buf_sva_mut_5_9, m_buf_sva_mut_5_10,
            STD_LOGIC_VECTOR'( and_dcpl_418 & and_dcpl_422 & and_dcpl_426 & and_dcpl_430
            & and_dcpl_433 & and_dcpl_437 & and_dcpl_441 & and_dcpl_444 & and_dcpl_447
            & mux_tmp_189));
        result_rem_12_cmp_5_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_5_2,
            base_buf_sva_mut_5_3, base_buf_sva_mut_5_4, base_buf_sva_mut_5_5, base_buf_sva_mut_5_6,
            base_buf_sva_mut_5_7, base_buf_sva_mut_5_8, base_buf_sva_mut_5_9, base_buf_sva_mut_5_10,
            STD_LOGIC_VECTOR'( and_dcpl_418 & and_dcpl_422 & and_dcpl_426 & and_dcpl_430
            & and_dcpl_433 & and_dcpl_437 & and_dcpl_441 & and_dcpl_444 & and_dcpl_447
            & mux_tmp_189));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_11_cse = '1' ) THEN
        result_rem_12_cmp_6_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_6_2,
            m_buf_sva_mut_6_3, m_buf_sva_mut_6_4, m_buf_sva_mut_6_5, m_buf_sva_mut_6_6,
            m_buf_sva_mut_6_7, m_buf_sva_mut_6_8, m_buf_sva_mut_6_9, m_buf_sva_mut_6_10,
            STD_LOGIC_VECTOR'( and_dcpl_452 & and_dcpl_455 & and_dcpl_458 & and_dcpl_462
            & and_dcpl_464 & and_dcpl_468 & and_dcpl_472 & and_dcpl_474 & and_dcpl_476
            & mux_tmp_227));
        result_rem_12_cmp_6_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_6_2,
            base_buf_sva_mut_6_3, base_buf_sva_mut_6_4, base_buf_sva_mut_6_5, base_buf_sva_mut_6_6,
            base_buf_sva_mut_6_7, base_buf_sva_mut_6_8, base_buf_sva_mut_6_9, base_buf_sva_mut_6_10,
            STD_LOGIC_VECTOR'( and_dcpl_452 & and_dcpl_455 & and_dcpl_458 & and_dcpl_462
            & and_dcpl_464 & and_dcpl_468 & and_dcpl_472 & and_dcpl_474 & and_dcpl_476
            & mux_tmp_227));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_13_cse = '1' ) THEN
        result_rem_12_cmp_7_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_7_2,
            m_buf_sva_mut_7_3, m_buf_sva_mut_7_4, m_buf_sva_mut_7_5, m_buf_sva_mut_7_6,
            m_buf_sva_mut_7_7, m_buf_sva_mut_7_8, m_buf_sva_mut_7_9, m_buf_sva_mut_7_10,
            STD_LOGIC_VECTOR'( and_dcpl_480 & and_dcpl_484 & and_dcpl_488 & and_dcpl_491
            & and_dcpl_493 & and_dcpl_496 & and_dcpl_499 & and_dcpl_501 & and_dcpl_503
            & mux_tmp_265));
        result_rem_12_cmp_7_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_7_2,
            base_buf_sva_mut_7_3, base_buf_sva_mut_7_4, base_buf_sva_mut_7_5, base_buf_sva_mut_7_6,
            base_buf_sva_mut_7_7, base_buf_sva_mut_7_8, base_buf_sva_mut_7_9, base_buf_sva_mut_7_10,
            STD_LOGIC_VECTOR'( and_dcpl_480 & and_dcpl_484 & and_dcpl_488 & and_dcpl_491
            & and_dcpl_493 & and_dcpl_496 & and_dcpl_499 & and_dcpl_501 & and_dcpl_503
            & mux_tmp_265));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_15_cse = '1' ) THEN
        result_rem_12_cmp_8_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_8_2,
            m_buf_sva_mut_8_3, m_buf_sva_mut_8_4, m_buf_sva_mut_8_5, m_buf_sva_mut_8_6,
            m_buf_sva_mut_8_7, m_buf_sva_mut_8_8, m_buf_sva_mut_8_9, m_buf_sva_mut_8_10,
            STD_LOGIC_VECTOR'( and_dcpl_507 & and_dcpl_510 & and_dcpl_513 & and_dcpl_516
            & and_dcpl_518 & and_dcpl_521 & and_dcpl_524 & and_dcpl_526 & and_dcpl_528
            & mux_tmp_303));
        result_rem_12_cmp_8_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_8_2,
            base_buf_sva_mut_8_3, base_buf_sva_mut_8_4, base_buf_sva_mut_8_5, base_buf_sva_mut_8_6,
            base_buf_sva_mut_8_7, base_buf_sva_mut_8_8, base_buf_sva_mut_8_9, base_buf_sva_mut_8_10,
            STD_LOGIC_VECTOR'( and_dcpl_507 & and_dcpl_510 & and_dcpl_513 & and_dcpl_516
            & and_dcpl_518 & and_dcpl_521 & and_dcpl_524 & and_dcpl_526 & and_dcpl_528
            & mux_tmp_303));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_17_cse = '1' ) THEN
        result_rem_12_cmp_9_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_9_2,
            m_buf_sva_mut_9_3, m_buf_sva_mut_9_4, m_buf_sva_mut_9_5, m_buf_sva_mut_9_6,
            m_buf_sva_mut_9_7, m_buf_sva_mut_9_8, m_buf_sva_mut_9_9, m_buf_sva_mut_9_10,
            STD_LOGIC_VECTOR'( and_dcpl_533 & and_dcpl_536 & and_dcpl_539 & and_dcpl_542
            & and_dcpl_546 & and_dcpl_549 & and_dcpl_552 & and_dcpl_556 & and_dcpl_560
            & mux_tmp_348));
        result_rem_12_cmp_9_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_9_2,
            base_buf_sva_mut_9_3, base_buf_sva_mut_9_4, base_buf_sva_mut_9_5, base_buf_sva_mut_9_6,
            base_buf_sva_mut_9_7, base_buf_sva_mut_9_8, base_buf_sva_mut_9_9, base_buf_sva_mut_9_10,
            STD_LOGIC_VECTOR'( and_dcpl_533 & and_dcpl_536 & and_dcpl_539 & and_dcpl_542
            & and_dcpl_546 & and_dcpl_549 & and_dcpl_552 & and_dcpl_556 & and_dcpl_560
            & mux_tmp_348));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_19_cse = '1' ) THEN
        result_rem_12_cmp_10_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_10_2,
            m_buf_sva_mut_10_3, m_buf_sva_mut_10_4, m_buf_sva_mut_10_5, m_buf_sva_mut_10_6,
            m_buf_sva_mut_10_7, m_buf_sva_mut_10_8, m_buf_sva_mut_10_9, m_buf_sva_mut_10_10,
            STD_LOGIC_VECTOR'( and_dcpl_566 & and_dcpl_568 & and_dcpl_570 & and_dcpl_572
            & and_dcpl_576 & and_dcpl_578 & and_dcpl_580 & and_dcpl_583 & and_dcpl_586
            & mux_tmp_393));
        result_rem_12_cmp_10_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_10_2,
            base_buf_sva_mut_10_3, base_buf_sva_mut_10_4, base_buf_sva_mut_10_5,
            base_buf_sva_mut_10_6, base_buf_sva_mut_10_7, base_buf_sva_mut_10_8,
            base_buf_sva_mut_10_9, base_buf_sva_mut_10_10, STD_LOGIC_VECTOR'( and_dcpl_566
            & and_dcpl_568 & and_dcpl_570 & and_dcpl_572 & and_dcpl_576 & and_dcpl_578
            & and_dcpl_580 & and_dcpl_583 & and_dcpl_586 & mux_tmp_393));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( result_and_21_cse = '1' ) THEN
        result_rem_12_cmp_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_2, m_buf_sva_mut_3,
            m_buf_sva_mut_4, m_buf_sva_mut_5, m_buf_sva_mut_6, m_buf_sva_mut_7, m_buf_sva_mut_8,
            m_buf_sva_mut_9, m_buf_sva_mut_10, STD_LOGIC_VECTOR'( and_dcpl_590 &
            and_dcpl_592 & and_dcpl_594 & and_dcpl_596 & and_dcpl_599 & and_dcpl_601
            & and_dcpl_603 & and_dcpl_607 & and_dcpl_611 & mux_tmp_438));
        result_rem_12_cmp_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_2,
            base_buf_sva_mut_3, base_buf_sva_mut_4, base_buf_sva_mut_5, base_buf_sva_mut_6,
            base_buf_sva_mut_7, base_buf_sva_mut_8, base_buf_sva_mut_9, base_buf_sva_mut_10,
            STD_LOGIC_VECTOR'( and_dcpl_590 & and_dcpl_592 & and_dcpl_594 & and_dcpl_596
            & and_dcpl_599 & and_dcpl_601 & and_dcpl_603 & and_dcpl_607 & and_dcpl_611
            & mux_tmp_438));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_cse = '1' ) THEN
        m_buf_sva_mut_1_10 <= m_buf_sva_mut_1_9;
        base_buf_sva_mut_1_10 <= base_buf_sva_mut_1_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_1_cse = '1' ) THEN
        m_buf_sva_mut_2_10 <= m_buf_sva_mut_2_9;
        base_buf_sva_mut_2_10 <= base_buf_sva_mut_2_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_2_cse = '1' ) THEN
        m_buf_sva_mut_3_10 <= m_buf_sva_mut_3_9;
        base_buf_sva_mut_3_10 <= base_buf_sva_mut_3_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_3_cse = '1' ) THEN
        m_buf_sva_mut_4_10 <= m_buf_sva_mut_4_9;
        base_buf_sva_mut_4_10 <= base_buf_sva_mut_4_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_4_cse = '1' ) THEN
        m_buf_sva_mut_5_10 <= m_buf_sva_mut_5_9;
        base_buf_sva_mut_5_10 <= base_buf_sva_mut_5_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_5_cse = '1' ) THEN
        m_buf_sva_mut_6_10 <= m_buf_sva_mut_6_9;
        base_buf_sva_mut_6_10 <= base_buf_sva_mut_6_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_6_cse = '1' ) THEN
        m_buf_sva_mut_7_10 <= m_buf_sva_mut_7_9;
        base_buf_sva_mut_7_10 <= base_buf_sva_mut_7_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_7_cse = '1' ) THEN
        m_buf_sva_mut_8_10 <= m_buf_sva_mut_8_9;
        base_buf_sva_mut_8_10 <= base_buf_sva_mut_8_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_8_cse = '1' ) THEN
        m_buf_sva_mut_9_10 <= m_buf_sva_mut_9_9;
        base_buf_sva_mut_9_10 <= base_buf_sva_mut_9_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_9_cse = '1' ) THEN
        m_buf_sva_mut_10_10 <= m_buf_sva_mut_10_9;
        base_buf_sva_mut_10_10 <= base_buf_sva_mut_10_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_10_cse = '1' ) THEN
        m_buf_sva_mut_10 <= m_buf_sva_mut_9;
        base_buf_sva_mut_10 <= base_buf_sva_mut_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_10 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_3) = '1' ) THEN
        result_rem_11cyc_st_10 <= result_rem_11cyc_st_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_11_cse = '1' ) THEN
        m_buf_sva_mut_1_9 <= m_buf_sva_mut_1_8;
        base_buf_sva_mut_1_9 <= base_buf_sva_mut_1_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_12_cse = '1' ) THEN
        m_buf_sva_mut_2_9 <= m_buf_sva_mut_2_8;
        base_buf_sva_mut_2_9 <= base_buf_sva_mut_2_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_13_cse = '1' ) THEN
        m_buf_sva_mut_3_9 <= m_buf_sva_mut_3_8;
        base_buf_sva_mut_3_9 <= base_buf_sva_mut_3_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_14_cse = '1' ) THEN
        m_buf_sva_mut_4_9 <= m_buf_sva_mut_4_8;
        base_buf_sva_mut_4_9 <= base_buf_sva_mut_4_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_15_cse = '1' ) THEN
        m_buf_sva_mut_5_9 <= m_buf_sva_mut_5_8;
        base_buf_sva_mut_5_9 <= base_buf_sva_mut_5_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_16_cse = '1' ) THEN
        m_buf_sva_mut_6_9 <= m_buf_sva_mut_6_8;
        base_buf_sva_mut_6_9 <= base_buf_sva_mut_6_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_17_cse = '1' ) THEN
        m_buf_sva_mut_7_9 <= m_buf_sva_mut_7_8;
        base_buf_sva_mut_7_9 <= base_buf_sva_mut_7_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_18_cse = '1' ) THEN
        m_buf_sva_mut_8_9 <= m_buf_sva_mut_8_8;
        base_buf_sva_mut_8_9 <= base_buf_sva_mut_8_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_19_cse = '1' ) THEN
        m_buf_sva_mut_9_9 <= m_buf_sva_mut_9_8;
        base_buf_sva_mut_9_9 <= base_buf_sva_mut_9_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_20_cse = '1' ) THEN
        m_buf_sva_mut_10_9 <= m_buf_sva_mut_10_8;
        base_buf_sva_mut_10_9 <= base_buf_sva_mut_10_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_21_cse = '1' ) THEN
        m_buf_sva_mut_9 <= m_buf_sva_mut_8;
        base_buf_sva_mut_9 <= base_buf_sva_mut_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_9 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_28) = '1' ) THEN
        result_rem_11cyc_st_9 <= result_rem_11cyc_st_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_22_cse = '1' ) THEN
        m_buf_sva_mut_1_8 <= m_buf_sva_mut_1_7;
        base_buf_sva_mut_1_8 <= base_buf_sva_mut_1_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_23_cse = '1' ) THEN
        m_buf_sva_mut_2_8 <= m_buf_sva_mut_2_7;
        base_buf_sva_mut_2_8 <= base_buf_sva_mut_2_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_24_cse = '1' ) THEN
        m_buf_sva_mut_3_8 <= m_buf_sva_mut_3_7;
        base_buf_sva_mut_3_8 <= base_buf_sva_mut_3_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_25_cse = '1' ) THEN
        m_buf_sva_mut_4_8 <= m_buf_sva_mut_4_7;
        base_buf_sva_mut_4_8 <= base_buf_sva_mut_4_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_26_cse = '1' ) THEN
        m_buf_sva_mut_5_8 <= m_buf_sva_mut_5_7;
        base_buf_sva_mut_5_8 <= base_buf_sva_mut_5_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_27_cse = '1' ) THEN
        m_buf_sva_mut_6_8 <= m_buf_sva_mut_6_7;
        base_buf_sva_mut_6_8 <= base_buf_sva_mut_6_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_28_cse = '1' ) THEN
        m_buf_sva_mut_7_8 <= m_buf_sva_mut_7_7;
        base_buf_sva_mut_7_8 <= base_buf_sva_mut_7_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_29_cse = '1' ) THEN
        m_buf_sva_mut_8_8 <= m_buf_sva_mut_8_7;
        base_buf_sva_mut_8_8 <= base_buf_sva_mut_8_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_30_cse = '1' ) THEN
        m_buf_sva_mut_9_8 <= m_buf_sva_mut_9_7;
        base_buf_sva_mut_9_8 <= base_buf_sva_mut_9_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_31_cse = '1' ) THEN
        m_buf_sva_mut_10_8 <= m_buf_sva_mut_10_7;
        base_buf_sva_mut_10_8 <= base_buf_sva_mut_10_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_32_cse = '1' ) THEN
        m_buf_sva_mut_8 <= m_buf_sva_mut_7;
        base_buf_sva_mut_8 <= base_buf_sva_mut_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_8 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_53) = '1' ) THEN
        result_rem_11cyc_st_8 <= result_rem_11cyc_st_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_33_cse = '1' ) THEN
        m_buf_sva_mut_1_7 <= m_buf_sva_mut_1_6;
        base_buf_sva_mut_1_7 <= base_buf_sva_mut_1_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_34_cse = '1' ) THEN
        m_buf_sva_mut_2_7 <= m_buf_sva_mut_2_6;
        base_buf_sva_mut_2_7 <= base_buf_sva_mut_2_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_35_cse = '1' ) THEN
        m_buf_sva_mut_3_7 <= m_buf_sva_mut_3_6;
        base_buf_sva_mut_3_7 <= base_buf_sva_mut_3_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_36_cse = '1' ) THEN
        m_buf_sva_mut_4_7 <= m_buf_sva_mut_4_6;
        base_buf_sva_mut_4_7 <= base_buf_sva_mut_4_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_37_cse = '1' ) THEN
        m_buf_sva_mut_5_7 <= m_buf_sva_mut_5_6;
        base_buf_sva_mut_5_7 <= base_buf_sva_mut_5_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_38_cse = '1' ) THEN
        m_buf_sva_mut_6_7 <= m_buf_sva_mut_6_6;
        base_buf_sva_mut_6_7 <= base_buf_sva_mut_6_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_39_cse = '1' ) THEN
        m_buf_sva_mut_7_7 <= m_buf_sva_mut_7_6;
        base_buf_sva_mut_7_7 <= base_buf_sva_mut_7_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_40_cse = '1' ) THEN
        m_buf_sva_mut_8_7 <= m_buf_sva_mut_8_6;
        base_buf_sva_mut_8_7 <= base_buf_sva_mut_8_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_41_cse = '1' ) THEN
        m_buf_sva_mut_9_7 <= m_buf_sva_mut_9_6;
        base_buf_sva_mut_9_7 <= base_buf_sva_mut_9_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_42_cse = '1' ) THEN
        m_buf_sva_mut_10_7 <= m_buf_sva_mut_10_6;
        base_buf_sva_mut_10_7 <= base_buf_sva_mut_10_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_43_cse = '1' ) THEN
        m_buf_sva_mut_7 <= m_buf_sva_mut_6;
        base_buf_sva_mut_7 <= base_buf_sva_mut_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_7 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_79) = '1' ) THEN
        result_rem_11cyc_st_7 <= result_rem_11cyc_st_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_44_cse = '1' ) THEN
        m_buf_sva_mut_1_6 <= m_buf_sva_mut_1_5;
        base_buf_sva_mut_1_6 <= base_buf_sva_mut_1_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_45_cse = '1' ) THEN
        m_buf_sva_mut_2_6 <= m_buf_sva_mut_2_5;
        base_buf_sva_mut_2_6 <= base_buf_sva_mut_2_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_46_cse = '1' ) THEN
        m_buf_sva_mut_3_6 <= m_buf_sva_mut_3_5;
        base_buf_sva_mut_3_6 <= base_buf_sva_mut_3_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_47_cse = '1' ) THEN
        m_buf_sva_mut_4_6 <= m_buf_sva_mut_4_5;
        base_buf_sva_mut_4_6 <= base_buf_sva_mut_4_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_48_cse = '1' ) THEN
        m_buf_sva_mut_5_6 <= m_buf_sva_mut_5_5;
        base_buf_sva_mut_5_6 <= base_buf_sva_mut_5_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_49_cse = '1' ) THEN
        m_buf_sva_mut_6_6 <= m_buf_sva_mut_6_5;
        base_buf_sva_mut_6_6 <= base_buf_sva_mut_6_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_50_cse = '1' ) THEN
        m_buf_sva_mut_7_6 <= m_buf_sva_mut_7_5;
        base_buf_sva_mut_7_6 <= base_buf_sva_mut_7_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_51_cse = '1' ) THEN
        m_buf_sva_mut_8_6 <= m_buf_sva_mut_8_5;
        base_buf_sva_mut_8_6 <= base_buf_sva_mut_8_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_52_cse = '1' ) THEN
        m_buf_sva_mut_9_6 <= m_buf_sva_mut_9_5;
        base_buf_sva_mut_9_6 <= base_buf_sva_mut_9_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_53_cse = '1' ) THEN
        m_buf_sva_mut_10_6 <= m_buf_sva_mut_10_5;
        base_buf_sva_mut_10_6 <= base_buf_sva_mut_10_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_54_cse = '1' ) THEN
        m_buf_sva_mut_6 <= m_buf_sva_mut_5;
        base_buf_sva_mut_6 <= base_buf_sva_mut_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_6 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_105) = '1' ) THEN
        result_rem_11cyc_st_6 <= result_rem_11cyc_st_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_55_cse = '1' ) THEN
        m_buf_sva_mut_1_5 <= m_buf_sva_mut_1_4;
        base_buf_sva_mut_1_5 <= base_buf_sva_mut_1_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_56_cse = '1' ) THEN
        m_buf_sva_mut_2_5 <= m_buf_sva_mut_2_4;
        base_buf_sva_mut_2_5 <= base_buf_sva_mut_2_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_57_cse = '1' ) THEN
        m_buf_sva_mut_3_5 <= m_buf_sva_mut_3_4;
        base_buf_sva_mut_3_5 <= base_buf_sva_mut_3_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_58_cse = '1' ) THEN
        m_buf_sva_mut_4_5 <= m_buf_sva_mut_4_4;
        base_buf_sva_mut_4_5 <= base_buf_sva_mut_4_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_59_cse = '1' ) THEN
        m_buf_sva_mut_5_5 <= m_buf_sva_mut_5_4;
        base_buf_sva_mut_5_5 <= base_buf_sva_mut_5_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_60_cse = '1' ) THEN
        m_buf_sva_mut_6_5 <= m_buf_sva_mut_6_4;
        base_buf_sva_mut_6_5 <= base_buf_sva_mut_6_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_61_cse = '1' ) THEN
        m_buf_sva_mut_7_5 <= m_buf_sva_mut_7_4;
        base_buf_sva_mut_7_5 <= base_buf_sva_mut_7_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_62_cse = '1' ) THEN
        m_buf_sva_mut_8_5 <= m_buf_sva_mut_8_4;
        base_buf_sva_mut_8_5 <= base_buf_sva_mut_8_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_63_cse = '1' ) THEN
        m_buf_sva_mut_9_5 <= m_buf_sva_mut_9_4;
        base_buf_sva_mut_9_5 <= base_buf_sva_mut_9_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_64_cse = '1' ) THEN
        m_buf_sva_mut_10_5 <= m_buf_sva_mut_10_4;
        base_buf_sva_mut_10_5 <= base_buf_sva_mut_10_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_65_cse = '1' ) THEN
        m_buf_sva_mut_5 <= m_buf_sva_mut_4;
        base_buf_sva_mut_5 <= base_buf_sva_mut_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_5 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_130) = '1' ) THEN
        result_rem_11cyc_st_5 <= result_rem_11cyc_st_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_66_cse = '1' ) THEN
        m_buf_sva_mut_1_4 <= m_buf_sva_mut_1_3;
        base_buf_sva_mut_1_4 <= base_buf_sva_mut_1_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_67_cse = '1' ) THEN
        m_buf_sva_mut_2_4 <= m_buf_sva_mut_2_3;
        base_buf_sva_mut_2_4 <= base_buf_sva_mut_2_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_68_cse = '1' ) THEN
        m_buf_sva_mut_3_4 <= m_buf_sva_mut_3_3;
        base_buf_sva_mut_3_4 <= base_buf_sva_mut_3_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_69_cse = '1' ) THEN
        m_buf_sva_mut_4_4 <= m_buf_sva_mut_4_3;
        base_buf_sva_mut_4_4 <= base_buf_sva_mut_4_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_70_cse = '1' ) THEN
        m_buf_sva_mut_5_4 <= m_buf_sva_mut_5_3;
        base_buf_sva_mut_5_4 <= base_buf_sva_mut_5_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_71_cse = '1' ) THEN
        m_buf_sva_mut_6_4 <= m_buf_sva_mut_6_3;
        base_buf_sva_mut_6_4 <= base_buf_sva_mut_6_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_72_cse = '1' ) THEN
        m_buf_sva_mut_7_4 <= m_buf_sva_mut_7_3;
        base_buf_sva_mut_7_4 <= base_buf_sva_mut_7_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_73_cse = '1' ) THEN
        m_buf_sva_mut_8_4 <= m_buf_sva_mut_8_3;
        base_buf_sva_mut_8_4 <= base_buf_sva_mut_8_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_74_cse = '1' ) THEN
        m_buf_sva_mut_9_4 <= m_buf_sva_mut_9_3;
        base_buf_sva_mut_9_4 <= base_buf_sva_mut_9_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_75_cse = '1' ) THEN
        m_buf_sva_mut_10_4 <= m_buf_sva_mut_10_3;
        base_buf_sva_mut_10_4 <= base_buf_sva_mut_10_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_76_cse = '1' ) THEN
        m_buf_sva_mut_4 <= m_buf_sva_mut_3;
        base_buf_sva_mut_4 <= base_buf_sva_mut_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_4 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_156) = '1' ) THEN
        result_rem_11cyc_st_4 <= result_rem_11cyc_st_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_77_cse = '1' ) THEN
        m_buf_sva_mut_1_3 <= m_buf_sva_mut_1_2;
        base_buf_sva_mut_1_3 <= base_buf_sva_mut_1_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_78_cse = '1' ) THEN
        m_buf_sva_mut_2_3 <= m_buf_sva_mut_2_2;
        base_buf_sva_mut_2_3 <= base_buf_sva_mut_2_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_79_cse = '1' ) THEN
        m_buf_sva_mut_3_3 <= m_buf_sva_mut_3_2;
        base_buf_sva_mut_3_3 <= base_buf_sva_mut_3_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_80_cse = '1' ) THEN
        m_buf_sva_mut_4_3 <= m_buf_sva_mut_4_2;
        base_buf_sva_mut_4_3 <= base_buf_sva_mut_4_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_81_cse = '1' ) THEN
        m_buf_sva_mut_5_3 <= m_buf_sva_mut_5_2;
        base_buf_sva_mut_5_3 <= base_buf_sva_mut_5_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_82_cse = '1' ) THEN
        m_buf_sva_mut_6_3 <= m_buf_sva_mut_6_2;
        base_buf_sva_mut_6_3 <= base_buf_sva_mut_6_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_83_cse = '1' ) THEN
        m_buf_sva_mut_7_3 <= m_buf_sva_mut_7_2;
        base_buf_sva_mut_7_3 <= base_buf_sva_mut_7_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_84_cse = '1' ) THEN
        m_buf_sva_mut_8_3 <= m_buf_sva_mut_8_2;
        base_buf_sva_mut_8_3 <= base_buf_sva_mut_8_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_85_cse = '1' ) THEN
        m_buf_sva_mut_9_3 <= m_buf_sva_mut_9_2;
        base_buf_sva_mut_9_3 <= base_buf_sva_mut_9_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_86_cse = '1' ) THEN
        m_buf_sva_mut_10_3 <= m_buf_sva_mut_10_2;
        base_buf_sva_mut_10_3 <= base_buf_sva_mut_10_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_87_cse = '1' ) THEN
        m_buf_sva_mut_3 <= m_buf_sva_mut_2;
        base_buf_sva_mut_3 <= base_buf_sva_mut_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_3 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_182) = '1' ) THEN
        result_rem_11cyc_st_3 <= result_rem_11cyc_st_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_88_cse = '1' ) THEN
        m_buf_sva_mut_1_2 <= result_rem_12_cmp_1_b;
        base_buf_sva_mut_1_2 <= result_rem_12_cmp_1_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_89_cse = '1' ) THEN
        m_buf_sva_mut_2_2 <= result_rem_12_cmp_2_b;
        base_buf_sva_mut_2_2 <= result_rem_12_cmp_2_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_90_cse = '1' ) THEN
        m_buf_sva_mut_3_2 <= result_rem_12_cmp_3_b;
        base_buf_sva_mut_3_2 <= result_rem_12_cmp_3_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_91_cse = '1' ) THEN
        m_buf_sva_mut_4_2 <= result_rem_12_cmp_4_b;
        base_buf_sva_mut_4_2 <= result_rem_12_cmp_4_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_92_cse = '1' ) THEN
        m_buf_sva_mut_5_2 <= result_rem_12_cmp_5_b;
        base_buf_sva_mut_5_2 <= result_rem_12_cmp_5_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_93_cse = '1' ) THEN
        m_buf_sva_mut_6_2 <= result_rem_12_cmp_6_b;
        base_buf_sva_mut_6_2 <= result_rem_12_cmp_6_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_94_cse = '1' ) THEN
        m_buf_sva_mut_7_2 <= result_rem_12_cmp_7_b;
        base_buf_sva_mut_7_2 <= result_rem_12_cmp_7_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_95_cse = '1' ) THEN
        m_buf_sva_mut_8_2 <= result_rem_12_cmp_8_b;
        base_buf_sva_mut_8_2 <= result_rem_12_cmp_8_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_96_cse = '1' ) THEN
        m_buf_sva_mut_9_2 <= result_rem_12_cmp_9_b;
        base_buf_sva_mut_9_2 <= result_rem_12_cmp_9_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_97_cse = '1' ) THEN
        m_buf_sva_mut_10_2 <= result_rem_12_cmp_10_b;
        base_buf_sva_mut_10_2 <= result_rem_12_cmp_10_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( m_and_98_cse = '1' ) THEN
        m_buf_sva_mut_2 <= result_rem_12_cmp_b;
        base_buf_sva_mut_2 <= result_rem_12_cmp_a;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc_st_2 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND and_dcpl_208) = '1' ) THEN
        result_rem_11cyc_st_2 <= result_rem_11cyc;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_rem_11cyc <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (ccs_ccore_en AND ccs_ccore_start_rsci_idat) = '1' ) THEN
        result_rem_11cyc <= result_result_acc_tmp;
      END IF;
    END IF;
  END PROCESS;
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    modulo_dev
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_dev IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_dev;

ARCHITECTURE v1 OF modulo_dev IS
  -- Default Constants

  COMPONENT modulo_dev_core
    PORT(
      base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_dev_core_inst_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_core_inst_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_core_inst_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  modulo_dev_core_inst : modulo_dev_core
    PORT MAP(
      base_rsc_dat => modulo_dev_core_inst_base_rsc_dat,
      m_rsc_dat => modulo_dev_core_inst_m_rsc_dat,
      return_rsc_z => modulo_dev_core_inst_return_rsc_z,
      ccs_ccore_start_rsc_dat => ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_srst => ccs_ccore_srst,
      ccs_ccore_en => ccs_ccore_en
    );
  modulo_dev_core_inst_base_rsc_dat <= base_rsc_dat;
  modulo_dev_core_inst_m_rsc_dat <= m_rsc_dat;
  return_rsc_z <= modulo_dev_core_inst_return_rsc_z;

END v1;




--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Fri Aug 27 10:18:00 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen;

ARCHITECTURE v14 OF inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    COMP_LOOP_C_28_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_56_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_84_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_112_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_140_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_168_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_196_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_224_tr0 : IN STD_LOGIC;
    VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_1_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIF_core_core_fsm;

ARCHITECTURE v14 OF inPlaceNTT_DIF_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIF_core_core_fsm_1
  TYPE inPlaceNTT_DIF_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, COMP_LOOP_C_0,
      COMP_LOOP_C_1, COMP_LOOP_C_2, COMP_LOOP_C_3, COMP_LOOP_C_4, COMP_LOOP_C_5,
      COMP_LOOP_C_6, COMP_LOOP_C_7, COMP_LOOP_C_8, COMP_LOOP_C_9, COMP_LOOP_C_10,
      COMP_LOOP_C_11, COMP_LOOP_C_12, COMP_LOOP_C_13, COMP_LOOP_C_14, COMP_LOOP_C_15,
      COMP_LOOP_C_16, COMP_LOOP_C_17, COMP_LOOP_C_18, COMP_LOOP_C_19, COMP_LOOP_C_20,
      COMP_LOOP_C_21, COMP_LOOP_C_22, COMP_LOOP_C_23, COMP_LOOP_C_24, COMP_LOOP_C_25,
      COMP_LOOP_C_26, COMP_LOOP_C_27, COMP_LOOP_C_28, COMP_LOOP_C_29, COMP_LOOP_C_30,
      COMP_LOOP_C_31, COMP_LOOP_C_32, COMP_LOOP_C_33, COMP_LOOP_C_34, COMP_LOOP_C_35,
      COMP_LOOP_C_36, COMP_LOOP_C_37, COMP_LOOP_C_38, COMP_LOOP_C_39, COMP_LOOP_C_40,
      COMP_LOOP_C_41, COMP_LOOP_C_42, COMP_LOOP_C_43, COMP_LOOP_C_44, COMP_LOOP_C_45,
      COMP_LOOP_C_46, COMP_LOOP_C_47, COMP_LOOP_C_48, COMP_LOOP_C_49, COMP_LOOP_C_50,
      COMP_LOOP_C_51, COMP_LOOP_C_52, COMP_LOOP_C_53, COMP_LOOP_C_54, COMP_LOOP_C_55,
      COMP_LOOP_C_56, COMP_LOOP_C_57, COMP_LOOP_C_58, COMP_LOOP_C_59, COMP_LOOP_C_60,
      COMP_LOOP_C_61, COMP_LOOP_C_62, COMP_LOOP_C_63, COMP_LOOP_C_64, COMP_LOOP_C_65,
      COMP_LOOP_C_66, COMP_LOOP_C_67, COMP_LOOP_C_68, COMP_LOOP_C_69, COMP_LOOP_C_70,
      COMP_LOOP_C_71, COMP_LOOP_C_72, COMP_LOOP_C_73, COMP_LOOP_C_74, COMP_LOOP_C_75,
      COMP_LOOP_C_76, COMP_LOOP_C_77, COMP_LOOP_C_78, COMP_LOOP_C_79, COMP_LOOP_C_80,
      COMP_LOOP_C_81, COMP_LOOP_C_82, COMP_LOOP_C_83, COMP_LOOP_C_84, COMP_LOOP_C_85,
      COMP_LOOP_C_86, COMP_LOOP_C_87, COMP_LOOP_C_88, COMP_LOOP_C_89, COMP_LOOP_C_90,
      COMP_LOOP_C_91, COMP_LOOP_C_92, COMP_LOOP_C_93, COMP_LOOP_C_94, COMP_LOOP_C_95,
      COMP_LOOP_C_96, COMP_LOOP_C_97, COMP_LOOP_C_98, COMP_LOOP_C_99, COMP_LOOP_C_100,
      COMP_LOOP_C_101, COMP_LOOP_C_102, COMP_LOOP_C_103, COMP_LOOP_C_104, COMP_LOOP_C_105,
      COMP_LOOP_C_106, COMP_LOOP_C_107, COMP_LOOP_C_108, COMP_LOOP_C_109, COMP_LOOP_C_110,
      COMP_LOOP_C_111, COMP_LOOP_C_112, COMP_LOOP_C_113, COMP_LOOP_C_114, COMP_LOOP_C_115,
      COMP_LOOP_C_116, COMP_LOOP_C_117, COMP_LOOP_C_118, COMP_LOOP_C_119, COMP_LOOP_C_120,
      COMP_LOOP_C_121, COMP_LOOP_C_122, COMP_LOOP_C_123, COMP_LOOP_C_124, COMP_LOOP_C_125,
      COMP_LOOP_C_126, COMP_LOOP_C_127, COMP_LOOP_C_128, COMP_LOOP_C_129, COMP_LOOP_C_130,
      COMP_LOOP_C_131, COMP_LOOP_C_132, COMP_LOOP_C_133, COMP_LOOP_C_134, COMP_LOOP_C_135,
      COMP_LOOP_C_136, COMP_LOOP_C_137, COMP_LOOP_C_138, COMP_LOOP_C_139, COMP_LOOP_C_140,
      COMP_LOOP_C_141, COMP_LOOP_C_142, COMP_LOOP_C_143, COMP_LOOP_C_144, COMP_LOOP_C_145,
      COMP_LOOP_C_146, COMP_LOOP_C_147, COMP_LOOP_C_148, COMP_LOOP_C_149, COMP_LOOP_C_150,
      COMP_LOOP_C_151, COMP_LOOP_C_152, COMP_LOOP_C_153, COMP_LOOP_C_154, COMP_LOOP_C_155,
      COMP_LOOP_C_156, COMP_LOOP_C_157, COMP_LOOP_C_158, COMP_LOOP_C_159, COMP_LOOP_C_160,
      COMP_LOOP_C_161, COMP_LOOP_C_162, COMP_LOOP_C_163, COMP_LOOP_C_164, COMP_LOOP_C_165,
      COMP_LOOP_C_166, COMP_LOOP_C_167, COMP_LOOP_C_168, COMP_LOOP_C_169, COMP_LOOP_C_170,
      COMP_LOOP_C_171, COMP_LOOP_C_172, COMP_LOOP_C_173, COMP_LOOP_C_174, COMP_LOOP_C_175,
      COMP_LOOP_C_176, COMP_LOOP_C_177, COMP_LOOP_C_178, COMP_LOOP_C_179, COMP_LOOP_C_180,
      COMP_LOOP_C_181, COMP_LOOP_C_182, COMP_LOOP_C_183, COMP_LOOP_C_184, COMP_LOOP_C_185,
      COMP_LOOP_C_186, COMP_LOOP_C_187, COMP_LOOP_C_188, COMP_LOOP_C_189, COMP_LOOP_C_190,
      COMP_LOOP_C_191, COMP_LOOP_C_192, COMP_LOOP_C_193, COMP_LOOP_C_194, COMP_LOOP_C_195,
      COMP_LOOP_C_196, COMP_LOOP_C_197, COMP_LOOP_C_198, COMP_LOOP_C_199, COMP_LOOP_C_200,
      COMP_LOOP_C_201, COMP_LOOP_C_202, COMP_LOOP_C_203, COMP_LOOP_C_204, COMP_LOOP_C_205,
      COMP_LOOP_C_206, COMP_LOOP_C_207, COMP_LOOP_C_208, COMP_LOOP_C_209, COMP_LOOP_C_210,
      COMP_LOOP_C_211, COMP_LOOP_C_212, COMP_LOOP_C_213, COMP_LOOP_C_214, COMP_LOOP_C_215,
      COMP_LOOP_C_216, COMP_LOOP_C_217, COMP_LOOP_C_218, COMP_LOOP_C_219, COMP_LOOP_C_220,
      COMP_LOOP_C_221, COMP_LOOP_C_222, COMP_LOOP_C_223, COMP_LOOP_C_224, VEC_LOOP_C_0,
      STAGE_LOOP_C_1, main_C_1);

  SIGNAL state_var : inPlaceNTT_DIF_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIF_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIF_core_core_fsm_1 : PROCESS (COMP_LOOP_C_28_tr0, COMP_LOOP_C_56_tr0,
      COMP_LOOP_C_84_tr0, COMP_LOOP_C_112_tr0, COMP_LOOP_C_140_tr0, COMP_LOOP_C_168_tr0,
      COMP_LOOP_C_196_tr0, COMP_LOOP_C_224_tr0, VEC_LOOP_C_0_tr0, STAGE_LOOP_C_1_tr0,
      state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001");
        state_var_NS <= COMP_LOOP_C_0;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011");
        state_var_NS <= COMP_LOOP_C_2;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101");
        state_var_NS <= COMP_LOOP_C_4;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110");
        state_var_NS <= COMP_LOOP_C_5;
      WHEN COMP_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111");
        state_var_NS <= COMP_LOOP_C_6;
      WHEN COMP_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000");
        state_var_NS <= COMP_LOOP_C_7;
      WHEN COMP_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001");
        state_var_NS <= COMP_LOOP_C_8;
      WHEN COMP_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010");
        state_var_NS <= COMP_LOOP_C_9;
      WHEN COMP_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011");
        state_var_NS <= COMP_LOOP_C_10;
      WHEN COMP_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100");
        state_var_NS <= COMP_LOOP_C_11;
      WHEN COMP_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101");
        state_var_NS <= COMP_LOOP_C_12;
      WHEN COMP_LOOP_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110");
        state_var_NS <= COMP_LOOP_C_13;
      WHEN COMP_LOOP_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111");
        state_var_NS <= COMP_LOOP_C_14;
      WHEN COMP_LOOP_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000");
        state_var_NS <= COMP_LOOP_C_15;
      WHEN COMP_LOOP_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001");
        state_var_NS <= COMP_LOOP_C_16;
      WHEN COMP_LOOP_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010");
        state_var_NS <= COMP_LOOP_C_17;
      WHEN COMP_LOOP_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011");
        state_var_NS <= COMP_LOOP_C_18;
      WHEN COMP_LOOP_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100");
        state_var_NS <= COMP_LOOP_C_19;
      WHEN COMP_LOOP_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101");
        state_var_NS <= COMP_LOOP_C_20;
      WHEN COMP_LOOP_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110");
        state_var_NS <= COMP_LOOP_C_21;
      WHEN COMP_LOOP_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111");
        state_var_NS <= COMP_LOOP_C_22;
      WHEN COMP_LOOP_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000");
        state_var_NS <= COMP_LOOP_C_23;
      WHEN COMP_LOOP_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001");
        state_var_NS <= COMP_LOOP_C_24;
      WHEN COMP_LOOP_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010");
        state_var_NS <= COMP_LOOP_C_25;
      WHEN COMP_LOOP_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011");
        state_var_NS <= COMP_LOOP_C_26;
      WHEN COMP_LOOP_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100");
        state_var_NS <= COMP_LOOP_C_27;
      WHEN COMP_LOOP_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101");
        state_var_NS <= COMP_LOOP_C_28;
      WHEN COMP_LOOP_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110");
        IF ( COMP_LOOP_C_28_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_29;
        END IF;
      WHEN COMP_LOOP_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111");
        state_var_NS <= COMP_LOOP_C_30;
      WHEN COMP_LOOP_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000");
        state_var_NS <= COMP_LOOP_C_31;
      WHEN COMP_LOOP_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001");
        state_var_NS <= COMP_LOOP_C_32;
      WHEN COMP_LOOP_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010");
        state_var_NS <= COMP_LOOP_C_33;
      WHEN COMP_LOOP_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011");
        state_var_NS <= COMP_LOOP_C_34;
      WHEN COMP_LOOP_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100");
        state_var_NS <= COMP_LOOP_C_35;
      WHEN COMP_LOOP_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101");
        state_var_NS <= COMP_LOOP_C_36;
      WHEN COMP_LOOP_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110");
        state_var_NS <= COMP_LOOP_C_37;
      WHEN COMP_LOOP_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111");
        state_var_NS <= COMP_LOOP_C_38;
      WHEN COMP_LOOP_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000");
        state_var_NS <= COMP_LOOP_C_39;
      WHEN COMP_LOOP_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001");
        state_var_NS <= COMP_LOOP_C_40;
      WHEN COMP_LOOP_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010");
        state_var_NS <= COMP_LOOP_C_41;
      WHEN COMP_LOOP_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011");
        state_var_NS <= COMP_LOOP_C_42;
      WHEN COMP_LOOP_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100");
        state_var_NS <= COMP_LOOP_C_43;
      WHEN COMP_LOOP_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101");
        state_var_NS <= COMP_LOOP_C_44;
      WHEN COMP_LOOP_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110");
        state_var_NS <= COMP_LOOP_C_45;
      WHEN COMP_LOOP_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111");
        state_var_NS <= COMP_LOOP_C_46;
      WHEN COMP_LOOP_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000");
        state_var_NS <= COMP_LOOP_C_47;
      WHEN COMP_LOOP_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001");
        state_var_NS <= COMP_LOOP_C_48;
      WHEN COMP_LOOP_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010");
        state_var_NS <= COMP_LOOP_C_49;
      WHEN COMP_LOOP_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011");
        state_var_NS <= COMP_LOOP_C_50;
      WHEN COMP_LOOP_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100");
        state_var_NS <= COMP_LOOP_C_51;
      WHEN COMP_LOOP_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101");
        state_var_NS <= COMP_LOOP_C_52;
      WHEN COMP_LOOP_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110");
        state_var_NS <= COMP_LOOP_C_53;
      WHEN COMP_LOOP_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111");
        state_var_NS <= COMP_LOOP_C_54;
      WHEN COMP_LOOP_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000");
        state_var_NS <= COMP_LOOP_C_55;
      WHEN COMP_LOOP_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001");
        state_var_NS <= COMP_LOOP_C_56;
      WHEN COMP_LOOP_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010");
        IF ( COMP_LOOP_C_56_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_57;
        END IF;
      WHEN COMP_LOOP_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011");
        state_var_NS <= COMP_LOOP_C_58;
      WHEN COMP_LOOP_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100");
        state_var_NS <= COMP_LOOP_C_59;
      WHEN COMP_LOOP_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101");
        state_var_NS <= COMP_LOOP_C_60;
      WHEN COMP_LOOP_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110");
        state_var_NS <= COMP_LOOP_C_61;
      WHEN COMP_LOOP_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111");
        state_var_NS <= COMP_LOOP_C_62;
      WHEN COMP_LOOP_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000");
        state_var_NS <= COMP_LOOP_C_63;
      WHEN COMP_LOOP_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001");
        state_var_NS <= COMP_LOOP_C_64;
      WHEN COMP_LOOP_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010");
        state_var_NS <= COMP_LOOP_C_65;
      WHEN COMP_LOOP_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011");
        state_var_NS <= COMP_LOOP_C_66;
      WHEN COMP_LOOP_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100");
        state_var_NS <= COMP_LOOP_C_67;
      WHEN COMP_LOOP_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101");
        state_var_NS <= COMP_LOOP_C_68;
      WHEN COMP_LOOP_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110");
        state_var_NS <= COMP_LOOP_C_69;
      WHEN COMP_LOOP_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111");
        state_var_NS <= COMP_LOOP_C_70;
      WHEN COMP_LOOP_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000");
        state_var_NS <= COMP_LOOP_C_71;
      WHEN COMP_LOOP_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001");
        state_var_NS <= COMP_LOOP_C_72;
      WHEN COMP_LOOP_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010");
        state_var_NS <= COMP_LOOP_C_73;
      WHEN COMP_LOOP_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011");
        state_var_NS <= COMP_LOOP_C_74;
      WHEN COMP_LOOP_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100");
        state_var_NS <= COMP_LOOP_C_75;
      WHEN COMP_LOOP_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101");
        state_var_NS <= COMP_LOOP_C_76;
      WHEN COMP_LOOP_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110");
        state_var_NS <= COMP_LOOP_C_77;
      WHEN COMP_LOOP_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111");
        state_var_NS <= COMP_LOOP_C_78;
      WHEN COMP_LOOP_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000");
        state_var_NS <= COMP_LOOP_C_79;
      WHEN COMP_LOOP_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001");
        state_var_NS <= COMP_LOOP_C_80;
      WHEN COMP_LOOP_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010");
        state_var_NS <= COMP_LOOP_C_81;
      WHEN COMP_LOOP_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011");
        state_var_NS <= COMP_LOOP_C_82;
      WHEN COMP_LOOP_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100");
        state_var_NS <= COMP_LOOP_C_83;
      WHEN COMP_LOOP_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101");
        state_var_NS <= COMP_LOOP_C_84;
      WHEN COMP_LOOP_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110");
        IF ( COMP_LOOP_C_84_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_85;
        END IF;
      WHEN COMP_LOOP_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111");
        state_var_NS <= COMP_LOOP_C_86;
      WHEN COMP_LOOP_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000");
        state_var_NS <= COMP_LOOP_C_87;
      WHEN COMP_LOOP_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001");
        state_var_NS <= COMP_LOOP_C_88;
      WHEN COMP_LOOP_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010");
        state_var_NS <= COMP_LOOP_C_89;
      WHEN COMP_LOOP_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011");
        state_var_NS <= COMP_LOOP_C_90;
      WHEN COMP_LOOP_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100");
        state_var_NS <= COMP_LOOP_C_91;
      WHEN COMP_LOOP_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101");
        state_var_NS <= COMP_LOOP_C_92;
      WHEN COMP_LOOP_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110");
        state_var_NS <= COMP_LOOP_C_93;
      WHEN COMP_LOOP_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111");
        state_var_NS <= COMP_LOOP_C_94;
      WHEN COMP_LOOP_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000");
        state_var_NS <= COMP_LOOP_C_95;
      WHEN COMP_LOOP_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001");
        state_var_NS <= COMP_LOOP_C_96;
      WHEN COMP_LOOP_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010");
        state_var_NS <= COMP_LOOP_C_97;
      WHEN COMP_LOOP_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011");
        state_var_NS <= COMP_LOOP_C_98;
      WHEN COMP_LOOP_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100");
        state_var_NS <= COMP_LOOP_C_99;
      WHEN COMP_LOOP_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101");
        state_var_NS <= COMP_LOOP_C_100;
      WHEN COMP_LOOP_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110");
        state_var_NS <= COMP_LOOP_C_101;
      WHEN COMP_LOOP_C_101 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111");
        state_var_NS <= COMP_LOOP_C_102;
      WHEN COMP_LOOP_C_102 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000");
        state_var_NS <= COMP_LOOP_C_103;
      WHEN COMP_LOOP_C_103 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001");
        state_var_NS <= COMP_LOOP_C_104;
      WHEN COMP_LOOP_C_104 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010");
        state_var_NS <= COMP_LOOP_C_105;
      WHEN COMP_LOOP_C_105 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011");
        state_var_NS <= COMP_LOOP_C_106;
      WHEN COMP_LOOP_C_106 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100");
        state_var_NS <= COMP_LOOP_C_107;
      WHEN COMP_LOOP_C_107 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101");
        state_var_NS <= COMP_LOOP_C_108;
      WHEN COMP_LOOP_C_108 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110");
        state_var_NS <= COMP_LOOP_C_109;
      WHEN COMP_LOOP_C_109 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111");
        state_var_NS <= COMP_LOOP_C_110;
      WHEN COMP_LOOP_C_110 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000");
        state_var_NS <= COMP_LOOP_C_111;
      WHEN COMP_LOOP_C_111 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001");
        state_var_NS <= COMP_LOOP_C_112;
      WHEN COMP_LOOP_C_112 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010");
        IF ( COMP_LOOP_C_112_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_113;
        END IF;
      WHEN COMP_LOOP_C_113 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011");
        state_var_NS <= COMP_LOOP_C_114;
      WHEN COMP_LOOP_C_114 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100");
        state_var_NS <= COMP_LOOP_C_115;
      WHEN COMP_LOOP_C_115 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101");
        state_var_NS <= COMP_LOOP_C_116;
      WHEN COMP_LOOP_C_116 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110");
        state_var_NS <= COMP_LOOP_C_117;
      WHEN COMP_LOOP_C_117 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111");
        state_var_NS <= COMP_LOOP_C_118;
      WHEN COMP_LOOP_C_118 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000");
        state_var_NS <= COMP_LOOP_C_119;
      WHEN COMP_LOOP_C_119 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001");
        state_var_NS <= COMP_LOOP_C_120;
      WHEN COMP_LOOP_C_120 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010");
        state_var_NS <= COMP_LOOP_C_121;
      WHEN COMP_LOOP_C_121 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011");
        state_var_NS <= COMP_LOOP_C_122;
      WHEN COMP_LOOP_C_122 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100");
        state_var_NS <= COMP_LOOP_C_123;
      WHEN COMP_LOOP_C_123 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101");
        state_var_NS <= COMP_LOOP_C_124;
      WHEN COMP_LOOP_C_124 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110");
        state_var_NS <= COMP_LOOP_C_125;
      WHEN COMP_LOOP_C_125 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111");
        state_var_NS <= COMP_LOOP_C_126;
      WHEN COMP_LOOP_C_126 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000");
        state_var_NS <= COMP_LOOP_C_127;
      WHEN COMP_LOOP_C_127 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001");
        state_var_NS <= COMP_LOOP_C_128;
      WHEN COMP_LOOP_C_128 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010");
        state_var_NS <= COMP_LOOP_C_129;
      WHEN COMP_LOOP_C_129 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011");
        state_var_NS <= COMP_LOOP_C_130;
      WHEN COMP_LOOP_C_130 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100");
        state_var_NS <= COMP_LOOP_C_131;
      WHEN COMP_LOOP_C_131 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101");
        state_var_NS <= COMP_LOOP_C_132;
      WHEN COMP_LOOP_C_132 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110");
        state_var_NS <= COMP_LOOP_C_133;
      WHEN COMP_LOOP_C_133 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111");
        state_var_NS <= COMP_LOOP_C_134;
      WHEN COMP_LOOP_C_134 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000");
        state_var_NS <= COMP_LOOP_C_135;
      WHEN COMP_LOOP_C_135 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001");
        state_var_NS <= COMP_LOOP_C_136;
      WHEN COMP_LOOP_C_136 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010");
        state_var_NS <= COMP_LOOP_C_137;
      WHEN COMP_LOOP_C_137 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011");
        state_var_NS <= COMP_LOOP_C_138;
      WHEN COMP_LOOP_C_138 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100");
        state_var_NS <= COMP_LOOP_C_139;
      WHEN COMP_LOOP_C_139 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101");
        state_var_NS <= COMP_LOOP_C_140;
      WHEN COMP_LOOP_C_140 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110");
        IF ( COMP_LOOP_C_140_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_141;
        END IF;
      WHEN COMP_LOOP_C_141 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111");
        state_var_NS <= COMP_LOOP_C_142;
      WHEN COMP_LOOP_C_142 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000");
        state_var_NS <= COMP_LOOP_C_143;
      WHEN COMP_LOOP_C_143 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001");
        state_var_NS <= COMP_LOOP_C_144;
      WHEN COMP_LOOP_C_144 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010");
        state_var_NS <= COMP_LOOP_C_145;
      WHEN COMP_LOOP_C_145 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011");
        state_var_NS <= COMP_LOOP_C_146;
      WHEN COMP_LOOP_C_146 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100");
        state_var_NS <= COMP_LOOP_C_147;
      WHEN COMP_LOOP_C_147 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101");
        state_var_NS <= COMP_LOOP_C_148;
      WHEN COMP_LOOP_C_148 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110");
        state_var_NS <= COMP_LOOP_C_149;
      WHEN COMP_LOOP_C_149 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111");
        state_var_NS <= COMP_LOOP_C_150;
      WHEN COMP_LOOP_C_150 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000");
        state_var_NS <= COMP_LOOP_C_151;
      WHEN COMP_LOOP_C_151 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001");
        state_var_NS <= COMP_LOOP_C_152;
      WHEN COMP_LOOP_C_152 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010");
        state_var_NS <= COMP_LOOP_C_153;
      WHEN COMP_LOOP_C_153 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011");
        state_var_NS <= COMP_LOOP_C_154;
      WHEN COMP_LOOP_C_154 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100");
        state_var_NS <= COMP_LOOP_C_155;
      WHEN COMP_LOOP_C_155 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101");
        state_var_NS <= COMP_LOOP_C_156;
      WHEN COMP_LOOP_C_156 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110");
        state_var_NS <= COMP_LOOP_C_157;
      WHEN COMP_LOOP_C_157 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111");
        state_var_NS <= COMP_LOOP_C_158;
      WHEN COMP_LOOP_C_158 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000");
        state_var_NS <= COMP_LOOP_C_159;
      WHEN COMP_LOOP_C_159 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001");
        state_var_NS <= COMP_LOOP_C_160;
      WHEN COMP_LOOP_C_160 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010");
        state_var_NS <= COMP_LOOP_C_161;
      WHEN COMP_LOOP_C_161 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011");
        state_var_NS <= COMP_LOOP_C_162;
      WHEN COMP_LOOP_C_162 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100");
        state_var_NS <= COMP_LOOP_C_163;
      WHEN COMP_LOOP_C_163 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101");
        state_var_NS <= COMP_LOOP_C_164;
      WHEN COMP_LOOP_C_164 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110");
        state_var_NS <= COMP_LOOP_C_165;
      WHEN COMP_LOOP_C_165 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111");
        state_var_NS <= COMP_LOOP_C_166;
      WHEN COMP_LOOP_C_166 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000");
        state_var_NS <= COMP_LOOP_C_167;
      WHEN COMP_LOOP_C_167 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001");
        state_var_NS <= COMP_LOOP_C_168;
      WHEN COMP_LOOP_C_168 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010");
        IF ( COMP_LOOP_C_168_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_169;
        END IF;
      WHEN COMP_LOOP_C_169 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011");
        state_var_NS <= COMP_LOOP_C_170;
      WHEN COMP_LOOP_C_170 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100");
        state_var_NS <= COMP_LOOP_C_171;
      WHEN COMP_LOOP_C_171 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101");
        state_var_NS <= COMP_LOOP_C_172;
      WHEN COMP_LOOP_C_172 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110");
        state_var_NS <= COMP_LOOP_C_173;
      WHEN COMP_LOOP_C_173 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111");
        state_var_NS <= COMP_LOOP_C_174;
      WHEN COMP_LOOP_C_174 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000");
        state_var_NS <= COMP_LOOP_C_175;
      WHEN COMP_LOOP_C_175 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001");
        state_var_NS <= COMP_LOOP_C_176;
      WHEN COMP_LOOP_C_176 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010");
        state_var_NS <= COMP_LOOP_C_177;
      WHEN COMP_LOOP_C_177 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011");
        state_var_NS <= COMP_LOOP_C_178;
      WHEN COMP_LOOP_C_178 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100");
        state_var_NS <= COMP_LOOP_C_179;
      WHEN COMP_LOOP_C_179 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101");
        state_var_NS <= COMP_LOOP_C_180;
      WHEN COMP_LOOP_C_180 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110");
        state_var_NS <= COMP_LOOP_C_181;
      WHEN COMP_LOOP_C_181 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111");
        state_var_NS <= COMP_LOOP_C_182;
      WHEN COMP_LOOP_C_182 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000");
        state_var_NS <= COMP_LOOP_C_183;
      WHEN COMP_LOOP_C_183 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001");
        state_var_NS <= COMP_LOOP_C_184;
      WHEN COMP_LOOP_C_184 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010");
        state_var_NS <= COMP_LOOP_C_185;
      WHEN COMP_LOOP_C_185 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011");
        state_var_NS <= COMP_LOOP_C_186;
      WHEN COMP_LOOP_C_186 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100");
        state_var_NS <= COMP_LOOP_C_187;
      WHEN COMP_LOOP_C_187 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111101");
        state_var_NS <= COMP_LOOP_C_188;
      WHEN COMP_LOOP_C_188 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111110");
        state_var_NS <= COMP_LOOP_C_189;
      WHEN COMP_LOOP_C_189 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111111");
        state_var_NS <= COMP_LOOP_C_190;
      WHEN COMP_LOOP_C_190 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000000");
        state_var_NS <= COMP_LOOP_C_191;
      WHEN COMP_LOOP_C_191 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000001");
        state_var_NS <= COMP_LOOP_C_192;
      WHEN COMP_LOOP_C_192 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000010");
        state_var_NS <= COMP_LOOP_C_193;
      WHEN COMP_LOOP_C_193 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000011");
        state_var_NS <= COMP_LOOP_C_194;
      WHEN COMP_LOOP_C_194 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000100");
        state_var_NS <= COMP_LOOP_C_195;
      WHEN COMP_LOOP_C_195 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000101");
        state_var_NS <= COMP_LOOP_C_196;
      WHEN COMP_LOOP_C_196 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000110");
        IF ( COMP_LOOP_C_196_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_197;
        END IF;
      WHEN COMP_LOOP_C_197 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11000111");
        state_var_NS <= COMP_LOOP_C_198;
      WHEN COMP_LOOP_C_198 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001000");
        state_var_NS <= COMP_LOOP_C_199;
      WHEN COMP_LOOP_C_199 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001001");
        state_var_NS <= COMP_LOOP_C_200;
      WHEN COMP_LOOP_C_200 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001010");
        state_var_NS <= COMP_LOOP_C_201;
      WHEN COMP_LOOP_C_201 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001011");
        state_var_NS <= COMP_LOOP_C_202;
      WHEN COMP_LOOP_C_202 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001100");
        state_var_NS <= COMP_LOOP_C_203;
      WHEN COMP_LOOP_C_203 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001101");
        state_var_NS <= COMP_LOOP_C_204;
      WHEN COMP_LOOP_C_204 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001110");
        state_var_NS <= COMP_LOOP_C_205;
      WHEN COMP_LOOP_C_205 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11001111");
        state_var_NS <= COMP_LOOP_C_206;
      WHEN COMP_LOOP_C_206 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010000");
        state_var_NS <= COMP_LOOP_C_207;
      WHEN COMP_LOOP_C_207 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010001");
        state_var_NS <= COMP_LOOP_C_208;
      WHEN COMP_LOOP_C_208 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010010");
        state_var_NS <= COMP_LOOP_C_209;
      WHEN COMP_LOOP_C_209 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010011");
        state_var_NS <= COMP_LOOP_C_210;
      WHEN COMP_LOOP_C_210 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010100");
        state_var_NS <= COMP_LOOP_C_211;
      WHEN COMP_LOOP_C_211 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010101");
        state_var_NS <= COMP_LOOP_C_212;
      WHEN COMP_LOOP_C_212 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010110");
        state_var_NS <= COMP_LOOP_C_213;
      WHEN COMP_LOOP_C_213 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11010111");
        state_var_NS <= COMP_LOOP_C_214;
      WHEN COMP_LOOP_C_214 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011000");
        state_var_NS <= COMP_LOOP_C_215;
      WHEN COMP_LOOP_C_215 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011001");
        state_var_NS <= COMP_LOOP_C_216;
      WHEN COMP_LOOP_C_216 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011010");
        state_var_NS <= COMP_LOOP_C_217;
      WHEN COMP_LOOP_C_217 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011011");
        state_var_NS <= COMP_LOOP_C_218;
      WHEN COMP_LOOP_C_218 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011100");
        state_var_NS <= COMP_LOOP_C_219;
      WHEN COMP_LOOP_C_219 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011101");
        state_var_NS <= COMP_LOOP_C_220;
      WHEN COMP_LOOP_C_220 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011110");
        state_var_NS <= COMP_LOOP_C_221;
      WHEN COMP_LOOP_C_221 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11011111");
        state_var_NS <= COMP_LOOP_C_222;
      WHEN COMP_LOOP_C_222 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100000");
        state_var_NS <= COMP_LOOP_C_223;
      WHEN COMP_LOOP_C_223 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100001");
        state_var_NS <= COMP_LOOP_C_224;
      WHEN COMP_LOOP_C_224 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100010");
        IF ( COMP_LOOP_C_224_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100011");
        IF ( VEC_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_1;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100100");
        IF ( STAGE_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "11100101");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS inPlaceNTT_DIF_core_core_fsm_1;

  inPlaceNTT_DIF_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIF_core_core_fsm_1_REG;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core_wait_dp IS
  PORT(
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : OUT STD_LOGIC
  );
END inPlaceNTT_DIF_core_wait_dp;

ARCHITECTURE v14 OF inPlaceNTT_DIF_core_wait_dp IS
  -- Default Constants

BEGIN
  COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en <= ensig_cgo OR ensig_cgo_iro;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_32_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_33_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_34_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_35_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_36_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_37_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_38_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_39_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_40_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_41_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_42_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_43_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_44_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_45_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_46_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_47_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_48_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_49_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_50_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_51_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_52_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_53_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_54_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_55_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_56_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_57_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_58_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_59_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_60_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_61_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_62_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_63_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_32_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_33_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_34_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_35_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_36_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_37_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_38_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_39_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_40_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_41_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_42_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_43_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_44_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_45_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_46_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_47_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_48_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_49_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_50_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_51_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_52_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_53_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_54_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_55_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_56_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_57_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_58_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_59_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_60_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_61_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_62_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_0_63_lz : OUT STD_LOGIC;
    vec_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_32_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_33_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_34_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_35_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_36_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_37_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_38_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_39_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_40_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_41_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_42_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_43_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_44_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_45_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_46_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_47_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_48_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_49_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_50_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_51_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_52_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_53_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_54_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_55_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_56_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_57_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_58_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_59_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_60_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_61_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_62_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_63_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_32_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_33_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_34_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_35_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_36_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_37_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_38_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_39_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_40_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_41_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_42_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_43_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_44_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_45_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_46_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_47_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_48_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_49_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_50_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_51_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_52_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_53_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_54_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_55_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_56_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_57_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_58_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_59_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_60_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_61_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_62_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_rsc_0_63_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_1_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_2_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_3_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_4_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_5_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_6_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_7_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_8_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_9_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_10_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_11_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_12_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_13_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_14_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_15_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_16_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_17_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_18_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_19_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_20_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_21_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_22_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_23_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_24_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_25_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_26_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_27_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_28_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_29_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_30_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_31_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_32_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_33_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_34_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_35_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_36_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_37_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_38_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_39_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_40_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_41_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_42_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_43_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_44_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_45_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_46_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_47_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_48_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_49_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_50_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_51_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_52_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_53_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_54_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_55_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_56_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_57_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_58_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_59_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_60_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_61_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_62_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_63_i_we_d_pff : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
  );
END inPlaceNTT_DIF_core;

ARCHITECTURE v14 OF inPlaceNTT_DIF_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : STD_LOGIC;
  SIGNAL fsm_output : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL nor_tmp_1 : STD_LOGIC;
  SIGNAL mux_tmp_6 : STD_LOGIC;
  SIGNAL and_dcpl_8 : STD_LOGIC;
  SIGNAL and_tmp_10 : STD_LOGIC;
  SIGNAL or_tmp_105 : STD_LOGIC;
  SIGNAL or_tmp_118 : STD_LOGIC;
  SIGNAL or_tmp_119 : STD_LOGIC;
  SIGNAL not_tmp_88 : STD_LOGIC;
  SIGNAL nor_tmp_99 : STD_LOGIC;
  SIGNAL mux_tmp_206 : STD_LOGIC;
  SIGNAL mux_tmp_293 : STD_LOGIC;
  SIGNAL mux_tmp_444 : STD_LOGIC;
  SIGNAL or_tmp_404 : STD_LOGIC;
  SIGNAL mux_tmp_656 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_59 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL and_dcpl_64 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_tmp_29 : STD_LOGIC;
  SIGNAL mux_tmp_720 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_73 : STD_LOGIC;
  SIGNAL and_dcpl_74 : STD_LOGIC;
  SIGNAL and_dcpl_75 : STD_LOGIC;
  SIGNAL and_dcpl_76 : STD_LOGIC;
  SIGNAL and_dcpl_77 : STD_LOGIC;
  SIGNAL and_dcpl_78 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL and_dcpl_80 : STD_LOGIC;
  SIGNAL and_dcpl_81 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_86 : STD_LOGIC;
  SIGNAL and_dcpl_87 : STD_LOGIC;
  SIGNAL and_dcpl_88 : STD_LOGIC;
  SIGNAL and_dcpl_90 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_95 : STD_LOGIC;
  SIGNAL and_dcpl_96 : STD_LOGIC;
  SIGNAL and_dcpl_97 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_101 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_106 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_113 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_116 : STD_LOGIC;
  SIGNAL and_dcpl_118 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL or_tmp_491 : STD_LOGIC;
  SIGNAL or_tmp_495 : STD_LOGIC;
  SIGNAL or_tmp_497 : STD_LOGIC;
  SIGNAL or_tmp_501 : STD_LOGIC;
  SIGNAL or_tmp_535 : STD_LOGIC;
  SIGNAL or_tmp_539 : STD_LOGIC;
  SIGNAL or_tmp_541 : STD_LOGIC;
  SIGNAL or_tmp_545 : STD_LOGIC;
  SIGNAL not_tmp_321 : STD_LOGIC;
  SIGNAL or_tmp_579 : STD_LOGIC;
  SIGNAL or_tmp_583 : STD_LOGIC;
  SIGNAL or_tmp_585 : STD_LOGIC;
  SIGNAL or_tmp_589 : STD_LOGIC;
  SIGNAL or_tmp_623 : STD_LOGIC;
  SIGNAL or_tmp_627 : STD_LOGIC;
  SIGNAL or_tmp_629 : STD_LOGIC;
  SIGNAL or_tmp_633 : STD_LOGIC;
  SIGNAL not_tmp_330 : STD_LOGIC;
  SIGNAL or_tmp_667 : STD_LOGIC;
  SIGNAL or_tmp_671 : STD_LOGIC;
  SIGNAL or_tmp_673 : STD_LOGIC;
  SIGNAL or_tmp_677 : STD_LOGIC;
  SIGNAL or_tmp_711 : STD_LOGIC;
  SIGNAL or_tmp_715 : STD_LOGIC;
  SIGNAL or_tmp_717 : STD_LOGIC;
  SIGNAL or_tmp_721 : STD_LOGIC;
  SIGNAL or_tmp_755 : STD_LOGIC;
  SIGNAL or_tmp_759 : STD_LOGIC;
  SIGNAL or_tmp_761 : STD_LOGIC;
  SIGNAL or_tmp_765 : STD_LOGIC;
  SIGNAL or_tmp_799 : STD_LOGIC;
  SIGNAL or_tmp_803 : STD_LOGIC;
  SIGNAL or_tmp_805 : STD_LOGIC;
  SIGNAL or_tmp_809 : STD_LOGIC;
  SIGNAL not_tmp_347 : STD_LOGIC;
  SIGNAL or_tmp_843 : STD_LOGIC;
  SIGNAL or_tmp_847 : STD_LOGIC;
  SIGNAL or_tmp_849 : STD_LOGIC;
  SIGNAL or_tmp_853 : STD_LOGIC;
  SIGNAL or_tmp_887 : STD_LOGIC;
  SIGNAL or_tmp_891 : STD_LOGIC;
  SIGNAL or_tmp_893 : STD_LOGIC;
  SIGNAL or_tmp_897 : STD_LOGIC;
  SIGNAL or_tmp_931 : STD_LOGIC;
  SIGNAL or_tmp_935 : STD_LOGIC;
  SIGNAL or_tmp_937 : STD_LOGIC;
  SIGNAL or_tmp_941 : STD_LOGIC;
  SIGNAL or_tmp_975 : STD_LOGIC;
  SIGNAL or_tmp_979 : STD_LOGIC;
  SIGNAL or_tmp_981 : STD_LOGIC;
  SIGNAL or_tmp_985 : STD_LOGIC;
  SIGNAL or_tmp_1019 : STD_LOGIC;
  SIGNAL or_tmp_1023 : STD_LOGIC;
  SIGNAL or_tmp_1025 : STD_LOGIC;
  SIGNAL or_tmp_1029 : STD_LOGIC;
  SIGNAL or_tmp_1063 : STD_LOGIC;
  SIGNAL or_tmp_1067 : STD_LOGIC;
  SIGNAL or_tmp_1069 : STD_LOGIC;
  SIGNAL or_tmp_1073 : STD_LOGIC;
  SIGNAL or_tmp_1107 : STD_LOGIC;
  SIGNAL or_tmp_1111 : STD_LOGIC;
  SIGNAL or_tmp_1113 : STD_LOGIC;
  SIGNAL or_tmp_1117 : STD_LOGIC;
  SIGNAL or_tmp_1151 : STD_LOGIC;
  SIGNAL or_tmp_1155 : STD_LOGIC;
  SIGNAL or_tmp_1157 : STD_LOGIC;
  SIGNAL or_tmp_1161 : STD_LOGIC;
  SIGNAL or_tmp_1195 : STD_LOGIC;
  SIGNAL or_tmp_1199 : STD_LOGIC;
  SIGNAL or_tmp_1201 : STD_LOGIC;
  SIGNAL or_tmp_1205 : STD_LOGIC;
  SIGNAL not_tmp_384 : STD_LOGIC;
  SIGNAL not_tmp_388 : STD_LOGIC;
  SIGNAL or_tmp_1239 : STD_LOGIC;
  SIGNAL or_tmp_1243 : STD_LOGIC;
  SIGNAL or_tmp_1245 : STD_LOGIC;
  SIGNAL or_tmp_1249 : STD_LOGIC;
  SIGNAL or_tmp_1283 : STD_LOGIC;
  SIGNAL or_tmp_1287 : STD_LOGIC;
  SIGNAL or_tmp_1289 : STD_LOGIC;
  SIGNAL or_tmp_1293 : STD_LOGIC;
  SIGNAL or_tmp_1327 : STD_LOGIC;
  SIGNAL or_tmp_1331 : STD_LOGIC;
  SIGNAL or_tmp_1333 : STD_LOGIC;
  SIGNAL or_tmp_1337 : STD_LOGIC;
  SIGNAL or_tmp_1371 : STD_LOGIC;
  SIGNAL or_tmp_1375 : STD_LOGIC;
  SIGNAL or_tmp_1377 : STD_LOGIC;
  SIGNAL or_tmp_1381 : STD_LOGIC;
  SIGNAL or_tmp_1415 : STD_LOGIC;
  SIGNAL or_tmp_1419 : STD_LOGIC;
  SIGNAL or_tmp_1421 : STD_LOGIC;
  SIGNAL or_tmp_1425 : STD_LOGIC;
  SIGNAL or_tmp_1459 : STD_LOGIC;
  SIGNAL or_tmp_1463 : STD_LOGIC;
  SIGNAL or_tmp_1465 : STD_LOGIC;
  SIGNAL or_tmp_1469 : STD_LOGIC;
  SIGNAL or_tmp_1503 : STD_LOGIC;
  SIGNAL or_tmp_1507 : STD_LOGIC;
  SIGNAL or_tmp_1509 : STD_LOGIC;
  SIGNAL or_tmp_1513 : STD_LOGIC;
  SIGNAL not_tmp_414 : STD_LOGIC;
  SIGNAL or_tmp_1547 : STD_LOGIC;
  SIGNAL or_tmp_1551 : STD_LOGIC;
  SIGNAL or_tmp_1553 : STD_LOGIC;
  SIGNAL or_tmp_1557 : STD_LOGIC;
  SIGNAL or_tmp_1591 : STD_LOGIC;
  SIGNAL or_tmp_1595 : STD_LOGIC;
  SIGNAL or_tmp_1597 : STD_LOGIC;
  SIGNAL or_tmp_1601 : STD_LOGIC;
  SIGNAL or_tmp_1635 : STD_LOGIC;
  SIGNAL or_tmp_1639 : STD_LOGIC;
  SIGNAL or_tmp_1641 : STD_LOGIC;
  SIGNAL or_tmp_1645 : STD_LOGIC;
  SIGNAL or_tmp_1679 : STD_LOGIC;
  SIGNAL or_tmp_1683 : STD_LOGIC;
  SIGNAL or_tmp_1685 : STD_LOGIC;
  SIGNAL or_tmp_1689 : STD_LOGIC;
  SIGNAL or_tmp_1723 : STD_LOGIC;
  SIGNAL or_tmp_1727 : STD_LOGIC;
  SIGNAL or_tmp_1729 : STD_LOGIC;
  SIGNAL or_tmp_1733 : STD_LOGIC;
  SIGNAL or_tmp_1767 : STD_LOGIC;
  SIGNAL or_tmp_1771 : STD_LOGIC;
  SIGNAL or_tmp_1773 : STD_LOGIC;
  SIGNAL or_tmp_1777 : STD_LOGIC;
  SIGNAL or_tmp_1811 : STD_LOGIC;
  SIGNAL or_tmp_1815 : STD_LOGIC;
  SIGNAL or_tmp_1817 : STD_LOGIC;
  SIGNAL or_tmp_1821 : STD_LOGIC;
  SIGNAL or_tmp_1855 : STD_LOGIC;
  SIGNAL or_tmp_1859 : STD_LOGIC;
  SIGNAL or_tmp_1861 : STD_LOGIC;
  SIGNAL or_tmp_1865 : STD_LOGIC;
  SIGNAL or_tmp_1898 : STD_LOGIC;
  SIGNAL or_tmp_1902 : STD_LOGIC;
  SIGNAL or_tmp_1904 : STD_LOGIC;
  SIGNAL not_tmp_452 : STD_LOGIC;
  SIGNAL not_tmp_453 : STD_LOGIC;
  SIGNAL or_tmp_1908 : STD_LOGIC;
  SIGNAL or_tmp_1942 : STD_LOGIC;
  SIGNAL or_tmp_1946 : STD_LOGIC;
  SIGNAL or_tmp_1948 : STD_LOGIC;
  SIGNAL not_tmp_458 : STD_LOGIC;
  SIGNAL or_tmp_1952 : STD_LOGIC;
  SIGNAL or_tmp_1986 : STD_LOGIC;
  SIGNAL or_tmp_1990 : STD_LOGIC;
  SIGNAL or_tmp_1992 : STD_LOGIC;
  SIGNAL or_tmp_1996 : STD_LOGIC;
  SIGNAL or_tmp_2030 : STD_LOGIC;
  SIGNAL or_tmp_2034 : STD_LOGIC;
  SIGNAL or_tmp_2036 : STD_LOGIC;
  SIGNAL not_tmp_467 : STD_LOGIC;
  SIGNAL or_tmp_2040 : STD_LOGIC;
  SIGNAL or_tmp_2074 : STD_LOGIC;
  SIGNAL or_tmp_2078 : STD_LOGIC;
  SIGNAL or_tmp_2080 : STD_LOGIC;
  SIGNAL or_tmp_2084 : STD_LOGIC;
  SIGNAL or_tmp_2118 : STD_LOGIC;
  SIGNAL or_tmp_2122 : STD_LOGIC;
  SIGNAL or_tmp_2124 : STD_LOGIC;
  SIGNAL or_tmp_2128 : STD_LOGIC;
  SIGNAL or_tmp_2162 : STD_LOGIC;
  SIGNAL or_tmp_2166 : STD_LOGIC;
  SIGNAL or_tmp_2168 : STD_LOGIC;
  SIGNAL or_tmp_2172 : STD_LOGIC;
  SIGNAL or_tmp_2206 : STD_LOGIC;
  SIGNAL or_tmp_2210 : STD_LOGIC;
  SIGNAL or_tmp_2212 : STD_LOGIC;
  SIGNAL not_tmp_484 : STD_LOGIC;
  SIGNAL or_tmp_2216 : STD_LOGIC;
  SIGNAL or_tmp_2250 : STD_LOGIC;
  SIGNAL or_tmp_2254 : STD_LOGIC;
  SIGNAL or_tmp_2256 : STD_LOGIC;
  SIGNAL or_tmp_2260 : STD_LOGIC;
  SIGNAL or_tmp_2294 : STD_LOGIC;
  SIGNAL or_tmp_2298 : STD_LOGIC;
  SIGNAL or_tmp_2300 : STD_LOGIC;
  SIGNAL or_tmp_2304 : STD_LOGIC;
  SIGNAL or_tmp_2338 : STD_LOGIC;
  SIGNAL or_tmp_2342 : STD_LOGIC;
  SIGNAL or_tmp_2344 : STD_LOGIC;
  SIGNAL or_tmp_2348 : STD_LOGIC;
  SIGNAL or_tmp_2382 : STD_LOGIC;
  SIGNAL or_tmp_2386 : STD_LOGIC;
  SIGNAL or_tmp_2388 : STD_LOGIC;
  SIGNAL or_tmp_2392 : STD_LOGIC;
  SIGNAL or_tmp_2426 : STD_LOGIC;
  SIGNAL or_tmp_2430 : STD_LOGIC;
  SIGNAL or_tmp_2432 : STD_LOGIC;
  SIGNAL or_tmp_2436 : STD_LOGIC;
  SIGNAL or_tmp_2470 : STD_LOGIC;
  SIGNAL or_tmp_2474 : STD_LOGIC;
  SIGNAL or_tmp_2476 : STD_LOGIC;
  SIGNAL or_tmp_2480 : STD_LOGIC;
  SIGNAL or_tmp_2514 : STD_LOGIC;
  SIGNAL or_tmp_2518 : STD_LOGIC;
  SIGNAL or_tmp_2520 : STD_LOGIC;
  SIGNAL or_tmp_2524 : STD_LOGIC;
  SIGNAL or_tmp_2558 : STD_LOGIC;
  SIGNAL or_tmp_2562 : STD_LOGIC;
  SIGNAL or_tmp_2564 : STD_LOGIC;
  SIGNAL or_tmp_2567 : STD_LOGIC;
  SIGNAL or_tmp_2601 : STD_LOGIC;
  SIGNAL or_tmp_2605 : STD_LOGIC;
  SIGNAL or_tmp_2607 : STD_LOGIC;
  SIGNAL not_tmp_522 : STD_LOGIC;
  SIGNAL or_tmp_2611 : STD_LOGIC;
  SIGNAL not_tmp_523 : STD_LOGIC;
  SIGNAL not_tmp_527 : STD_LOGIC;
  SIGNAL or_tmp_2645 : STD_LOGIC;
  SIGNAL or_tmp_2649 : STD_LOGIC;
  SIGNAL or_tmp_2651 : STD_LOGIC;
  SIGNAL or_tmp_2655 : STD_LOGIC;
  SIGNAL or_tmp_2689 : STD_LOGIC;
  SIGNAL or_tmp_2693 : STD_LOGIC;
  SIGNAL or_tmp_2695 : STD_LOGIC;
  SIGNAL or_tmp_2699 : STD_LOGIC;
  SIGNAL or_tmp_2733 : STD_LOGIC;
  SIGNAL or_tmp_2737 : STD_LOGIC;
  SIGNAL or_tmp_2739 : STD_LOGIC;
  SIGNAL or_tmp_2743 : STD_LOGIC;
  SIGNAL or_tmp_2777 : STD_LOGIC;
  SIGNAL or_tmp_2781 : STD_LOGIC;
  SIGNAL or_tmp_2783 : STD_LOGIC;
  SIGNAL or_tmp_2787 : STD_LOGIC;
  SIGNAL not_tmp_544 : STD_LOGIC;
  SIGNAL or_tmp_2821 : STD_LOGIC;
  SIGNAL or_tmp_2825 : STD_LOGIC;
  SIGNAL or_tmp_2827 : STD_LOGIC;
  SIGNAL or_tmp_2831 : STD_LOGIC;
  SIGNAL not_tmp_549 : STD_LOGIC;
  SIGNAL or_tmp_2865 : STD_LOGIC;
  SIGNAL or_tmp_2869 : STD_LOGIC;
  SIGNAL or_tmp_2871 : STD_LOGIC;
  SIGNAL or_tmp_2875 : STD_LOGIC;
  SIGNAL or_tmp_2909 : STD_LOGIC;
  SIGNAL or_tmp_2913 : STD_LOGIC;
  SIGNAL or_tmp_2915 : STD_LOGIC;
  SIGNAL or_tmp_2919 : STD_LOGIC;
  SIGNAL or_tmp_2953 : STD_LOGIC;
  SIGNAL or_tmp_2957 : STD_LOGIC;
  SIGNAL or_tmp_2959 : STD_LOGIC;
  SIGNAL not_tmp_559 : STD_LOGIC;
  SIGNAL or_tmp_2963 : STD_LOGIC;
  SIGNAL not_tmp_560 : STD_LOGIC;
  SIGNAL or_tmp_2997 : STD_LOGIC;
  SIGNAL or_tmp_3001 : STD_LOGIC;
  SIGNAL or_tmp_3003 : STD_LOGIC;
  SIGNAL not_tmp_565 : STD_LOGIC;
  SIGNAL or_tmp_3007 : STD_LOGIC;
  SIGNAL or_tmp_3041 : STD_LOGIC;
  SIGNAL or_tmp_3045 : STD_LOGIC;
  SIGNAL or_tmp_3047 : STD_LOGIC;
  SIGNAL or_tmp_3051 : STD_LOGIC;
  SIGNAL not_tmp_570 : STD_LOGIC;
  SIGNAL or_tmp_3085 : STD_LOGIC;
  SIGNAL or_tmp_3089 : STD_LOGIC;
  SIGNAL or_tmp_3091 : STD_LOGIC;
  SIGNAL not_tmp_575 : STD_LOGIC;
  SIGNAL or_tmp_3094 : STD_LOGIC;
  SIGNAL or_tmp_3128 : STD_LOGIC;
  SIGNAL or_tmp_3132 : STD_LOGIC;
  SIGNAL or_tmp_3134 : STD_LOGIC;
  SIGNAL or_tmp_3138 : STD_LOGIC;
  SIGNAL or_tmp_3172 : STD_LOGIC;
  SIGNAL or_tmp_3176 : STD_LOGIC;
  SIGNAL or_tmp_3178 : STD_LOGIC;
  SIGNAL or_tmp_3182 : STD_LOGIC;
  SIGNAL or_tmp_3215 : STD_LOGIC;
  SIGNAL or_tmp_3219 : STD_LOGIC;
  SIGNAL or_tmp_3221 : STD_LOGIC;
  SIGNAL or_tmp_3225 : STD_LOGIC;
  SIGNAL or_tmp_3258 : STD_LOGIC;
  SIGNAL or_tmp_3262 : STD_LOGIC;
  SIGNAL or_tmp_3264 : STD_LOGIC;
  SIGNAL nor_tmp_306 : STD_LOGIC;
  SIGNAL nor_tmp_307 : STD_LOGIC;
  SIGNAL and_dcpl_258 : STD_LOGIC;
  SIGNAL and_dcpl_259 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL and_dcpl_261 : STD_LOGIC;
  SIGNAL and_dcpl_262 : STD_LOGIC;
  SIGNAL and_dcpl_263 : STD_LOGIC;
  SIGNAL and_dcpl_264 : STD_LOGIC;
  SIGNAL and_dcpl_265 : STD_LOGIC;
  SIGNAL and_dcpl_268 : STD_LOGIC;
  SIGNAL mux_tmp_2924 : STD_LOGIC;
  SIGNAL or_tmp_3717 : STD_LOGIC;
  SIGNAL mux_tmp_2927 : STD_LOGIC;
  SIGNAL or_tmp_3718 : STD_LOGIC;
  SIGNAL and_dcpl_340 : STD_LOGIC;
  SIGNAL or_tmp_3721 : STD_LOGIC;
  SIGNAL and_dcpl_343 : STD_LOGIC;
  SIGNAL and_dcpl_344 : STD_LOGIC;
  SIGNAL and_dcpl_346 : STD_LOGIC;
  SIGNAL and_dcpl_347 : STD_LOGIC;
  SIGNAL and_dcpl_349 : STD_LOGIC;
  SIGNAL and_dcpl_351 : STD_LOGIC;
  SIGNAL and_dcpl_353 : STD_LOGIC;
  SIGNAL and_dcpl_354 : STD_LOGIC;
  SIGNAL and_dcpl_355 : STD_LOGIC;
  SIGNAL and_dcpl_357 : STD_LOGIC;
  SIGNAL and_dcpl_359 : STD_LOGIC;
  SIGNAL nand_tmp_142 : STD_LOGIC;
  SIGNAL mux_tmp_2939 : STD_LOGIC;
  SIGNAL or_tmp_3734 : STD_LOGIC;
  SIGNAL and_dcpl_365 : STD_LOGIC;
  SIGNAL or_dcpl_122 : STD_LOGIC;
  SIGNAL or_dcpl_125 : STD_LOGIC;
  SIGNAL mux_tmp_2953 : STD_LOGIC;
  SIGNAL mux_tmp_2955 : STD_LOGIC;
  SIGNAL mux_tmp_2956 : STD_LOGIC;
  SIGNAL mux_tmp_2959 : STD_LOGIC;
  SIGNAL mux_tmp_2960 : STD_LOGIC;
  SIGNAL mux_tmp_2961 : STD_LOGIC;
  SIGNAL mux_tmp_2965 : STD_LOGIC;
  SIGNAL mux_tmp_2966 : STD_LOGIC;
  SIGNAL mux_tmp_2968 : STD_LOGIC;
  SIGNAL and_dcpl_370 : STD_LOGIC;
  SIGNAL mux_tmp_2971 : STD_LOGIC;
  SIGNAL or_tmp_3744 : STD_LOGIC;
  SIGNAL mux_tmp_2975 : STD_LOGIC;
  SIGNAL or_tmp_3746 : STD_LOGIC;
  SIGNAL mux_tmp_2976 : STD_LOGIC;
  SIGNAL and_dcpl_375 : STD_LOGIC;
  SIGNAL or_tmp_3747 : STD_LOGIC;
  SIGNAL and_dcpl_377 : STD_LOGIC;
  SIGNAL and_dcpl_382 : STD_LOGIC;
  SIGNAL and_dcpl_384 : STD_LOGIC;
  SIGNAL mux_tmp_2993 : STD_LOGIC;
  SIGNAL mux_tmp_2994 : STD_LOGIC;
  SIGNAL or_tmp_3757 : STD_LOGIC;
  SIGNAL or_tmp_3760 : STD_LOGIC;
  SIGNAL mux_tmp_3001 : STD_LOGIC;
  SIGNAL mux_tmp_3003 : STD_LOGIC;
  SIGNAL mux_tmp_3009 : STD_LOGIC;
  SIGNAL mux_tmp_3012 : STD_LOGIC;
  SIGNAL mux_tmp_3013 : STD_LOGIC;
  SIGNAL mux_tmp_3016 : STD_LOGIC;
  SIGNAL and_dcpl_387 : STD_LOGIC;
  SIGNAL or_tmp_3773 : STD_LOGIC;
  SIGNAL and_dcpl_388 : STD_LOGIC;
  SIGNAL mux_tmp_3042 : STD_LOGIC;
  SIGNAL and_tmp_31 : STD_LOGIC;
  SIGNAL mux_tmp_3049 : STD_LOGIC;
  SIGNAL and_dcpl_390 : STD_LOGIC;
  SIGNAL and_dcpl_392 : STD_LOGIC;
  SIGNAL and_dcpl_396 : STD_LOGIC;
  SIGNAL and_dcpl_399 : STD_LOGIC;
  SIGNAL and_dcpl_402 : STD_LOGIC;
  SIGNAL mux_tmp_3069 : STD_LOGIC;
  SIGNAL mux_tmp_3070 : STD_LOGIC;
  SIGNAL mux_tmp_3078 : STD_LOGIC;
  SIGNAL and_dcpl_403 : STD_LOGIC;
  SIGNAL and_dcpl_404 : STD_LOGIC;
  SIGNAL and_dcpl_406 : STD_LOGIC;
  SIGNAL and_dcpl_407 : STD_LOGIC;
  SIGNAL mux_tmp_3098 : STD_LOGIC;
  SIGNAL mux_tmp_3100 : STD_LOGIC;
  SIGNAL mux_tmp_3101 : STD_LOGIC;
  SIGNAL mux_tmp_3102 : STD_LOGIC;
  SIGNAL and_dcpl_410 : STD_LOGIC;
  SIGNAL and_dcpl_411 : STD_LOGIC;
  SIGNAL mux_tmp_3119 : STD_LOGIC;
  SIGNAL not_tmp_811 : STD_LOGIC;
  SIGNAL mux_tmp_3133 : STD_LOGIC;
  SIGNAL or_tmp_3801 : STD_LOGIC;
  SIGNAL and_tmp_33 : STD_LOGIC;
  SIGNAL and_dcpl_421 : STD_LOGIC;
  SIGNAL mux_tmp_3169 : STD_LOGIC;
  SIGNAL mux_tmp_3193 : STD_LOGIC;
  SIGNAL mux_tmp_3196 : STD_LOGIC;
  SIGNAL and_tmp_35 : STD_LOGIC;
  SIGNAL mux_tmp_3210 : STD_LOGIC;
  SIGNAL and_tmp_36 : STD_LOGIC;
  SIGNAL mux_tmp_3213 : STD_LOGIC;
  SIGNAL mux_tmp_3214 : STD_LOGIC;
  SIGNAL mux_tmp_3218 : STD_LOGIC;
  SIGNAL or_dcpl_134 : STD_LOGIC;
  SIGNAL and_dcpl_432 : STD_LOGIC;
  SIGNAL or_tmp_3833 : STD_LOGIC;
  SIGNAL nor_tmp_391 : STD_LOGIC;
  SIGNAL mux_tmp_3280 : STD_LOGIC;
  SIGNAL not_tmp_868 : STD_LOGIC;
  SIGNAL or_dcpl_150 : STD_LOGIC;
  SIGNAL mux_tmp_3288 : STD_LOGIC;
  SIGNAL COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_14_psp_sva_1 : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL VEC_LOOP_j_10_0_sva_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_k_10_3_sva_6_0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_315_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_289_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_313_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_326_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_319_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_521_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_767_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_760_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_734_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_970_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_969_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_984_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_964_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_961_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_955_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_962_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_957_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_976_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_958_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_998_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_972_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_987_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_985_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_991_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1185_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1211_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1209_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1196_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1208_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1186_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1182_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1222_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1188_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1215_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1194_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1193_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1435_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1446_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1439_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1420_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1432_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1424_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1410_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1403_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1663_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1659_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1633_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1642_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1648_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1630_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1670_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1629_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_2_tmp_mul_idiv_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_2_tmp_lshift_ncse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_3_tmp_lshift_ncse_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_206_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_151_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_119_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_109_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1106_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_102_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_117_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1370_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_122_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_1_cse_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_3_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_14_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_7_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_psp_sva : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_1_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_13_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_5_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_5_tmp_mul_idiv_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_psp_sva_mx0w0 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva_1 : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_274_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_276_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_280_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_288_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_304_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_243_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_245_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_249_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_257_rgt : STD_LOGIC;
  SIGNAL mux_3360_tmp : STD_LOGIC;
  SIGNAL and_478_m1c : STD_LOGIC;
  SIGNAL nor_tmp_396 : STD_LOGIC;
  SIGNAL and_476_tmp : STD_LOGIC;
  SIGNAL nor_1579_tmp : STD_LOGIC;
  SIGNAL and_474_tmp : STD_LOGIC;
  SIGNAL reg_COMP_LOOP_k_10_3_ftd : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL nand_191_cse : STD_LOGIC;
  SIGNAL nand_190_cse : STD_LOGIC;
  SIGNAL nand_188_cse : STD_LOGIC;
  SIGNAL nand_174_cse : STD_LOGIC;
  SIGNAL nand_175_cse : STD_LOGIC;
  SIGNAL nand_184_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_0_63_obj_ld_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL or_595_cse : STD_LOGIC;
  SIGNAL and_507_cse : STD_LOGIC;
  SIGNAL or_341_cse : STD_LOGIC;
  SIGNAL or_359_cse : STD_LOGIC;
  SIGNAL mux_297_cse : STD_LOGIC;
  SIGNAL or_4057_cse : STD_LOGIC;
  SIGNAL and_677_cse : STD_LOGIC;
  SIGNAL nor_358_cse : STD_LOGIC;
  SIGNAL nor_412_cse : STD_LOGIC;
  SIGNAL and_493_cse : STD_LOGIC;
  SIGNAL and_640_cse : STD_LOGIC;
  SIGNAL or_564_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_5_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_36_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_43_cse : STD_LOGIC;
  SIGNAL nor_399_cse : STD_LOGIC;
  SIGNAL or_4007_cse : STD_LOGIC;
  SIGNAL or_80_cse : STD_LOGIC;
  SIGNAL and_705_cse : STD_LOGIC;
  SIGNAL nor_1683_cse : STD_LOGIC;
  SIGNAL and_673_cse : STD_LOGIC;
  SIGNAL and_639_cse : STD_LOGIC;
  SIGNAL and_735_cse : STD_LOGIC;
  SIGNAL or_364_cse : STD_LOGIC;
  SIGNAL and_763_cse : STD_LOGIC;
  SIGNAL or_477_cse : STD_LOGIC;
  SIGNAL nor_1674_cse : STD_LOGIC;
  SIGNAL and_808_cse : STD_LOGIC;
  SIGNAL or_150_cse : STD_LOGIC;
  SIGNAL nor_398_cse : STD_LOGIC;
  SIGNAL mux_742_cse : STD_LOGIC;
  SIGNAL and_779_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm : STD_LOGIC;
  SIGNAL and_655_cse : STD_LOGIC;
  SIGNAL or_4050_cse : STD_LOGIC;
  SIGNAL and_78_cse : STD_LOGIC;
  SIGNAL mux_180_cse : STD_LOGIC;
  SIGNAL mux_221_cse : STD_LOGIC;
  SIGNAL and_736_cse : STD_LOGIC;
  SIGNAL mux_3095_cse : STD_LOGIC;
  SIGNAL mux_2997_rmff : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_8_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_1_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_2_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_3_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_4_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_5_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_mux1h_6_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_3025_itm : STD_LOGIC;
  SIGNAL mux_3058_itm : STD_LOGIC;
  SIGNAL mux_3114_itm : STD_LOGIC;
  SIGNAL mux_3175_itm : STD_LOGIC;
  SIGNAL mux_3185_itm : STD_LOGIC;
  SIGNAL mux_3187_itm : STD_LOGIC;
  SIGNAL mux_3201_itm : STD_LOGIC;
  SIGNAL mux_3305_itm : STD_LOGIC;
  SIGNAL z_out : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL and_dcpl_477 : STD_LOGIC;
  SIGNAL and_dcpl_488 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL and_dcpl_501 : STD_LOGIC;
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_dcpl_503 : STD_LOGIC;
  SIGNAL and_dcpl_509 : STD_LOGIC;
  SIGNAL and_dcpl_513 : STD_LOGIC;
  SIGNAL and_dcpl_514 : STD_LOGIC;
  SIGNAL and_dcpl_519 : STD_LOGIC;
  SIGNAL and_dcpl_526 : STD_LOGIC;
  SIGNAL and_dcpl_570 : STD_LOGIC;
  SIGNAL and_dcpl_573 : STD_LOGIC;
  SIGNAL and_dcpl_574 : STD_LOGIC;
  SIGNAL and_dcpl_576 : STD_LOGIC;
  SIGNAL and_dcpl_577 : STD_LOGIC;
  SIGNAL and_dcpl_579 : STD_LOGIC;
  SIGNAL and_dcpl_580 : STD_LOGIC;
  SIGNAL and_dcpl_582 : STD_LOGIC;
  SIGNAL and_dcpl_583 : STD_LOGIC;
  SIGNAL and_dcpl_588 : STD_LOGIC;
  SIGNAL and_dcpl_589 : STD_LOGIC;
  SIGNAL and_dcpl_590 : STD_LOGIC;
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_599 : STD_LOGIC;
  SIGNAL and_dcpl_602 : STD_LOGIC;
  SIGNAL and_dcpl_605 : STD_LOGIC;
  SIGNAL and_dcpl_608 : STD_LOGIC;
  SIGNAL and_dcpl_611 : STD_LOGIC;
  SIGNAL and_dcpl_612 : STD_LOGIC;
  SIGNAL and_dcpl_614 : STD_LOGIC;
  SIGNAL and_dcpl_615 : STD_LOGIC;
  SIGNAL and_dcpl_617 : STD_LOGIC;
  SIGNAL and_dcpl_618 : STD_LOGIC;
  SIGNAL and_dcpl_619 : STD_LOGIC;
  SIGNAL and_dcpl_620 : STD_LOGIC;
  SIGNAL and_dcpl_623 : STD_LOGIC;
  SIGNAL and_dcpl_625 : STD_LOGIC;
  SIGNAL z_out_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_dcpl_632 : STD_LOGIC;
  SIGNAL and_dcpl_636 : STD_LOGIC;
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_acc_cse_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tmp_21_sva_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_11 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_13 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_14 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_15 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_17 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_18 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_19 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_21 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_22 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_23 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_25 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_26 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_27 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_29 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_30 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_31 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_33 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_34 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_35 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_37 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_38 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_39 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_41 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_42 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_43 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_45 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_46 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_47 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_49 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_50 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_51 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_53 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_54 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_55 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_57 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_58 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_59 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_61 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_62 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_21_sva_63 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_18_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_20_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_21_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_22_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_23_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_24_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_25_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_26_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_27_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_28_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_29_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_30_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_34_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_36_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_37_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_38_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_39_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_40_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_41_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_42_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_43_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_44_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_45_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_46_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_47_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_48_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_49_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_50_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_51_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_52_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_53_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_54_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_55_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_56_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_57_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_58_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_59_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_60_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_61_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_62_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_73_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_74_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_75_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_100_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_101_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_103_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_104_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_105_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_106_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_107_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_108_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_110_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_115_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_116_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_118_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_120_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_121_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_123_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_124_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_125_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_258_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_260_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_261_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_262_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_264_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_268_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_270_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_272_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_284_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_285_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_286_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_288_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_281_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_282_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_284_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_288_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_296_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_333_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_334_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_335_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_336_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_337_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_338_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_339_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_340_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_341_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_342_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_343_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_344_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_345_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_311_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_347_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_349_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_351_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_352_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_353_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_355_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_356_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_357_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_358_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_359_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_360_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_361_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_363_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_364_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_365_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_366_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_367_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_368_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_369_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_370_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_371_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_372_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_373_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_374_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_375_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_376_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_377_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_509_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_510_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_522_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_505_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_506_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_569_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_508_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_571_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_572_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_573_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_512_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_575_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_576_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_577_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_578_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_579_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_580_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_581_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_520_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_583_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_584_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_585_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_586_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_587_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_588_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_589_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_590_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_591_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_592_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_593_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_594_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_595_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_596_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_597_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_535_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_599_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_600_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_601_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_602_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_603_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_604_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_605_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_606_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_607_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_608_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_609_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_610_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_611_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_612_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_613_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_614_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_615_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_616_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_617_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_618_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_619_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_620_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_621_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_622_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_623_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_624_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_625_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_626_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_627_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_628_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_629_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_760_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_761_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_729_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_730_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_821_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_732_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_823_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_825_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_736_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_827_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_828_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_829_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_830_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_831_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_832_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_833_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_744_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_835_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_836_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_837_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_838_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_839_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_840_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_841_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_842_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_843_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_844_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_845_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_846_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_847_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_848_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_849_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_759_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_852_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_853_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_854_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_855_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_856_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_857_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_859_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_860_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_861_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_862_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_863_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_864_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_865_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_866_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_867_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_868_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_869_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_870_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_871_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_872_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_873_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_874_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_875_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_876_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_877_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_878_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_879_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_880_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_881_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_17_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_953_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_954_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_956_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1077_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_960_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1081_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1083_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1084_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1085_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_968_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1089_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1091_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1092_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1093_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1095_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1096_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1097_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1098_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1099_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1100_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1101_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_983_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1104_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1105_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1107_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1108_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1109_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1110_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1111_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1112_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1113_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1114_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1115_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1116_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1117_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1118_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1119_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1120_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1121_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1122_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1123_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1124_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1125_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1126_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1127_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1128_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1129_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1130_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1131_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1132_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1133_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_141_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_166_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_143_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_168_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_169_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_170_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_146_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_172_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_173_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_175_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_176_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_177_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_178_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_21_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1177_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1178_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1325_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1180_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1327_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1329_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1184_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1333_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1335_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1336_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1337_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1192_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1341_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1343_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1344_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1345_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1346_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1347_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1348_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1349_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1350_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1351_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1352_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1353_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1207_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1357_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1359_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1360_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1361_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1363_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1364_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1365_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1366_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1367_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1368_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1369_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1371_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1372_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1373_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1374_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1375_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1376_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1377_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1378_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1379_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1380_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1381_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1382_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1383_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1384_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1385_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_153_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_157_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_165_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_180_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1518_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_25_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1401_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1402_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1577_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1404_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1579_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1580_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1581_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1408_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1583_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1584_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1585_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1586_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1587_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1588_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1589_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1416_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1591_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1592_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1593_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1594_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1595_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1596_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1597_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1598_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1599_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1600_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1601_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1602_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1603_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1604_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1605_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1431_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1607_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1608_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1609_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1610_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1611_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1612_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1613_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1614_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1615_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1616_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1617_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1618_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1619_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1620_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1621_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1622_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1623_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1624_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1625_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1626_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1627_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1628_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1629_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1630_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1631_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1632_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1633_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1634_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1635_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1636_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1637_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_207_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_209_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_213_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_220_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_29_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1625_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1626_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1829_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1628_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1831_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1832_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1833_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1632_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1835_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1836_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1837_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1838_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1839_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1840_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1841_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1640_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1843_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1844_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1845_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1846_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1847_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1848_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1849_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1850_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1851_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1852_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1853_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1854_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1855_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1856_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1857_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_1655_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1859_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1860_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1861_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1862_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1863_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1864_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1865_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1866_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1867_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1868_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1869_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1870_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1871_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1872_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1873_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1874_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1875_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1876_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1877_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1878_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1879_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1880_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1881_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1882_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1883_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1884_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1885_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1886_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1887_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1888_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1889_itm : STD_LOGIC;
  SIGNAL STAGE_LOOP_i_3_0_sva_mx0c1 : STD_LOGIC;
  SIGNAL VEC_LOOP_j_10_0_sva_9_0_mx0c0 : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_8_itm_mx0c4 : STD_LOGIC;
  SIGNAL COMP_LOOP_1_tmp_mul_idiv_sva_2_0 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL COMP_LOOP_3_tmp_mul_idiv_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_or_120_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_or_110_rgt : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_27_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_28_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_29_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_30_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_31_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_32_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_33_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_76_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_77_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_78_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_79_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_80_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_81_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_82_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_83_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_23_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_140_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_24_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_141_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_25_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_244_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_208_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_63_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_64_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_65_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_67_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_68_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_69_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_70_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_71_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_72_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_61_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_150_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_74_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_151_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_153_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_10_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_18_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_65_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_67_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_68_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_69_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_34_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_35_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_37_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_nor_41_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_92_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_96_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_98_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_99_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse : STD_LOGIC;
  SIGNAL nor_746_cse : STD_LOGIC;
  SIGNAL nor_740_cse : STD_LOGIC;
  SIGNAL nor_735_cse : STD_LOGIC;
  SIGNAL nor_734_cse : STD_LOGIC;
  SIGNAL nor_730_cse : STD_LOGIC;
  SIGNAL nor_719_cse : STD_LOGIC;
  SIGNAL nor_714_cse : STD_LOGIC;
  SIGNAL nor_713_cse : STD_LOGIC;
  SIGNAL nor_709_cse : STD_LOGIC;
  SIGNAL nor_703_cse : STD_LOGIC;
  SIGNAL nor_697_cse : STD_LOGIC;
  SIGNAL nor_692_cse : STD_LOGIC;
  SIGNAL nor_691_cse : STD_LOGIC;
  SIGNAL nor_687_cse : STD_LOGIC;
  SIGNAL nor_676_cse : STD_LOGIC;
  SIGNAL nor_671_cse : STD_LOGIC;
  SIGNAL nor_670_cse : STD_LOGIC;
  SIGNAL nor_666_cse : STD_LOGIC;
  SIGNAL nor_660_cse : STD_LOGIC;
  SIGNAL nor_654_cse : STD_LOGIC;
  SIGNAL nor_649_cse : STD_LOGIC;
  SIGNAL nor_648_cse : STD_LOGIC;
  SIGNAL nor_644_cse : STD_LOGIC;
  SIGNAL nor_633_cse : STD_LOGIC;
  SIGNAL nor_628_cse : STD_LOGIC;
  SIGNAL nor_627_cse : STD_LOGIC;
  SIGNAL nor_623_cse : STD_LOGIC;
  SIGNAL nor_617_cse : STD_LOGIC;
  SIGNAL nor_611_cse : STD_LOGIC;
  SIGNAL nor_606_cse : STD_LOGIC;
  SIGNAL nor_605_cse : STD_LOGIC;
  SIGNAL nor_601_cse : STD_LOGIC;
  SIGNAL nor_590_cse : STD_LOGIC;
  SIGNAL nor_585_cse : STD_LOGIC;
  SIGNAL nor_584_cse : STD_LOGIC;
  SIGNAL and_533_cse : STD_LOGIC;
  SIGNAL nor_576_cse : STD_LOGIC;
  SIGNAL nor_570_cse : STD_LOGIC;
  SIGNAL nor_565_cse : STD_LOGIC;
  SIGNAL nor_564_cse : STD_LOGIC;
  SIGNAL nor_560_cse : STD_LOGIC;
  SIGNAL nor_549_cse : STD_LOGIC;
  SIGNAL nor_544_cse : STD_LOGIC;
  SIGNAL nor_543_cse : STD_LOGIC;
  SIGNAL nor_539_cse : STD_LOGIC;
  SIGNAL nor_533_cse : STD_LOGIC;
  SIGNAL nor_527_cse : STD_LOGIC;
  SIGNAL nor_522_cse : STD_LOGIC;
  SIGNAL nor_521_cse : STD_LOGIC;
  SIGNAL nor_517_cse : STD_LOGIC;
  SIGNAL nor_506_cse : STD_LOGIC;
  SIGNAL nor_501_cse : STD_LOGIC;
  SIGNAL nor_500_cse : STD_LOGIC;
  SIGNAL and_531_cse : STD_LOGIC;
  SIGNAL nor_492_cse : STD_LOGIC;
  SIGNAL nor_486_cse : STD_LOGIC;
  SIGNAL nor_481_cse : STD_LOGIC;
  SIGNAL nor_480_cse : STD_LOGIC;
  SIGNAL nor_476_cse : STD_LOGIC;
  SIGNAL nor_465_cse : STD_LOGIC;
  SIGNAL nor_460_cse : STD_LOGIC;
  SIGNAL nor_459_cse : STD_LOGIC;
  SIGNAL and_529_cse : STD_LOGIC;
  SIGNAL nor_451_cse : STD_LOGIC;
  SIGNAL nor_446_cse : STD_LOGIC;
  SIGNAL nor_441_cse : STD_LOGIC;
  SIGNAL nor_440_cse : STD_LOGIC;
  SIGNAL and_526_cse : STD_LOGIC;
  SIGNAL and_523_cse : STD_LOGIC;
  SIGNAL and_519_cse : STD_LOGIC;
  SIGNAL and_518_cse : STD_LOGIC;
  SIGNAL and_515_cse : STD_LOGIC;
  SIGNAL nor_1716_cse : STD_LOGIC;
  SIGNAL nor_1715_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_121_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_126_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_135_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_151_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_153_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_49_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_50_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_52_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_56_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_57_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_58_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_59_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_60_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_62_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_63_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_64_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_66_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_74_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_75_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_76_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_78_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_79_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_87_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_88_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_89_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_90_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_91_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_93_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_94_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_95_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_97_cse : STD_LOGIC;
  SIGNAL and_907_cse : STD_LOGIC;
  SIGNAL and_918_cse : STD_LOGIC;
  SIGNAL and_903_cse : STD_LOGIC;
  SIGNAL and_910_cse : STD_LOGIC;
  SIGNAL and_914_cse : STD_LOGIC;
  SIGNAL and_920_cse : STD_LOGIC;
  SIGNAL nor_1744_cse : STD_LOGIC;
  SIGNAL and_1046_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_or_68_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_or_65_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_83_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_2_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_3_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_4_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_5_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_6_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_7_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_8_acc_10_itm_10_1_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_or_54_ssc : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_724_cse : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_nor_300_cse : STD_LOGIC;

  SIGNAL nor_1423_nl : STD_LOGIC;
  SIGNAL mux_789_nl : STD_LOGIC;
  SIGNAL mux_788_nl : STD_LOGIC;
  SIGNAL mux_2996_nl : STD_LOGIC;
  SIGNAL mux_2995_nl : STD_LOGIC;
  SIGNAL mux_2993_nl : STD_LOGIC;
  SIGNAL mux_2992_nl : STD_LOGIC;
  SIGNAL nor_425_nl : STD_LOGIC;
  SIGNAL VEC_LOOP_j_not_1_nl : STD_LOGIC;
  SIGNAL nor_422_nl : STD_LOGIC;
  SIGNAL nand_480_nl : STD_LOGIC;
  SIGNAL mux_781_nl : STD_LOGIC;
  SIGNAL nor_1426_nl : STD_LOGIC;
  SIGNAL and_637_nl : STD_LOGIC;
  SIGNAL or_4159_nl : STD_LOGIC;
  SIGNAL nand_493_nl : STD_LOGIC;
  SIGNAL mux_3365_nl : STD_LOGIC;
  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL nor_1745_nl : STD_LOGIC;
  SIGNAL or_4154_nl : STD_LOGIC;
  SIGNAL mux_3031_nl : STD_LOGIC;
  SIGNAL mux_3030_nl : STD_LOGIC;
  SIGNAL mux_3029_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_73_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_824_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_74_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_851_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_75_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_858_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_100_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_323_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1073_nl : STD_LOGIC;
  SIGNAL mux_3037_nl : STD_LOGIC;
  SIGNAL mux_3036_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_101_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_348_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1075_nl : STD_LOGIC;
  SIGNAL and_403_nl : STD_LOGIC;
  SIGNAL mux_3039_nl : STD_LOGIC;
  SIGNAL nor_420_nl : STD_LOGIC;
  SIGNAL mux_3045_nl : STD_LOGIC;
  SIGNAL mux_3044_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_102_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1076_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_103_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_350_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1079_nl : STD_LOGIC;
  SIGNAL mux_3046_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_104_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_354_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1080_nl : STD_LOGIC;
  SIGNAL and_409_nl : STD_LOGIC;
  SIGNAL mux_3047_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_105_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_362_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1082_nl : STD_LOGIC;
  SIGNAL mux_3048_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_106_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1087_nl : STD_LOGIC;
  SIGNAL and_411_nl : STD_LOGIC;
  SIGNAL mux_3053_nl : STD_LOGIC;
  SIGNAL mux_3052_nl : STD_LOGIC;
  SIGNAL mux_3051_nl : STD_LOGIC;
  SIGNAL or_3878_nl : STD_LOGIC;
  SIGNAL or_3877_nl : STD_LOGIC;
  SIGNAL mux_3050_nl : STD_LOGIC;
  SIGNAL mux_3049_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL or_3874_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_107_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1088_nl : STD_LOGIC;
  SIGNAL mux_3059_nl : STD_LOGIC;
  SIGNAL mux_3056_nl : STD_LOGIC;
  SIGNAL mux_3055_nl : STD_LOGIC;
  SIGNAL mux_3054_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_108_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1090_nl : STD_LOGIC;
  SIGNAL mux_3063_nl : STD_LOGIC;
  SIGNAL mux_3062_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_109_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1094_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_110_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1103_nl : STD_LOGIC;
  SIGNAL mux_3064_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_115_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1328_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_116_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1331_nl : STD_LOGIC;
  SIGNAL mux_3073_nl : STD_LOGIC;
  SIGNAL or_3889_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_117_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1332_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_118_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1334_nl : STD_LOGIC;
  SIGNAL mux_3081_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_119_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1339_nl : STD_LOGIC;
  SIGNAL mux_3085_nl : STD_LOGIC;
  SIGNAL mux_3084_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_120_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1340_nl : STD_LOGIC;
  SIGNAL mux_3092_nl : STD_LOGIC;
  SIGNAL mux_3091_nl : STD_LOGIC;
  SIGNAL mux_3090_nl : STD_LOGIC;
  SIGNAL mux_3089_nl : STD_LOGIC;
  SIGNAL mux_3087_nl : STD_LOGIC;
  SIGNAL mux_3094_nl : STD_LOGIC;
  SIGNAL or_3900_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_121_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1342_nl : STD_LOGIC;
  SIGNAL mux_3097_nl : STD_LOGIC;
  SIGNAL mux_3096_nl : STD_LOGIC;
  SIGNAL and_503_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_122_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1355_nl : STD_LOGIC;
  SIGNAL or_560_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_123_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1356_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_124_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1358_nl : STD_LOGIC;
  SIGNAL mux_3102_nl : STD_LOGIC;
  SIGNAL or_3904_nl : STD_LOGIC;
  SIGNAL nand_145_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_125_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1362_nl : STD_LOGIC;
  SIGNAL mux_3107_nl : STD_LOGIC;
  SIGNAL mux_3106_nl : STD_LOGIC;
  SIGNAL mux_3105_nl : STD_LOGIC;
  SIGNAL mux_3104_nl : STD_LOGIC;
  SIGNAL mux_3111_nl : STD_LOGIC;
  SIGNAL mux_3110_nl : STD_LOGIC;
  SIGNAL mux_3115_nl : STD_LOGIC;
  SIGNAL mux_3113_nl : STD_LOGIC;
  SIGNAL mux_3123_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_3_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_3124_nl : STD_LOGIC;
  SIGNAL nand_149_nl : STD_LOGIC;
  SIGNAL mux_3126_nl : STD_LOGIC;
  SIGNAL mux_3125_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_12_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL mux_3128_nl : STD_LOGIC;
  SIGNAL mux_3127_nl : STD_LOGIC;
  SIGNAL mux_3130_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_5_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_3132_nl : STD_LOGIC;
  SIGNAL mux_3131_nl : STD_LOGIC;
  SIGNAL mux_3140_nl : STD_LOGIC;
  SIGNAL mux_3139_nl : STD_LOGIC;
  SIGNAL mux_3138_nl : STD_LOGIC;
  SIGNAL and_497_nl : STD_LOGIC;
  SIGNAL mux_3143_nl : STD_LOGIC;
  SIGNAL mux_3142_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_6_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_3146_nl : STD_LOGIC;
  SIGNAL mux_3152_nl : STD_LOGIC;
  SIGNAL mux_212_nl : STD_LOGIC;
  SIGNAL mux_3160_nl : STD_LOGIC;
  SIGNAL mux_219_nl : STD_LOGIC;
  SIGNAL or_154_nl : STD_LOGIC;
  SIGNAL mux_3163_nl : STD_LOGIC;
  SIGNAL mux_3162_nl : STD_LOGIC;
  SIGNAL mux_3161_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL and_491_nl : STD_LOGIC;
  SIGNAL and_492_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_7_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_3171_nl : STD_LOGIC;
  SIGNAL mux_3182_nl : STD_LOGIC;
  SIGNAL mux_3181_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_15_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL mux_3188_nl : STD_LOGIC;
  SIGNAL nand_148_nl : STD_LOGIC;
  SIGNAL mux_3192_nl : STD_LOGIC;
  SIGNAL mux_361_nl : STD_LOGIC;
  SIGNAL mux_359_nl : STD_LOGIC;
  SIGNAL mux_3193_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_3197_nl : STD_LOGIC;
  SIGNAL mux_3205_nl : STD_LOGIC;
  SIGNAL mux_3204_nl : STD_LOGIC;
  SIGNAL mux_3203_nl : STD_LOGIC;
  SIGNAL and_489_nl : STD_LOGIC;
  SIGNAL mux_3202_nl : STD_LOGIC;
  SIGNAL mux_3210_nl : STD_LOGIC;
  SIGNAL mux_3209_nl : STD_LOGIC;
  SIGNAL mux_3208_nl : STD_LOGIC;
  SIGNAL and_449_nl : STD_LOGIC;
  SIGNAL mux_3207_nl : STD_LOGIC;
  SIGNAL mux_3206_nl : STD_LOGIC;
  SIGNAL mux_3216_nl : STD_LOGIC;
  SIGNAL mux_3215_nl : STD_LOGIC;
  SIGNAL mux_3214_nl : STD_LOGIC;
  SIGNAL mux_3213_nl : STD_LOGIC;
  SIGNAL mux_3212_nl : STD_LOGIC;
  SIGNAL mux_3211_nl : STD_LOGIC;
  SIGNAL mux_3219_nl : STD_LOGIC;
  SIGNAL mux_435_nl : STD_LOGIC;
  SIGNAL mux_434_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_111_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1104_nl : STD_LOGIC;
  SIGNAL mux_3223_nl : STD_LOGIC;
  SIGNAL mux_3222_nl : STD_LOGIC;
  SIGNAL mux_3221_nl : STD_LOGIC;
  SIGNAL or_3932_nl : STD_LOGIC;
  SIGNAL mux_3220_nl : STD_LOGIC;
  SIGNAL or_3929_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_112_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1106_nl : STD_LOGIC;
  SIGNAL mux_3226_nl : STD_LOGIC;
  SIGNAL mux_3225_nl : STD_LOGIC;
  SIGNAL mux_3224_nl : STD_LOGIC;
  SIGNAL or_3934_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_113_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1110_nl : STD_LOGIC;
  SIGNAL mux_3227_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_114_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1118_nl : STD_LOGIC;
  SIGNAL mux_3229_nl : STD_LOGIC;
  SIGNAL mux_3228_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_65_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1370_nl : STD_LOGIC;
  SIGNAL mux_3231_nl : STD_LOGIC;
  SIGNAL mux_3230_nl : STD_LOGIC;
  SIGNAL mux_3234_nl : STD_LOGIC;
  SIGNAL mux_3233_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_67_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1577_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_68_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1584_nl : STD_LOGIC;
  SIGNAL mux_3238_nl : STD_LOGIC;
  SIGNAL mux_3237_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_317_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1594_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_319_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1598_nl : STD_LOGIC;
  SIGNAL mux_3243_nl : STD_LOGIC;
  SIGNAL mux_3242_nl : STD_LOGIC;
  SIGNAL mux_3241_nl : STD_LOGIC;
  SIGNAL nor_403_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL mux_3240_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_320_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1607_nl : STD_LOGIC;
  SIGNAL and_458_nl : STD_LOGIC;
  SIGNAL mux_3246_nl : STD_LOGIC;
  SIGNAL mux_3245_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_321_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1610_nl : STD_LOGIC;
  SIGNAL mux_3253_nl : STD_LOGIC;
  SIGNAL mux_3252_nl : STD_LOGIC;
  SIGNAL mux_3251_nl : STD_LOGIC;
  SIGNAL or_3946_nl : STD_LOGIC;
  SIGNAL mux_582_nl : STD_LOGIC;
  SIGNAL mux_3249_nl : STD_LOGIC;
  SIGNAL mux_3248_nl : STD_LOGIC;
  SIGNAL or_3943_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_324_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1614_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_325_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1622_nl : STD_LOGIC;
  SIGNAL and_459_nl : STD_LOGIC;
  SIGNAL mux_3256_nl : STD_LOGIC;
  SIGNAL mux_3255_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_69_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1831_nl : STD_LOGIC;
  SIGNAL mux_3264_nl : STD_LOGIC;
  SIGNAL mux_3261_nl : STD_LOGIC;
  SIGNAL mux_3259_nl : STD_LOGIC;
  SIGNAL mux_3258_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_326_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1832_nl : STD_LOGIC;
  SIGNAL and_461_nl : STD_LOGIC;
  SIGNAL mux_3274_nl : STD_LOGIC;
  SIGNAL mux_3273_nl : STD_LOGIC;
  SIGNAL mux_3272_nl : STD_LOGIC;
  SIGNAL mux_3271_nl : STD_LOGIC;
  SIGNAL mux_3270_nl : STD_LOGIC;
  SIGNAL mux_3269_nl : STD_LOGIC;
  SIGNAL mux_3268_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL mux_3267_nl : STD_LOGIC;
  SIGNAL nor_384_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_327_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1835_nl : STD_LOGIC;
  SIGNAL and_463_nl : STD_LOGIC;
  SIGNAL mux_3283_nl : STD_LOGIC;
  SIGNAL mux_3282_nl : STD_LOGIC;
  SIGNAL mux_3279_nl : STD_LOGIC;
  SIGNAL mux_3278_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_328_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1844_nl : STD_LOGIC;
  SIGNAL mux_3286_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_329_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1850_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_331_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1862_nl : STD_LOGIC;
  SIGNAL and_465_nl : STD_LOGIC;
  SIGNAL mux_3292_nl : STD_LOGIC;
  SIGNAL mux_3291_nl : STD_LOGIC;
  SIGNAL and_464_nl : STD_LOGIC;
  SIGNAL mux_3290_nl : STD_LOGIC;
  SIGNAL mux_3289_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_332_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1866_nl : STD_LOGIC;
  SIGNAL and_468_nl : STD_LOGIC;
  SIGNAL mux_3298_nl : STD_LOGIC;
  SIGNAL mux_3297_nl : STD_LOGIC;
  SIGNAL mux_3296_nl : STD_LOGIC;
  SIGNAL and_73_nl : STD_LOGIC;
  SIGNAL mux_3295_nl : STD_LOGIC;
  SIGNAL mux_3294_nl : STD_LOGIC;
  SIGNAL and_466_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_71_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1874_nl : STD_LOGIC;
  SIGNAL mux_3302_nl : STD_LOGIC;
  SIGNAL mux_3301_nl : STD_LOGIC;
  SIGNAL mux_3300_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_72_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_583_nl : STD_LOGIC;
  SIGNAL mux_3306_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_nor_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_76_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_77_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_79_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_80_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_81_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_82_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_83_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_84_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_85_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_86_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_87_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_88_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_89_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_90_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_91_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_92_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_93_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_95_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_96_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_97_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_98_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_99_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_57_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_58_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_60_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_64_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_72_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_87_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_17_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_mux_21_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_or_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_23_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_24_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_25_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_28_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_30_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_31_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_32_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_33_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_34_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_35_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_36_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_37_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_38_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_39_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_40_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_41_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_42_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_43_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_44_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_45_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_46_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_47_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_48_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_49_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_50_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_51_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_52_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_53_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_54_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_55_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_56_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_57_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_58_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_59_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_60_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_61_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_62_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_63_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_249_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_250_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_251_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_252_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_253_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_254_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_255_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_256_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_257_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_258_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_259_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_260_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_261_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_262_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_263_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_264_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_265_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_266_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_267_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_268_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_269_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_270_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_271_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_272_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_273_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_274_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_275_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_276_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_277_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_278_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_279_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_280_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_281_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_282_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_283_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_284_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_285_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_286_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_287_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_288_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_289_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_290_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_291_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_292_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_293_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_294_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_295_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_296_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_297_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_298_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_299_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_300_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_301_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_302_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_303_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_304_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_305_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_306_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_222_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_70_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_71_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_223_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_73_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_224_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_225_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_226_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_77_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_227_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_228_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_229_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_230_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_231_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_232_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_233_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_234_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_235_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_236_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_237_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_238_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_239_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_240_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_241_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_242_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_243_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_244_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_245_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_246_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_247_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_248_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_164_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_102_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_165_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_166_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_167_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_168_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_169_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_170_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_171_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_172_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_173_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_174_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_175_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_176_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_177_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_178_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_179_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_180_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_181_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_182_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_183_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_184_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_185_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_186_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_187_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_188_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_189_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_190_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_191_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_192_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_193_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_194_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_195_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_196_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_197_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_198_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_199_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_200_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_201_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_202_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_203_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_204_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_205_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_206_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_207_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_208_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_209_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_210_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_211_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_212_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_213_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_214_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_215_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_216_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_217_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_218_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_219_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_220_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_221_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_152_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_164_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_165_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_153_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_167_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_154_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_155_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_156_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_171_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_157_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_158_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_159_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_160_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_161_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_162_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_163_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_89_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_90_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_91_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_92_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_93_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_94_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_95_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_96_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_97_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_98_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_99_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_100_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_101_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_102_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_103_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_104_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_105_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_106_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_107_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_108_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_109_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_110_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_111_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_112_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_113_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_114_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_115_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_116_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_117_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_118_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_119_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_120_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_121_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_122_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_123_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_124_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_125_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_126_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_127_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_128_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_129_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_130_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_131_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_132_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_133_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_134_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_135_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_136_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_137_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_138_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_139_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_140_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_141_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_142_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_143_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_144_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_145_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_146_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_147_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_148_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_149_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_150_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_151_nl : STD_LOGIC;
  SIGNAL mux_3353_nl : STD_LOGIC;
  SIGNAL mux_3352_nl : STD_LOGIC;
  SIGNAL mux_3351_nl : STD_LOGIC;
  SIGNAL mux_3350_nl : STD_LOGIC;
  SIGNAL mux_3349_nl : STD_LOGIC;
  SIGNAL mux_3348_nl : STD_LOGIC;
  SIGNAL mux_3359_nl : STD_LOGIC;
  SIGNAL mux_3358_nl : STD_LOGIC;
  SIGNAL mux_3357_nl : STD_LOGIC;
  SIGNAL mux_3356_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_31_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_179_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_180_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_32_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_182_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_33_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_34_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_35_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_186_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_36_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_37_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_38_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_39_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_40_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_41_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_42_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_194_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_43_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_44_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_45_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_46_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_47_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_48_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_49_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_50_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_51_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_52_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_53_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_54_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_55_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_56_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_57_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_210_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_58_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_59_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_60_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_61_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_62_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_63_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_64_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_65_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_66_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_67_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_68_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_69_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_70_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_71_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_72_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_73_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_74_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_75_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_76_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_77_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_78_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_79_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_80_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_81_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_82_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_83_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_84_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_85_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_86_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_87_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_88_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_2_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_5_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_22_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_23_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_24_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_25_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_26_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_27_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_28_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_29_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_30_nl : STD_LOGIC;
  SIGNAL mux_3364_nl : STD_LOGIC;
  SIGNAL mux_3363_nl : STD_LOGIC;
  SIGNAL mux_3362_nl : STD_LOGIC;
  SIGNAL mux_3361_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_2_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_3_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_4_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_5_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_6_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_7_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_8_acc_10_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL mux_510_nl : STD_LOGIC;
  SIGNAL or_201_nl : STD_LOGIC;
  SIGNAL mux_3004_nl : STD_LOGIC;
  SIGNAL mux_522_nl : STD_LOGIC;
  SIGNAL or_3843_nl : STD_LOGIC;
  SIGNAL mux_3024_nl : STD_LOGIC;
  SIGNAL mux_3021_nl : STD_LOGIC;
  SIGNAL mux_3034_nl : STD_LOGIC;
  SIGNAL mux_3041_nl : STD_LOGIC;
  SIGNAL mux_3057_nl : STD_LOGIC;
  SIGNAL or_3880_nl : STD_LOGIC;
  SIGNAL or_3887_nl : STD_LOGIC;
  SIGNAL mux_3069_nl : STD_LOGIC;
  SIGNAL mux_3067_nl : STD_LOGIC;
  SIGNAL mux_3065_nl : STD_LOGIC;
  SIGNAL or_3884_nl : STD_LOGIC;
  SIGNAL mux_3075_nl : STD_LOGIC;
  SIGNAL or_3906_nl : STD_LOGIC;
  SIGNAL mux_3119_nl : STD_LOGIC;
  SIGNAL mux_3118_nl : STD_LOGIC;
  SIGNAL mux_3117_nl : STD_LOGIC;
  SIGNAL mux_3122_nl : STD_LOGIC;
  SIGNAL mux_67_nl : STD_LOGIC;
  SIGNAL mux_3129_nl : STD_LOGIC;
  SIGNAL mux_3135_nl : STD_LOGIC;
  SIGNAL mux_3134_nl : STD_LOGIC;
  SIGNAL mux_3133_nl : STD_LOGIC;
  SIGNAL nor_1425_nl : STD_LOGIC;
  SIGNAL mux_3148_nl : STD_LOGIC;
  SIGNAL mux_3150_nl : STD_LOGIC;
  SIGNAL mux_210_nl : STD_LOGIC;
  SIGNAL mux_3156_nl : STD_LOGIC;
  SIGNAL mux_215_nl : STD_LOGIC;
  SIGNAL mux_214_nl : STD_LOGIC;
  SIGNAL mux_3158_nl : STD_LOGIC;
  SIGNAL mux_217_nl : STD_LOGIC;
  SIGNAL mux_3166_nl : STD_LOGIC;
  SIGNAL mux_3174_nl : STD_LOGIC;
  SIGNAL mux_3173_nl : STD_LOGIC;
  SIGNAL mux_3178_nl : STD_LOGIC;
  SIGNAL mux_3177_nl : STD_LOGIC;
  SIGNAL mux_3176_nl : STD_LOGIC;
  SIGNAL mux_3180_nl : STD_LOGIC;
  SIGNAL mux_3179_nl : STD_LOGIC;
  SIGNAL mux_3184_nl : STD_LOGIC;
  SIGNAL nor_1524_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL mux_3199_nl : STD_LOGIC;
  SIGNAL mux_3262_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL nor_1474_nl : STD_LOGIC;
  SIGNAL mux_75_nl : STD_LOGIC;
  SIGNAL mux_3314_nl : STD_LOGIC;
  SIGNAL nor_1709_nl : STD_LOGIC;
  SIGNAL nor_1710_nl : STD_LOGIC;
  SIGNAL mux_3354_nl : STD_LOGIC;
  SIGNAL mux_3320_nl : STD_LOGIC;
  SIGNAL mux_3319_nl : STD_LOGIC;
  SIGNAL mux_3318_nl : STD_LOGIC;
  SIGNAL mux_3317_nl : STD_LOGIC;
  SIGNAL mux_3316_nl : STD_LOGIC;
  SIGNAL or_3973_nl : STD_LOGIC;
  SIGNAL mux_3315_nl : STD_LOGIC;
  SIGNAL mux_3340_nl : STD_LOGIC;
  SIGNAL mux_3343_nl : STD_LOGIC;
  SIGNAL mux_3342_nl : STD_LOGIC;
  SIGNAL mux_104_nl : STD_LOGIC;
  SIGNAL mux_3346_nl : STD_LOGIC;
  SIGNAL mux_3345_nl : STD_LOGIC;
  SIGNAL mux_3344_nl : STD_LOGIC;
  SIGNAL and_102_nl : STD_LOGIC;
  SIGNAL and_114_nl : STD_LOGIC;
  SIGNAL and_120_nl : STD_LOGIC;
  SIGNAL and_124_nl : STD_LOGIC;
  SIGNAL and_129_nl : STD_LOGIC;
  SIGNAL and_133_nl : STD_LOGIC;
  SIGNAL and_136_nl : STD_LOGIC;
  SIGNAL and_138_nl : STD_LOGIC;
  SIGNAL and_142_nl : STD_LOGIC;
  SIGNAL and_145_nl : STD_LOGIC;
  SIGNAL and_148_nl : STD_LOGIC;
  SIGNAL and_151_nl : STD_LOGIC;
  SIGNAL and_152_nl : STD_LOGIC;
  SIGNAL and_153_nl : STD_LOGIC;
  SIGNAL and_154_nl : STD_LOGIC;
  SIGNAL and_155_nl : STD_LOGIC;
  SIGNAL and_156_nl : STD_LOGIC;
  SIGNAL and_157_nl : STD_LOGIC;
  SIGNAL and_158_nl : STD_LOGIC;
  SIGNAL and_159_nl : STD_LOGIC;
  SIGNAL and_160_nl : STD_LOGIC;
  SIGNAL mux_805_nl : STD_LOGIC;
  SIGNAL nand_469_nl : STD_LOGIC;
  SIGNAL mux_804_nl : STD_LOGIC;
  SIGNAL mux_803_nl : STD_LOGIC;
  SIGNAL mux_802_nl : STD_LOGIC;
  SIGNAL nor_1414_nl : STD_LOGIC;
  SIGNAL nor_1415_nl : STD_LOGIC;
  SIGNAL mux_801_nl : STD_LOGIC;
  SIGNAL nor_1416_nl : STD_LOGIC;
  SIGNAL nor_1417_nl : STD_LOGIC;
  SIGNAL mux_800_nl : STD_LOGIC;
  SIGNAL mux_799_nl : STD_LOGIC;
  SIGNAL nor_1418_nl : STD_LOGIC;
  SIGNAL nor_1419_nl : STD_LOGIC;
  SIGNAL mux_798_nl : STD_LOGIC;
  SIGNAL nor_1420_nl : STD_LOGIC;
  SIGNAL nor_1421_nl : STD_LOGIC;
  SIGNAL or_4142_nl : STD_LOGIC;
  SIGNAL mux_797_nl : STD_LOGIC;
  SIGNAL mux_796_nl : STD_LOGIC;
  SIGNAL mux_795_nl : STD_LOGIC;
  SIGNAL or_615_nl : STD_LOGIC;
  SIGNAL mux_794_nl : STD_LOGIC;
  SIGNAL or_612_nl : STD_LOGIC;
  SIGNAL mux_793_nl : STD_LOGIC;
  SIGNAL mux_792_nl : STD_LOGIC;
  SIGNAL or_609_nl : STD_LOGIC;
  SIGNAL mux_791_nl : STD_LOGIC;
  SIGNAL or_606_nl : STD_LOGIC;
  SIGNAL mux_820_nl : STD_LOGIC;
  SIGNAL mux_819_nl : STD_LOGIC;
  SIGNAL or_649_nl : STD_LOGIC;
  SIGNAL mux_818_nl : STD_LOGIC;
  SIGNAL or_648_nl : STD_LOGIC;
  SIGNAL or_647_nl : STD_LOGIC;
  SIGNAL mux_817_nl : STD_LOGIC;
  SIGNAL mux_816_nl : STD_LOGIC;
  SIGNAL mux_815_nl : STD_LOGIC;
  SIGNAL or_645_nl : STD_LOGIC;
  SIGNAL mux_814_nl : STD_LOGIC;
  SIGNAL or_643_nl : STD_LOGIC;
  SIGNAL mux_813_nl : STD_LOGIC;
  SIGNAL mux_812_nl : STD_LOGIC;
  SIGNAL or_642_nl : STD_LOGIC;
  SIGNAL mux_811_nl : STD_LOGIC;
  SIGNAL or_640_nl : STD_LOGIC;
  SIGNAL or_639_nl : STD_LOGIC;
  SIGNAL mux_810_nl : STD_LOGIC;
  SIGNAL mux_809_nl : STD_LOGIC;
  SIGNAL mux_808_nl : STD_LOGIC;
  SIGNAL or_638_nl : STD_LOGIC;
  SIGNAL or_636_nl : STD_LOGIC;
  SIGNAL mux_807_nl : STD_LOGIC;
  SIGNAL or_634_nl : STD_LOGIC;
  SIGNAL or_633_nl : STD_LOGIC;
  SIGNAL nand_15_nl : STD_LOGIC;
  SIGNAL mux_806_nl : STD_LOGIC;
  SIGNAL nor_1412_nl : STD_LOGIC;
  SIGNAL nor_1413_nl : STD_LOGIC;
  SIGNAL mux_835_nl : STD_LOGIC;
  SIGNAL nand_468_nl : STD_LOGIC;
  SIGNAL mux_834_nl : STD_LOGIC;
  SIGNAL mux_833_nl : STD_LOGIC;
  SIGNAL mux_832_nl : STD_LOGIC;
  SIGNAL nor_1403_nl : STD_LOGIC;
  SIGNAL nor_1404_nl : STD_LOGIC;
  SIGNAL mux_831_nl : STD_LOGIC;
  SIGNAL nor_1405_nl : STD_LOGIC;
  SIGNAL nor_1406_nl : STD_LOGIC;
  SIGNAL mux_830_nl : STD_LOGIC;
  SIGNAL mux_829_nl : STD_LOGIC;
  SIGNAL nor_1407_nl : STD_LOGIC;
  SIGNAL nor_1408_nl : STD_LOGIC;
  SIGNAL mux_828_nl : STD_LOGIC;
  SIGNAL nor_1409_nl : STD_LOGIC;
  SIGNAL nor_1410_nl : STD_LOGIC;
  SIGNAL or_4141_nl : STD_LOGIC;
  SIGNAL mux_827_nl : STD_LOGIC;
  SIGNAL mux_826_nl : STD_LOGIC;
  SIGNAL mux_825_nl : STD_LOGIC;
  SIGNAL or_659_nl : STD_LOGIC;
  SIGNAL mux_824_nl : STD_LOGIC;
  SIGNAL or_656_nl : STD_LOGIC;
  SIGNAL mux_823_nl : STD_LOGIC;
  SIGNAL mux_822_nl : STD_LOGIC;
  SIGNAL or_653_nl : STD_LOGIC;
  SIGNAL mux_821_nl : STD_LOGIC;
  SIGNAL or_650_nl : STD_LOGIC;
  SIGNAL mux_850_nl : STD_LOGIC;
  SIGNAL mux_849_nl : STD_LOGIC;
  SIGNAL or_693_nl : STD_LOGIC;
  SIGNAL mux_848_nl : STD_LOGIC;
  SIGNAL or_692_nl : STD_LOGIC;
  SIGNAL or_691_nl : STD_LOGIC;
  SIGNAL mux_847_nl : STD_LOGIC;
  SIGNAL mux_846_nl : STD_LOGIC;
  SIGNAL mux_845_nl : STD_LOGIC;
  SIGNAL or_689_nl : STD_LOGIC;
  SIGNAL mux_844_nl : STD_LOGIC;
  SIGNAL or_687_nl : STD_LOGIC;
  SIGNAL mux_843_nl : STD_LOGIC;
  SIGNAL mux_842_nl : STD_LOGIC;
  SIGNAL or_686_nl : STD_LOGIC;
  SIGNAL mux_841_nl : STD_LOGIC;
  SIGNAL or_684_nl : STD_LOGIC;
  SIGNAL or_683_nl : STD_LOGIC;
  SIGNAL mux_840_nl : STD_LOGIC;
  SIGNAL mux_839_nl : STD_LOGIC;
  SIGNAL mux_838_nl : STD_LOGIC;
  SIGNAL or_682_nl : STD_LOGIC;
  SIGNAL or_680_nl : STD_LOGIC;
  SIGNAL mux_837_nl : STD_LOGIC;
  SIGNAL or_678_nl : STD_LOGIC;
  SIGNAL or_677_nl : STD_LOGIC;
  SIGNAL nand_17_nl : STD_LOGIC;
  SIGNAL mux_836_nl : STD_LOGIC;
  SIGNAL nor_1401_nl : STD_LOGIC;
  SIGNAL nor_1402_nl : STD_LOGIC;
  SIGNAL mux_865_nl : STD_LOGIC;
  SIGNAL nand_467_nl : STD_LOGIC;
  SIGNAL mux_864_nl : STD_LOGIC;
  SIGNAL mux_863_nl : STD_LOGIC;
  SIGNAL mux_862_nl : STD_LOGIC;
  SIGNAL nor_1392_nl : STD_LOGIC;
  SIGNAL nor_1393_nl : STD_LOGIC;
  SIGNAL mux_861_nl : STD_LOGIC;
  SIGNAL nor_1394_nl : STD_LOGIC;
  SIGNAL nor_1395_nl : STD_LOGIC;
  SIGNAL mux_860_nl : STD_LOGIC;
  SIGNAL mux_859_nl : STD_LOGIC;
  SIGNAL nor_1396_nl : STD_LOGIC;
  SIGNAL nor_1397_nl : STD_LOGIC;
  SIGNAL mux_858_nl : STD_LOGIC;
  SIGNAL nor_1398_nl : STD_LOGIC;
  SIGNAL nor_1399_nl : STD_LOGIC;
  SIGNAL or_4140_nl : STD_LOGIC;
  SIGNAL mux_857_nl : STD_LOGIC;
  SIGNAL mux_856_nl : STD_LOGIC;
  SIGNAL mux_855_nl : STD_LOGIC;
  SIGNAL or_703_nl : STD_LOGIC;
  SIGNAL mux_854_nl : STD_LOGIC;
  SIGNAL or_700_nl : STD_LOGIC;
  SIGNAL mux_853_nl : STD_LOGIC;
  SIGNAL mux_852_nl : STD_LOGIC;
  SIGNAL or_697_nl : STD_LOGIC;
  SIGNAL mux_851_nl : STD_LOGIC;
  SIGNAL or_694_nl : STD_LOGIC;
  SIGNAL mux_880_nl : STD_LOGIC;
  SIGNAL mux_879_nl : STD_LOGIC;
  SIGNAL or_737_nl : STD_LOGIC;
  SIGNAL mux_878_nl : STD_LOGIC;
  SIGNAL or_736_nl : STD_LOGIC;
  SIGNAL or_735_nl : STD_LOGIC;
  SIGNAL mux_877_nl : STD_LOGIC;
  SIGNAL mux_876_nl : STD_LOGIC;
  SIGNAL mux_875_nl : STD_LOGIC;
  SIGNAL or_733_nl : STD_LOGIC;
  SIGNAL mux_874_nl : STD_LOGIC;
  SIGNAL or_731_nl : STD_LOGIC;
  SIGNAL mux_873_nl : STD_LOGIC;
  SIGNAL mux_872_nl : STD_LOGIC;
  SIGNAL or_730_nl : STD_LOGIC;
  SIGNAL mux_871_nl : STD_LOGIC;
  SIGNAL or_728_nl : STD_LOGIC;
  SIGNAL or_727_nl : STD_LOGIC;
  SIGNAL mux_870_nl : STD_LOGIC;
  SIGNAL mux_869_nl : STD_LOGIC;
  SIGNAL mux_868_nl : STD_LOGIC;
  SIGNAL or_726_nl : STD_LOGIC;
  SIGNAL or_724_nl : STD_LOGIC;
  SIGNAL mux_867_nl : STD_LOGIC;
  SIGNAL or_722_nl : STD_LOGIC;
  SIGNAL or_721_nl : STD_LOGIC;
  SIGNAL nand_19_nl : STD_LOGIC;
  SIGNAL mux_866_nl : STD_LOGIC;
  SIGNAL nor_1390_nl : STD_LOGIC;
  SIGNAL nor_1391_nl : STD_LOGIC;
  SIGNAL mux_895_nl : STD_LOGIC;
  SIGNAL nand_466_nl : STD_LOGIC;
  SIGNAL mux_894_nl : STD_LOGIC;
  SIGNAL mux_893_nl : STD_LOGIC;
  SIGNAL mux_892_nl : STD_LOGIC;
  SIGNAL nor_1381_nl : STD_LOGIC;
  SIGNAL nor_1382_nl : STD_LOGIC;
  SIGNAL mux_891_nl : STD_LOGIC;
  SIGNAL nor_1383_nl : STD_LOGIC;
  SIGNAL nor_1384_nl : STD_LOGIC;
  SIGNAL mux_890_nl : STD_LOGIC;
  SIGNAL mux_889_nl : STD_LOGIC;
  SIGNAL nor_1385_nl : STD_LOGIC;
  SIGNAL nor_1386_nl : STD_LOGIC;
  SIGNAL mux_888_nl : STD_LOGIC;
  SIGNAL nor_1387_nl : STD_LOGIC;
  SIGNAL nor_1388_nl : STD_LOGIC;
  SIGNAL or_4139_nl : STD_LOGIC;
  SIGNAL mux_887_nl : STD_LOGIC;
  SIGNAL mux_886_nl : STD_LOGIC;
  SIGNAL mux_885_nl : STD_LOGIC;
  SIGNAL or_747_nl : STD_LOGIC;
  SIGNAL mux_884_nl : STD_LOGIC;
  SIGNAL or_744_nl : STD_LOGIC;
  SIGNAL mux_883_nl : STD_LOGIC;
  SIGNAL mux_882_nl : STD_LOGIC;
  SIGNAL or_741_nl : STD_LOGIC;
  SIGNAL mux_881_nl : STD_LOGIC;
  SIGNAL or_738_nl : STD_LOGIC;
  SIGNAL mux_910_nl : STD_LOGIC;
  SIGNAL mux_909_nl : STD_LOGIC;
  SIGNAL or_781_nl : STD_LOGIC;
  SIGNAL mux_908_nl : STD_LOGIC;
  SIGNAL or_780_nl : STD_LOGIC;
  SIGNAL or_779_nl : STD_LOGIC;
  SIGNAL mux_907_nl : STD_LOGIC;
  SIGNAL mux_906_nl : STD_LOGIC;
  SIGNAL mux_905_nl : STD_LOGIC;
  SIGNAL or_777_nl : STD_LOGIC;
  SIGNAL mux_904_nl : STD_LOGIC;
  SIGNAL or_775_nl : STD_LOGIC;
  SIGNAL mux_903_nl : STD_LOGIC;
  SIGNAL mux_902_nl : STD_LOGIC;
  SIGNAL or_774_nl : STD_LOGIC;
  SIGNAL mux_901_nl : STD_LOGIC;
  SIGNAL or_772_nl : STD_LOGIC;
  SIGNAL or_771_nl : STD_LOGIC;
  SIGNAL mux_900_nl : STD_LOGIC;
  SIGNAL mux_899_nl : STD_LOGIC;
  SIGNAL mux_898_nl : STD_LOGIC;
  SIGNAL or_770_nl : STD_LOGIC;
  SIGNAL or_768_nl : STD_LOGIC;
  SIGNAL mux_897_nl : STD_LOGIC;
  SIGNAL or_766_nl : STD_LOGIC;
  SIGNAL or_765_nl : STD_LOGIC;
  SIGNAL nand_21_nl : STD_LOGIC;
  SIGNAL mux_896_nl : STD_LOGIC;
  SIGNAL nor_1379_nl : STD_LOGIC;
  SIGNAL nor_1380_nl : STD_LOGIC;
  SIGNAL mux_925_nl : STD_LOGIC;
  SIGNAL nand_465_nl : STD_LOGIC;
  SIGNAL mux_924_nl : STD_LOGIC;
  SIGNAL mux_923_nl : STD_LOGIC;
  SIGNAL mux_922_nl : STD_LOGIC;
  SIGNAL nor_1370_nl : STD_LOGIC;
  SIGNAL nor_1371_nl : STD_LOGIC;
  SIGNAL mux_921_nl : STD_LOGIC;
  SIGNAL nor_1372_nl : STD_LOGIC;
  SIGNAL nor_1373_nl : STD_LOGIC;
  SIGNAL mux_920_nl : STD_LOGIC;
  SIGNAL mux_919_nl : STD_LOGIC;
  SIGNAL nor_1374_nl : STD_LOGIC;
  SIGNAL nor_1375_nl : STD_LOGIC;
  SIGNAL mux_918_nl : STD_LOGIC;
  SIGNAL nor_1376_nl : STD_LOGIC;
  SIGNAL nor_1377_nl : STD_LOGIC;
  SIGNAL or_4138_nl : STD_LOGIC;
  SIGNAL mux_917_nl : STD_LOGIC;
  SIGNAL mux_916_nl : STD_LOGIC;
  SIGNAL mux_915_nl : STD_LOGIC;
  SIGNAL or_791_nl : STD_LOGIC;
  SIGNAL mux_914_nl : STD_LOGIC;
  SIGNAL or_788_nl : STD_LOGIC;
  SIGNAL mux_913_nl : STD_LOGIC;
  SIGNAL mux_912_nl : STD_LOGIC;
  SIGNAL or_785_nl : STD_LOGIC;
  SIGNAL mux_911_nl : STD_LOGIC;
  SIGNAL or_782_nl : STD_LOGIC;
  SIGNAL mux_940_nl : STD_LOGIC;
  SIGNAL mux_939_nl : STD_LOGIC;
  SIGNAL or_825_nl : STD_LOGIC;
  SIGNAL mux_938_nl : STD_LOGIC;
  SIGNAL or_824_nl : STD_LOGIC;
  SIGNAL or_823_nl : STD_LOGIC;
  SIGNAL mux_937_nl : STD_LOGIC;
  SIGNAL mux_936_nl : STD_LOGIC;
  SIGNAL mux_935_nl : STD_LOGIC;
  SIGNAL or_821_nl : STD_LOGIC;
  SIGNAL mux_934_nl : STD_LOGIC;
  SIGNAL or_819_nl : STD_LOGIC;
  SIGNAL mux_933_nl : STD_LOGIC;
  SIGNAL mux_932_nl : STD_LOGIC;
  SIGNAL or_818_nl : STD_LOGIC;
  SIGNAL mux_931_nl : STD_LOGIC;
  SIGNAL or_816_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL mux_930_nl : STD_LOGIC;
  SIGNAL mux_929_nl : STD_LOGIC;
  SIGNAL mux_928_nl : STD_LOGIC;
  SIGNAL or_814_nl : STD_LOGIC;
  SIGNAL or_812_nl : STD_LOGIC;
  SIGNAL mux_927_nl : STD_LOGIC;
  SIGNAL or_810_nl : STD_LOGIC;
  SIGNAL or_809_nl : STD_LOGIC;
  SIGNAL nand_23_nl : STD_LOGIC;
  SIGNAL mux_926_nl : STD_LOGIC;
  SIGNAL nor_1368_nl : STD_LOGIC;
  SIGNAL nor_1369_nl : STD_LOGIC;
  SIGNAL mux_955_nl : STD_LOGIC;
  SIGNAL nand_464_nl : STD_LOGIC;
  SIGNAL mux_954_nl : STD_LOGIC;
  SIGNAL mux_953_nl : STD_LOGIC;
  SIGNAL mux_952_nl : STD_LOGIC;
  SIGNAL nor_1359_nl : STD_LOGIC;
  SIGNAL nor_1360_nl : STD_LOGIC;
  SIGNAL mux_951_nl : STD_LOGIC;
  SIGNAL nor_1361_nl : STD_LOGIC;
  SIGNAL nor_1362_nl : STD_LOGIC;
  SIGNAL mux_950_nl : STD_LOGIC;
  SIGNAL mux_949_nl : STD_LOGIC;
  SIGNAL nor_1363_nl : STD_LOGIC;
  SIGNAL nor_1364_nl : STD_LOGIC;
  SIGNAL mux_948_nl : STD_LOGIC;
  SIGNAL nor_1365_nl : STD_LOGIC;
  SIGNAL nor_1366_nl : STD_LOGIC;
  SIGNAL or_4137_nl : STD_LOGIC;
  SIGNAL mux_947_nl : STD_LOGIC;
  SIGNAL mux_946_nl : STD_LOGIC;
  SIGNAL mux_945_nl : STD_LOGIC;
  SIGNAL or_835_nl : STD_LOGIC;
  SIGNAL mux_944_nl : STD_LOGIC;
  SIGNAL or_832_nl : STD_LOGIC;
  SIGNAL mux_943_nl : STD_LOGIC;
  SIGNAL mux_942_nl : STD_LOGIC;
  SIGNAL or_829_nl : STD_LOGIC;
  SIGNAL mux_941_nl : STD_LOGIC;
  SIGNAL or_826_nl : STD_LOGIC;
  SIGNAL mux_970_nl : STD_LOGIC;
  SIGNAL mux_969_nl : STD_LOGIC;
  SIGNAL or_869_nl : STD_LOGIC;
  SIGNAL mux_968_nl : STD_LOGIC;
  SIGNAL or_868_nl : STD_LOGIC;
  SIGNAL or_867_nl : STD_LOGIC;
  SIGNAL mux_967_nl : STD_LOGIC;
  SIGNAL mux_966_nl : STD_LOGIC;
  SIGNAL mux_965_nl : STD_LOGIC;
  SIGNAL or_865_nl : STD_LOGIC;
  SIGNAL mux_964_nl : STD_LOGIC;
  SIGNAL or_863_nl : STD_LOGIC;
  SIGNAL mux_963_nl : STD_LOGIC;
  SIGNAL mux_962_nl : STD_LOGIC;
  SIGNAL or_862_nl : STD_LOGIC;
  SIGNAL mux_961_nl : STD_LOGIC;
  SIGNAL or_860_nl : STD_LOGIC;
  SIGNAL or_859_nl : STD_LOGIC;
  SIGNAL mux_960_nl : STD_LOGIC;
  SIGNAL mux_959_nl : STD_LOGIC;
  SIGNAL mux_958_nl : STD_LOGIC;
  SIGNAL or_858_nl : STD_LOGIC;
  SIGNAL or_856_nl : STD_LOGIC;
  SIGNAL mux_957_nl : STD_LOGIC;
  SIGNAL or_854_nl : STD_LOGIC;
  SIGNAL or_853_nl : STD_LOGIC;
  SIGNAL nand_25_nl : STD_LOGIC;
  SIGNAL mux_956_nl : STD_LOGIC;
  SIGNAL nor_1357_nl : STD_LOGIC;
  SIGNAL nor_1358_nl : STD_LOGIC;
  SIGNAL mux_985_nl : STD_LOGIC;
  SIGNAL nand_463_nl : STD_LOGIC;
  SIGNAL mux_984_nl : STD_LOGIC;
  SIGNAL mux_983_nl : STD_LOGIC;
  SIGNAL mux_982_nl : STD_LOGIC;
  SIGNAL nor_1348_nl : STD_LOGIC;
  SIGNAL nor_1349_nl : STD_LOGIC;
  SIGNAL mux_981_nl : STD_LOGIC;
  SIGNAL nor_1350_nl : STD_LOGIC;
  SIGNAL nor_1351_nl : STD_LOGIC;
  SIGNAL mux_980_nl : STD_LOGIC;
  SIGNAL mux_979_nl : STD_LOGIC;
  SIGNAL nor_1352_nl : STD_LOGIC;
  SIGNAL nor_1353_nl : STD_LOGIC;
  SIGNAL mux_978_nl : STD_LOGIC;
  SIGNAL nor_1354_nl : STD_LOGIC;
  SIGNAL nor_1355_nl : STD_LOGIC;
  SIGNAL or_4136_nl : STD_LOGIC;
  SIGNAL mux_977_nl : STD_LOGIC;
  SIGNAL mux_976_nl : STD_LOGIC;
  SIGNAL mux_975_nl : STD_LOGIC;
  SIGNAL or_879_nl : STD_LOGIC;
  SIGNAL mux_974_nl : STD_LOGIC;
  SIGNAL or_876_nl : STD_LOGIC;
  SIGNAL mux_973_nl : STD_LOGIC;
  SIGNAL mux_972_nl : STD_LOGIC;
  SIGNAL or_873_nl : STD_LOGIC;
  SIGNAL mux_971_nl : STD_LOGIC;
  SIGNAL or_870_nl : STD_LOGIC;
  SIGNAL mux_1000_nl : STD_LOGIC;
  SIGNAL mux_999_nl : STD_LOGIC;
  SIGNAL or_913_nl : STD_LOGIC;
  SIGNAL mux_998_nl : STD_LOGIC;
  SIGNAL or_912_nl : STD_LOGIC;
  SIGNAL or_911_nl : STD_LOGIC;
  SIGNAL mux_997_nl : STD_LOGIC;
  SIGNAL mux_996_nl : STD_LOGIC;
  SIGNAL mux_995_nl : STD_LOGIC;
  SIGNAL or_909_nl : STD_LOGIC;
  SIGNAL mux_994_nl : STD_LOGIC;
  SIGNAL or_907_nl : STD_LOGIC;
  SIGNAL mux_993_nl : STD_LOGIC;
  SIGNAL mux_992_nl : STD_LOGIC;
  SIGNAL or_906_nl : STD_LOGIC;
  SIGNAL mux_991_nl : STD_LOGIC;
  SIGNAL or_904_nl : STD_LOGIC;
  SIGNAL or_903_nl : STD_LOGIC;
  SIGNAL mux_990_nl : STD_LOGIC;
  SIGNAL mux_989_nl : STD_LOGIC;
  SIGNAL mux_988_nl : STD_LOGIC;
  SIGNAL or_902_nl : STD_LOGIC;
  SIGNAL or_900_nl : STD_LOGIC;
  SIGNAL mux_987_nl : STD_LOGIC;
  SIGNAL or_898_nl : STD_LOGIC;
  SIGNAL or_897_nl : STD_LOGIC;
  SIGNAL nand_27_nl : STD_LOGIC;
  SIGNAL mux_986_nl : STD_LOGIC;
  SIGNAL nor_1346_nl : STD_LOGIC;
  SIGNAL nor_1347_nl : STD_LOGIC;
  SIGNAL mux_1015_nl : STD_LOGIC;
  SIGNAL nand_462_nl : STD_LOGIC;
  SIGNAL mux_1014_nl : STD_LOGIC;
  SIGNAL mux_1013_nl : STD_LOGIC;
  SIGNAL mux_1012_nl : STD_LOGIC;
  SIGNAL nor_1337_nl : STD_LOGIC;
  SIGNAL nor_1338_nl : STD_LOGIC;
  SIGNAL mux_1011_nl : STD_LOGIC;
  SIGNAL nor_1339_nl : STD_LOGIC;
  SIGNAL nor_1340_nl : STD_LOGIC;
  SIGNAL mux_1010_nl : STD_LOGIC;
  SIGNAL mux_1009_nl : STD_LOGIC;
  SIGNAL nor_1341_nl : STD_LOGIC;
  SIGNAL nor_1342_nl : STD_LOGIC;
  SIGNAL mux_1008_nl : STD_LOGIC;
  SIGNAL nor_1343_nl : STD_LOGIC;
  SIGNAL nor_1344_nl : STD_LOGIC;
  SIGNAL or_4135_nl : STD_LOGIC;
  SIGNAL mux_1007_nl : STD_LOGIC;
  SIGNAL mux_1006_nl : STD_LOGIC;
  SIGNAL mux_1005_nl : STD_LOGIC;
  SIGNAL or_923_nl : STD_LOGIC;
  SIGNAL mux_1004_nl : STD_LOGIC;
  SIGNAL or_920_nl : STD_LOGIC;
  SIGNAL mux_1003_nl : STD_LOGIC;
  SIGNAL mux_1002_nl : STD_LOGIC;
  SIGNAL or_917_nl : STD_LOGIC;
  SIGNAL mux_1001_nl : STD_LOGIC;
  SIGNAL or_914_nl : STD_LOGIC;
  SIGNAL mux_1030_nl : STD_LOGIC;
  SIGNAL mux_1029_nl : STD_LOGIC;
  SIGNAL or_957_nl : STD_LOGIC;
  SIGNAL mux_1028_nl : STD_LOGIC;
  SIGNAL or_956_nl : STD_LOGIC;
  SIGNAL or_955_nl : STD_LOGIC;
  SIGNAL mux_1027_nl : STD_LOGIC;
  SIGNAL mux_1026_nl : STD_LOGIC;
  SIGNAL mux_1025_nl : STD_LOGIC;
  SIGNAL or_953_nl : STD_LOGIC;
  SIGNAL mux_1024_nl : STD_LOGIC;
  SIGNAL or_951_nl : STD_LOGIC;
  SIGNAL mux_1023_nl : STD_LOGIC;
  SIGNAL mux_1022_nl : STD_LOGIC;
  SIGNAL or_950_nl : STD_LOGIC;
  SIGNAL mux_1021_nl : STD_LOGIC;
  SIGNAL or_948_nl : STD_LOGIC;
  SIGNAL or_947_nl : STD_LOGIC;
  SIGNAL mux_1020_nl : STD_LOGIC;
  SIGNAL mux_1019_nl : STD_LOGIC;
  SIGNAL mux_1018_nl : STD_LOGIC;
  SIGNAL or_946_nl : STD_LOGIC;
  SIGNAL or_944_nl : STD_LOGIC;
  SIGNAL mux_1017_nl : STD_LOGIC;
  SIGNAL or_942_nl : STD_LOGIC;
  SIGNAL or_941_nl : STD_LOGIC;
  SIGNAL nand_29_nl : STD_LOGIC;
  SIGNAL mux_1016_nl : STD_LOGIC;
  SIGNAL nor_1335_nl : STD_LOGIC;
  SIGNAL nor_1336_nl : STD_LOGIC;
  SIGNAL mux_1045_nl : STD_LOGIC;
  SIGNAL nand_461_nl : STD_LOGIC;
  SIGNAL mux_1044_nl : STD_LOGIC;
  SIGNAL mux_1043_nl : STD_LOGIC;
  SIGNAL mux_1042_nl : STD_LOGIC;
  SIGNAL nor_1326_nl : STD_LOGIC;
  SIGNAL nor_1327_nl : STD_LOGIC;
  SIGNAL mux_1041_nl : STD_LOGIC;
  SIGNAL nor_1328_nl : STD_LOGIC;
  SIGNAL nor_1329_nl : STD_LOGIC;
  SIGNAL mux_1040_nl : STD_LOGIC;
  SIGNAL mux_1039_nl : STD_LOGIC;
  SIGNAL nor_1330_nl : STD_LOGIC;
  SIGNAL nor_1331_nl : STD_LOGIC;
  SIGNAL mux_1038_nl : STD_LOGIC;
  SIGNAL nor_1332_nl : STD_LOGIC;
  SIGNAL nor_1333_nl : STD_LOGIC;
  SIGNAL or_4134_nl : STD_LOGIC;
  SIGNAL mux_1037_nl : STD_LOGIC;
  SIGNAL mux_1036_nl : STD_LOGIC;
  SIGNAL mux_1035_nl : STD_LOGIC;
  SIGNAL or_967_nl : STD_LOGIC;
  SIGNAL mux_1034_nl : STD_LOGIC;
  SIGNAL or_964_nl : STD_LOGIC;
  SIGNAL mux_1033_nl : STD_LOGIC;
  SIGNAL mux_1032_nl : STD_LOGIC;
  SIGNAL or_961_nl : STD_LOGIC;
  SIGNAL mux_1031_nl : STD_LOGIC;
  SIGNAL or_958_nl : STD_LOGIC;
  SIGNAL mux_1060_nl : STD_LOGIC;
  SIGNAL mux_1059_nl : STD_LOGIC;
  SIGNAL or_1001_nl : STD_LOGIC;
  SIGNAL mux_1058_nl : STD_LOGIC;
  SIGNAL or_1000_nl : STD_LOGIC;
  SIGNAL or_999_nl : STD_LOGIC;
  SIGNAL mux_1057_nl : STD_LOGIC;
  SIGNAL mux_1056_nl : STD_LOGIC;
  SIGNAL mux_1055_nl : STD_LOGIC;
  SIGNAL or_997_nl : STD_LOGIC;
  SIGNAL mux_1054_nl : STD_LOGIC;
  SIGNAL or_995_nl : STD_LOGIC;
  SIGNAL mux_1053_nl : STD_LOGIC;
  SIGNAL mux_1052_nl : STD_LOGIC;
  SIGNAL or_994_nl : STD_LOGIC;
  SIGNAL mux_1051_nl : STD_LOGIC;
  SIGNAL or_992_nl : STD_LOGIC;
  SIGNAL or_991_nl : STD_LOGIC;
  SIGNAL mux_1050_nl : STD_LOGIC;
  SIGNAL mux_1049_nl : STD_LOGIC;
  SIGNAL mux_1048_nl : STD_LOGIC;
  SIGNAL or_990_nl : STD_LOGIC;
  SIGNAL or_988_nl : STD_LOGIC;
  SIGNAL mux_1047_nl : STD_LOGIC;
  SIGNAL or_986_nl : STD_LOGIC;
  SIGNAL or_985_nl : STD_LOGIC;
  SIGNAL nand_31_nl : STD_LOGIC;
  SIGNAL mux_1046_nl : STD_LOGIC;
  SIGNAL nor_1324_nl : STD_LOGIC;
  SIGNAL nor_1325_nl : STD_LOGIC;
  SIGNAL mux_1075_nl : STD_LOGIC;
  SIGNAL nand_460_nl : STD_LOGIC;
  SIGNAL mux_1074_nl : STD_LOGIC;
  SIGNAL mux_1073_nl : STD_LOGIC;
  SIGNAL mux_1072_nl : STD_LOGIC;
  SIGNAL nor_1315_nl : STD_LOGIC;
  SIGNAL nor_1316_nl : STD_LOGIC;
  SIGNAL mux_1071_nl : STD_LOGIC;
  SIGNAL nor_1317_nl : STD_LOGIC;
  SIGNAL nor_1318_nl : STD_LOGIC;
  SIGNAL mux_1070_nl : STD_LOGIC;
  SIGNAL mux_1069_nl : STD_LOGIC;
  SIGNAL nor_1319_nl : STD_LOGIC;
  SIGNAL nor_1320_nl : STD_LOGIC;
  SIGNAL mux_1068_nl : STD_LOGIC;
  SIGNAL nor_1321_nl : STD_LOGIC;
  SIGNAL nor_1322_nl : STD_LOGIC;
  SIGNAL or_4133_nl : STD_LOGIC;
  SIGNAL mux_1067_nl : STD_LOGIC;
  SIGNAL mux_1066_nl : STD_LOGIC;
  SIGNAL mux_1065_nl : STD_LOGIC;
  SIGNAL or_1011_nl : STD_LOGIC;
  SIGNAL mux_1064_nl : STD_LOGIC;
  SIGNAL or_1008_nl : STD_LOGIC;
  SIGNAL mux_1063_nl : STD_LOGIC;
  SIGNAL mux_1062_nl : STD_LOGIC;
  SIGNAL or_1005_nl : STD_LOGIC;
  SIGNAL mux_1061_nl : STD_LOGIC;
  SIGNAL or_1002_nl : STD_LOGIC;
  SIGNAL mux_1090_nl : STD_LOGIC;
  SIGNAL mux_1089_nl : STD_LOGIC;
  SIGNAL or_1045_nl : STD_LOGIC;
  SIGNAL mux_1088_nl : STD_LOGIC;
  SIGNAL or_1044_nl : STD_LOGIC;
  SIGNAL or_1043_nl : STD_LOGIC;
  SIGNAL mux_1087_nl : STD_LOGIC;
  SIGNAL mux_1086_nl : STD_LOGIC;
  SIGNAL mux_1085_nl : STD_LOGIC;
  SIGNAL or_1041_nl : STD_LOGIC;
  SIGNAL mux_1084_nl : STD_LOGIC;
  SIGNAL or_1039_nl : STD_LOGIC;
  SIGNAL mux_1083_nl : STD_LOGIC;
  SIGNAL mux_1082_nl : STD_LOGIC;
  SIGNAL or_1038_nl : STD_LOGIC;
  SIGNAL mux_1081_nl : STD_LOGIC;
  SIGNAL or_1036_nl : STD_LOGIC;
  SIGNAL or_1035_nl : STD_LOGIC;
  SIGNAL mux_1080_nl : STD_LOGIC;
  SIGNAL mux_1079_nl : STD_LOGIC;
  SIGNAL mux_1078_nl : STD_LOGIC;
  SIGNAL or_1034_nl : STD_LOGIC;
  SIGNAL or_1032_nl : STD_LOGIC;
  SIGNAL mux_1077_nl : STD_LOGIC;
  SIGNAL or_1030_nl : STD_LOGIC;
  SIGNAL or_1029_nl : STD_LOGIC;
  SIGNAL nand_33_nl : STD_LOGIC;
  SIGNAL mux_1076_nl : STD_LOGIC;
  SIGNAL nor_1313_nl : STD_LOGIC;
  SIGNAL nor_1314_nl : STD_LOGIC;
  SIGNAL mux_1105_nl : STD_LOGIC;
  SIGNAL nand_459_nl : STD_LOGIC;
  SIGNAL mux_1104_nl : STD_LOGIC;
  SIGNAL mux_1103_nl : STD_LOGIC;
  SIGNAL mux_1102_nl : STD_LOGIC;
  SIGNAL nor_1304_nl : STD_LOGIC;
  SIGNAL nor_1305_nl : STD_LOGIC;
  SIGNAL mux_1101_nl : STD_LOGIC;
  SIGNAL nor_1306_nl : STD_LOGIC;
  SIGNAL nor_1307_nl : STD_LOGIC;
  SIGNAL mux_1100_nl : STD_LOGIC;
  SIGNAL mux_1099_nl : STD_LOGIC;
  SIGNAL nor_1308_nl : STD_LOGIC;
  SIGNAL nor_1309_nl : STD_LOGIC;
  SIGNAL mux_1098_nl : STD_LOGIC;
  SIGNAL nor_1310_nl : STD_LOGIC;
  SIGNAL nor_1311_nl : STD_LOGIC;
  SIGNAL or_4132_nl : STD_LOGIC;
  SIGNAL mux_1097_nl : STD_LOGIC;
  SIGNAL mux_1096_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL or_1055_nl : STD_LOGIC;
  SIGNAL mux_1094_nl : STD_LOGIC;
  SIGNAL or_1052_nl : STD_LOGIC;
  SIGNAL mux_1093_nl : STD_LOGIC;
  SIGNAL mux_1092_nl : STD_LOGIC;
  SIGNAL or_1049_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL or_1046_nl : STD_LOGIC;
  SIGNAL mux_1120_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL or_1089_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL or_1088_nl : STD_LOGIC;
  SIGNAL or_1087_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL mux_1116_nl : STD_LOGIC;
  SIGNAL mux_1115_nl : STD_LOGIC;
  SIGNAL or_1085_nl : STD_LOGIC;
  SIGNAL mux_1114_nl : STD_LOGIC;
  SIGNAL or_1083_nl : STD_LOGIC;
  SIGNAL mux_1113_nl : STD_LOGIC;
  SIGNAL mux_1112_nl : STD_LOGIC;
  SIGNAL or_1082_nl : STD_LOGIC;
  SIGNAL mux_1111_nl : STD_LOGIC;
  SIGNAL or_1080_nl : STD_LOGIC;
  SIGNAL or_1079_nl : STD_LOGIC;
  SIGNAL mux_1110_nl : STD_LOGIC;
  SIGNAL mux_1109_nl : STD_LOGIC;
  SIGNAL mux_1108_nl : STD_LOGIC;
  SIGNAL or_1078_nl : STD_LOGIC;
  SIGNAL or_1076_nl : STD_LOGIC;
  SIGNAL mux_1107_nl : STD_LOGIC;
  SIGNAL or_1074_nl : STD_LOGIC;
  SIGNAL or_1073_nl : STD_LOGIC;
  SIGNAL nand_35_nl : STD_LOGIC;
  SIGNAL mux_1106_nl : STD_LOGIC;
  SIGNAL nor_1302_nl : STD_LOGIC;
  SIGNAL nor_1303_nl : STD_LOGIC;
  SIGNAL mux_1135_nl : STD_LOGIC;
  SIGNAL nand_458_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL mux_1132_nl : STD_LOGIC;
  SIGNAL nor_1293_nl : STD_LOGIC;
  SIGNAL nor_1294_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL nor_1295_nl : STD_LOGIC;
  SIGNAL nor_1296_nl : STD_LOGIC;
  SIGNAL mux_1130_nl : STD_LOGIC;
  SIGNAL mux_1129_nl : STD_LOGIC;
  SIGNAL nor_1297_nl : STD_LOGIC;
  SIGNAL nor_1298_nl : STD_LOGIC;
  SIGNAL mux_1128_nl : STD_LOGIC;
  SIGNAL nor_1299_nl : STD_LOGIC;
  SIGNAL nor_1300_nl : STD_LOGIC;
  SIGNAL or_4131_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL mux_1125_nl : STD_LOGIC;
  SIGNAL or_1099_nl : STD_LOGIC;
  SIGNAL mux_1124_nl : STD_LOGIC;
  SIGNAL or_1096_nl : STD_LOGIC;
  SIGNAL mux_1123_nl : STD_LOGIC;
  SIGNAL mux_1122_nl : STD_LOGIC;
  SIGNAL or_1093_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL or_1090_nl : STD_LOGIC;
  SIGNAL mux_1150_nl : STD_LOGIC;
  SIGNAL mux_1149_nl : STD_LOGIC;
  SIGNAL or_1133_nl : STD_LOGIC;
  SIGNAL mux_1148_nl : STD_LOGIC;
  SIGNAL or_1132_nl : STD_LOGIC;
  SIGNAL or_1131_nl : STD_LOGIC;
  SIGNAL mux_1147_nl : STD_LOGIC;
  SIGNAL mux_1146_nl : STD_LOGIC;
  SIGNAL mux_1145_nl : STD_LOGIC;
  SIGNAL or_1129_nl : STD_LOGIC;
  SIGNAL mux_1144_nl : STD_LOGIC;
  SIGNAL or_1127_nl : STD_LOGIC;
  SIGNAL mux_1143_nl : STD_LOGIC;
  SIGNAL mux_1142_nl : STD_LOGIC;
  SIGNAL or_1126_nl : STD_LOGIC;
  SIGNAL mux_1141_nl : STD_LOGIC;
  SIGNAL or_1124_nl : STD_LOGIC;
  SIGNAL or_1123_nl : STD_LOGIC;
  SIGNAL mux_1140_nl : STD_LOGIC;
  SIGNAL mux_1139_nl : STD_LOGIC;
  SIGNAL mux_1138_nl : STD_LOGIC;
  SIGNAL or_1122_nl : STD_LOGIC;
  SIGNAL or_1120_nl : STD_LOGIC;
  SIGNAL mux_1137_nl : STD_LOGIC;
  SIGNAL or_1118_nl : STD_LOGIC;
  SIGNAL or_1117_nl : STD_LOGIC;
  SIGNAL nand_37_nl : STD_LOGIC;
  SIGNAL mux_1136_nl : STD_LOGIC;
  SIGNAL nor_1291_nl : STD_LOGIC;
  SIGNAL nor_1292_nl : STD_LOGIC;
  SIGNAL mux_1165_nl : STD_LOGIC;
  SIGNAL nand_457_nl : STD_LOGIC;
  SIGNAL mux_1164_nl : STD_LOGIC;
  SIGNAL mux_1163_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL nor_1282_nl : STD_LOGIC;
  SIGNAL nor_1283_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL nor_1284_nl : STD_LOGIC;
  SIGNAL nor_1285_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL mux_1159_nl : STD_LOGIC;
  SIGNAL nor_1286_nl : STD_LOGIC;
  SIGNAL nor_1287_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL nor_1288_nl : STD_LOGIC;
  SIGNAL nor_1289_nl : STD_LOGIC;
  SIGNAL or_4130_nl : STD_LOGIC;
  SIGNAL mux_1157_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL mux_1155_nl : STD_LOGIC;
  SIGNAL or_1143_nl : STD_LOGIC;
  SIGNAL mux_1154_nl : STD_LOGIC;
  SIGNAL or_1140_nl : STD_LOGIC;
  SIGNAL mux_1153_nl : STD_LOGIC;
  SIGNAL mux_1152_nl : STD_LOGIC;
  SIGNAL or_1137_nl : STD_LOGIC;
  SIGNAL mux_1151_nl : STD_LOGIC;
  SIGNAL or_1134_nl : STD_LOGIC;
  SIGNAL mux_1180_nl : STD_LOGIC;
  SIGNAL mux_1179_nl : STD_LOGIC;
  SIGNAL or_1177_nl : STD_LOGIC;
  SIGNAL mux_1178_nl : STD_LOGIC;
  SIGNAL or_1176_nl : STD_LOGIC;
  SIGNAL or_1175_nl : STD_LOGIC;
  SIGNAL mux_1177_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL mux_1175_nl : STD_LOGIC;
  SIGNAL or_1173_nl : STD_LOGIC;
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL or_1171_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL mux_1172_nl : STD_LOGIC;
  SIGNAL or_1170_nl : STD_LOGIC;
  SIGNAL mux_1171_nl : STD_LOGIC;
  SIGNAL or_1168_nl : STD_LOGIC;
  SIGNAL or_1167_nl : STD_LOGIC;
  SIGNAL mux_1170_nl : STD_LOGIC;
  SIGNAL mux_1169_nl : STD_LOGIC;
  SIGNAL mux_1168_nl : STD_LOGIC;
  SIGNAL or_1166_nl : STD_LOGIC;
  SIGNAL or_1164_nl : STD_LOGIC;
  SIGNAL mux_1167_nl : STD_LOGIC;
  SIGNAL or_1162_nl : STD_LOGIC;
  SIGNAL or_1161_nl : STD_LOGIC;
  SIGNAL nand_39_nl : STD_LOGIC;
  SIGNAL mux_1166_nl : STD_LOGIC;
  SIGNAL nor_1280_nl : STD_LOGIC;
  SIGNAL nor_1281_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL nand_456_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL nor_1271_nl : STD_LOGIC;
  SIGNAL nor_1272_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL nor_1273_nl : STD_LOGIC;
  SIGNAL nor_1274_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL nor_1275_nl : STD_LOGIC;
  SIGNAL nor_1276_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL nor_1277_nl : STD_LOGIC;
  SIGNAL nor_1278_nl : STD_LOGIC;
  SIGNAL or_4129_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL mux_1185_nl : STD_LOGIC;
  SIGNAL or_1187_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL or_1184_nl : STD_LOGIC;
  SIGNAL mux_1183_nl : STD_LOGIC;
  SIGNAL mux_1182_nl : STD_LOGIC;
  SIGNAL or_1181_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL or_1178_nl : STD_LOGIC;
  SIGNAL mux_1210_nl : STD_LOGIC;
  SIGNAL mux_1209_nl : STD_LOGIC;
  SIGNAL or_1221_nl : STD_LOGIC;
  SIGNAL mux_1208_nl : STD_LOGIC;
  SIGNAL or_1220_nl : STD_LOGIC;
  SIGNAL or_1219_nl : STD_LOGIC;
  SIGNAL mux_1207_nl : STD_LOGIC;
  SIGNAL mux_1206_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL or_1217_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL or_1215_nl : STD_LOGIC;
  SIGNAL mux_1203_nl : STD_LOGIC;
  SIGNAL mux_1202_nl : STD_LOGIC;
  SIGNAL or_1214_nl : STD_LOGIC;
  SIGNAL mux_1201_nl : STD_LOGIC;
  SIGNAL or_1212_nl : STD_LOGIC;
  SIGNAL or_1211_nl : STD_LOGIC;
  SIGNAL mux_1200_nl : STD_LOGIC;
  SIGNAL mux_1199_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL or_1210_nl : STD_LOGIC;
  SIGNAL or_1208_nl : STD_LOGIC;
  SIGNAL mux_1197_nl : STD_LOGIC;
  SIGNAL or_1206_nl : STD_LOGIC;
  SIGNAL or_1205_nl : STD_LOGIC;
  SIGNAL nand_41_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL nor_1269_nl : STD_LOGIC;
  SIGNAL nor_1270_nl : STD_LOGIC;
  SIGNAL mux_1225_nl : STD_LOGIC;
  SIGNAL nand_455_nl : STD_LOGIC;
  SIGNAL mux_1224_nl : STD_LOGIC;
  SIGNAL mux_1223_nl : STD_LOGIC;
  SIGNAL mux_1222_nl : STD_LOGIC;
  SIGNAL nor_1260_nl : STD_LOGIC;
  SIGNAL nor_1261_nl : STD_LOGIC;
  SIGNAL mux_1221_nl : STD_LOGIC;
  SIGNAL nor_1262_nl : STD_LOGIC;
  SIGNAL nor_1263_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL mux_1219_nl : STD_LOGIC;
  SIGNAL nor_1264_nl : STD_LOGIC;
  SIGNAL nor_1265_nl : STD_LOGIC;
  SIGNAL mux_1218_nl : STD_LOGIC;
  SIGNAL nor_1266_nl : STD_LOGIC;
  SIGNAL nor_1267_nl : STD_LOGIC;
  SIGNAL or_4128_nl : STD_LOGIC;
  SIGNAL mux_1217_nl : STD_LOGIC;
  SIGNAL mux_1216_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL or_1231_nl : STD_LOGIC;
  SIGNAL mux_1214_nl : STD_LOGIC;
  SIGNAL or_1228_nl : STD_LOGIC;
  SIGNAL mux_1213_nl : STD_LOGIC;
  SIGNAL mux_1212_nl : STD_LOGIC;
  SIGNAL or_1225_nl : STD_LOGIC;
  SIGNAL mux_1211_nl : STD_LOGIC;
  SIGNAL or_1222_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL mux_1239_nl : STD_LOGIC;
  SIGNAL or_1265_nl : STD_LOGIC;
  SIGNAL mux_1238_nl : STD_LOGIC;
  SIGNAL or_1264_nl : STD_LOGIC;
  SIGNAL or_1263_nl : STD_LOGIC;
  SIGNAL mux_1237_nl : STD_LOGIC;
  SIGNAL mux_1236_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL or_1261_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL or_1259_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL mux_1232_nl : STD_LOGIC;
  SIGNAL or_1258_nl : STD_LOGIC;
  SIGNAL mux_1231_nl : STD_LOGIC;
  SIGNAL or_1256_nl : STD_LOGIC;
  SIGNAL or_1255_nl : STD_LOGIC;
  SIGNAL mux_1230_nl : STD_LOGIC;
  SIGNAL mux_1229_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL or_1254_nl : STD_LOGIC;
  SIGNAL or_1252_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL or_1250_nl : STD_LOGIC;
  SIGNAL or_1249_nl : STD_LOGIC;
  SIGNAL nand_43_nl : STD_LOGIC;
  SIGNAL mux_1226_nl : STD_LOGIC;
  SIGNAL nor_1258_nl : STD_LOGIC;
  SIGNAL nor_1259_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL nand_454_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL and_618_nl : STD_LOGIC;
  SIGNAL nor_1250_nl : STD_LOGIC;
  SIGNAL mux_1251_nl : STD_LOGIC;
  SIGNAL nor_1251_nl : STD_LOGIC;
  SIGNAL nor_1252_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL nor_1253_nl : STD_LOGIC;
  SIGNAL nor_1254_nl : STD_LOGIC;
  SIGNAL mux_1248_nl : STD_LOGIC;
  SIGNAL nor_1255_nl : STD_LOGIC;
  SIGNAL nor_1256_nl : STD_LOGIC;
  SIGNAL or_4127_nl : STD_LOGIC;
  SIGNAL mux_1247_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL mux_1245_nl : STD_LOGIC;
  SIGNAL nand_332_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL or_1272_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL or_1269_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL or_1266_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL or_1309_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL or_1308_nl : STD_LOGIC;
  SIGNAL or_1307_nl : STD_LOGIC;
  SIGNAL mux_1267_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL nand_330_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL or_1303_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL or_1302_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL or_1300_nl : STD_LOGIC;
  SIGNAL or_1299_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL or_1298_nl : STD_LOGIC;
  SIGNAL nand_331_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL or_1294_nl : STD_LOGIC;
  SIGNAL or_1293_nl : STD_LOGIC;
  SIGNAL nand_45_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL nor_1248_nl : STD_LOGIC;
  SIGNAL nor_1249_nl : STD_LOGIC;
  SIGNAL mux_1285_nl : STD_LOGIC;
  SIGNAL nand_453_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL mux_1283_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL nor_1239_nl : STD_LOGIC;
  SIGNAL nor_1240_nl : STD_LOGIC;
  SIGNAL mux_1281_nl : STD_LOGIC;
  SIGNAL nor_1241_nl : STD_LOGIC;
  SIGNAL nor_1242_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL nor_1243_nl : STD_LOGIC;
  SIGNAL nor_1244_nl : STD_LOGIC;
  SIGNAL mux_1278_nl : STD_LOGIC;
  SIGNAL nor_1245_nl : STD_LOGIC;
  SIGNAL nor_1246_nl : STD_LOGIC;
  SIGNAL or_4126_nl : STD_LOGIC;
  SIGNAL mux_1277_nl : STD_LOGIC;
  SIGNAL mux_1276_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL or_1319_nl : STD_LOGIC;
  SIGNAL mux_1274_nl : STD_LOGIC;
  SIGNAL or_1316_nl : STD_LOGIC;
  SIGNAL mux_1273_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL or_1313_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL or_1310_nl : STD_LOGIC;
  SIGNAL mux_1300_nl : STD_LOGIC;
  SIGNAL mux_1299_nl : STD_LOGIC;
  SIGNAL or_1353_nl : STD_LOGIC;
  SIGNAL mux_1298_nl : STD_LOGIC;
  SIGNAL or_1352_nl : STD_LOGIC;
  SIGNAL or_1351_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL mux_1296_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL or_1349_nl : STD_LOGIC;
  SIGNAL mux_1294_nl : STD_LOGIC;
  SIGNAL or_1347_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL mux_1292_nl : STD_LOGIC;
  SIGNAL or_1346_nl : STD_LOGIC;
  SIGNAL mux_1291_nl : STD_LOGIC;
  SIGNAL or_1344_nl : STD_LOGIC;
  SIGNAL or_1343_nl : STD_LOGIC;
  SIGNAL mux_1290_nl : STD_LOGIC;
  SIGNAL mux_1289_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL or_1342_nl : STD_LOGIC;
  SIGNAL or_1340_nl : STD_LOGIC;
  SIGNAL mux_1287_nl : STD_LOGIC;
  SIGNAL or_1338_nl : STD_LOGIC;
  SIGNAL or_1337_nl : STD_LOGIC;
  SIGNAL nand_47_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL nor_1237_nl : STD_LOGIC;
  SIGNAL nor_1238_nl : STD_LOGIC;
  SIGNAL mux_1315_nl : STD_LOGIC;
  SIGNAL nand_452_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL nor_1228_nl : STD_LOGIC;
  SIGNAL nor_1229_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL nor_1230_nl : STD_LOGIC;
  SIGNAL nor_1231_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL mux_1309_nl : STD_LOGIC;
  SIGNAL nor_1232_nl : STD_LOGIC;
  SIGNAL nor_1233_nl : STD_LOGIC;
  SIGNAL mux_1308_nl : STD_LOGIC;
  SIGNAL nor_1234_nl : STD_LOGIC;
  SIGNAL nor_1235_nl : STD_LOGIC;
  SIGNAL or_4125_nl : STD_LOGIC;
  SIGNAL mux_1307_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL mux_1305_nl : STD_LOGIC;
  SIGNAL or_1363_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL or_1360_nl : STD_LOGIC;
  SIGNAL mux_1303_nl : STD_LOGIC;
  SIGNAL mux_1302_nl : STD_LOGIC;
  SIGNAL or_1357_nl : STD_LOGIC;
  SIGNAL mux_1301_nl : STD_LOGIC;
  SIGNAL or_1354_nl : STD_LOGIC;
  SIGNAL mux_1330_nl : STD_LOGIC;
  SIGNAL mux_1329_nl : STD_LOGIC;
  SIGNAL or_1397_nl : STD_LOGIC;
  SIGNAL mux_1328_nl : STD_LOGIC;
  SIGNAL or_1396_nl : STD_LOGIC;
  SIGNAL or_1395_nl : STD_LOGIC;
  SIGNAL mux_1327_nl : STD_LOGIC;
  SIGNAL mux_1326_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL or_1393_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL or_1391_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL or_1390_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL or_1388_nl : STD_LOGIC;
  SIGNAL or_1387_nl : STD_LOGIC;
  SIGNAL mux_1320_nl : STD_LOGIC;
  SIGNAL mux_1319_nl : STD_LOGIC;
  SIGNAL mux_1318_nl : STD_LOGIC;
  SIGNAL or_1386_nl : STD_LOGIC;
  SIGNAL or_1384_nl : STD_LOGIC;
  SIGNAL mux_1317_nl : STD_LOGIC;
  SIGNAL or_1382_nl : STD_LOGIC;
  SIGNAL or_1381_nl : STD_LOGIC;
  SIGNAL nand_49_nl : STD_LOGIC;
  SIGNAL mux_1316_nl : STD_LOGIC;
  SIGNAL nor_1226_nl : STD_LOGIC;
  SIGNAL nor_1227_nl : STD_LOGIC;
  SIGNAL mux_1345_nl : STD_LOGIC;
  SIGNAL nand_451_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL mux_1343_nl : STD_LOGIC;
  SIGNAL mux_1342_nl : STD_LOGIC;
  SIGNAL nor_1217_nl : STD_LOGIC;
  SIGNAL nor_1218_nl : STD_LOGIC;
  SIGNAL mux_1341_nl : STD_LOGIC;
  SIGNAL nor_1219_nl : STD_LOGIC;
  SIGNAL nor_1220_nl : STD_LOGIC;
  SIGNAL mux_1340_nl : STD_LOGIC;
  SIGNAL mux_1339_nl : STD_LOGIC;
  SIGNAL nor_1221_nl : STD_LOGIC;
  SIGNAL nor_1222_nl : STD_LOGIC;
  SIGNAL mux_1338_nl : STD_LOGIC;
  SIGNAL nor_1223_nl : STD_LOGIC;
  SIGNAL nor_1224_nl : STD_LOGIC;
  SIGNAL or_4124_nl : STD_LOGIC;
  SIGNAL mux_1337_nl : STD_LOGIC;
  SIGNAL mux_1336_nl : STD_LOGIC;
  SIGNAL mux_1335_nl : STD_LOGIC;
  SIGNAL or_1407_nl : STD_LOGIC;
  SIGNAL mux_1334_nl : STD_LOGIC;
  SIGNAL or_1404_nl : STD_LOGIC;
  SIGNAL mux_1333_nl : STD_LOGIC;
  SIGNAL mux_1332_nl : STD_LOGIC;
  SIGNAL or_1401_nl : STD_LOGIC;
  SIGNAL mux_1331_nl : STD_LOGIC;
  SIGNAL or_1398_nl : STD_LOGIC;
  SIGNAL mux_1360_nl : STD_LOGIC;
  SIGNAL mux_1359_nl : STD_LOGIC;
  SIGNAL or_1441_nl : STD_LOGIC;
  SIGNAL mux_1358_nl : STD_LOGIC;
  SIGNAL or_1440_nl : STD_LOGIC;
  SIGNAL or_1439_nl : STD_LOGIC;
  SIGNAL mux_1357_nl : STD_LOGIC;
  SIGNAL mux_1356_nl : STD_LOGIC;
  SIGNAL mux_1355_nl : STD_LOGIC;
  SIGNAL or_1437_nl : STD_LOGIC;
  SIGNAL mux_1354_nl : STD_LOGIC;
  SIGNAL or_1435_nl : STD_LOGIC;
  SIGNAL mux_1353_nl : STD_LOGIC;
  SIGNAL mux_1352_nl : STD_LOGIC;
  SIGNAL or_1434_nl : STD_LOGIC;
  SIGNAL mux_1351_nl : STD_LOGIC;
  SIGNAL or_1432_nl : STD_LOGIC;
  SIGNAL or_1431_nl : STD_LOGIC;
  SIGNAL mux_1350_nl : STD_LOGIC;
  SIGNAL mux_1349_nl : STD_LOGIC;
  SIGNAL mux_1348_nl : STD_LOGIC;
  SIGNAL or_1430_nl : STD_LOGIC;
  SIGNAL or_1428_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL or_1426_nl : STD_LOGIC;
  SIGNAL or_1425_nl : STD_LOGIC;
  SIGNAL nand_51_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL nor_1215_nl : STD_LOGIC;
  SIGNAL nor_1216_nl : STD_LOGIC;
  SIGNAL mux_1375_nl : STD_LOGIC;
  SIGNAL nand_450_nl : STD_LOGIC;
  SIGNAL mux_1374_nl : STD_LOGIC;
  SIGNAL mux_1373_nl : STD_LOGIC;
  SIGNAL mux_1372_nl : STD_LOGIC;
  SIGNAL nor_1206_nl : STD_LOGIC;
  SIGNAL nor_1207_nl : STD_LOGIC;
  SIGNAL mux_1371_nl : STD_LOGIC;
  SIGNAL nor_1208_nl : STD_LOGIC;
  SIGNAL nor_1209_nl : STD_LOGIC;
  SIGNAL mux_1370_nl : STD_LOGIC;
  SIGNAL mux_1369_nl : STD_LOGIC;
  SIGNAL nor_1210_nl : STD_LOGIC;
  SIGNAL nor_1211_nl : STD_LOGIC;
  SIGNAL mux_1368_nl : STD_LOGIC;
  SIGNAL nor_1212_nl : STD_LOGIC;
  SIGNAL nor_1213_nl : STD_LOGIC;
  SIGNAL or_4123_nl : STD_LOGIC;
  SIGNAL mux_1367_nl : STD_LOGIC;
  SIGNAL mux_1366_nl : STD_LOGIC;
  SIGNAL mux_1365_nl : STD_LOGIC;
  SIGNAL or_1451_nl : STD_LOGIC;
  SIGNAL mux_1364_nl : STD_LOGIC;
  SIGNAL or_1448_nl : STD_LOGIC;
  SIGNAL mux_1363_nl : STD_LOGIC;
  SIGNAL mux_1362_nl : STD_LOGIC;
  SIGNAL or_1445_nl : STD_LOGIC;
  SIGNAL mux_1361_nl : STD_LOGIC;
  SIGNAL or_1442_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL mux_1389_nl : STD_LOGIC;
  SIGNAL or_1485_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL or_1484_nl : STD_LOGIC;
  SIGNAL or_1483_nl : STD_LOGIC;
  SIGNAL mux_1387_nl : STD_LOGIC;
  SIGNAL mux_1386_nl : STD_LOGIC;
  SIGNAL mux_1385_nl : STD_LOGIC;
  SIGNAL or_1481_nl : STD_LOGIC;
  SIGNAL mux_1384_nl : STD_LOGIC;
  SIGNAL or_1479_nl : STD_LOGIC;
  SIGNAL mux_1383_nl : STD_LOGIC;
  SIGNAL mux_1382_nl : STD_LOGIC;
  SIGNAL or_1478_nl : STD_LOGIC;
  SIGNAL mux_1381_nl : STD_LOGIC;
  SIGNAL or_1476_nl : STD_LOGIC;
  SIGNAL or_1475_nl : STD_LOGIC;
  SIGNAL mux_1380_nl : STD_LOGIC;
  SIGNAL mux_1379_nl : STD_LOGIC;
  SIGNAL mux_1378_nl : STD_LOGIC;
  SIGNAL or_1474_nl : STD_LOGIC;
  SIGNAL or_1472_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL or_1470_nl : STD_LOGIC;
  SIGNAL or_1469_nl : STD_LOGIC;
  SIGNAL nand_53_nl : STD_LOGIC;
  SIGNAL mux_1376_nl : STD_LOGIC;
  SIGNAL nor_1204_nl : STD_LOGIC;
  SIGNAL nor_1205_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL nand_449_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL nor_1195_nl : STD_LOGIC;
  SIGNAL nor_1196_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL nor_1197_nl : STD_LOGIC;
  SIGNAL nor_1198_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL nor_1199_nl : STD_LOGIC;
  SIGNAL nor_1200_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL nor_1201_nl : STD_LOGIC;
  SIGNAL nor_1202_nl : STD_LOGIC;
  SIGNAL or_4122_nl : STD_LOGIC;
  SIGNAL mux_1397_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL or_1495_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL or_1492_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL or_1489_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL or_1486_nl : STD_LOGIC;
  SIGNAL mux_1420_nl : STD_LOGIC;
  SIGNAL mux_1419_nl : STD_LOGIC;
  SIGNAL or_1529_nl : STD_LOGIC;
  SIGNAL mux_1418_nl : STD_LOGIC;
  SIGNAL or_1528_nl : STD_LOGIC;
  SIGNAL or_1527_nl : STD_LOGIC;
  SIGNAL mux_1417_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL or_1525_nl : STD_LOGIC;
  SIGNAL mux_1414_nl : STD_LOGIC;
  SIGNAL or_1523_nl : STD_LOGIC;
  SIGNAL mux_1413_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL or_1522_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL or_1520_nl : STD_LOGIC;
  SIGNAL or_1519_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL or_1518_nl : STD_LOGIC;
  SIGNAL or_1516_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL or_1514_nl : STD_LOGIC;
  SIGNAL or_1513_nl : STD_LOGIC;
  SIGNAL nand_55_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL nor_1193_nl : STD_LOGIC;
  SIGNAL nor_1194_nl : STD_LOGIC;
  SIGNAL mux_1435_nl : STD_LOGIC;
  SIGNAL nand_448_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL nor_1184_nl : STD_LOGIC;
  SIGNAL nor_1185_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL nor_1186_nl : STD_LOGIC;
  SIGNAL nor_1187_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL nor_1188_nl : STD_LOGIC;
  SIGNAL nor_1189_nl : STD_LOGIC;
  SIGNAL mux_1428_nl : STD_LOGIC;
  SIGNAL nor_1190_nl : STD_LOGIC;
  SIGNAL nor_1191_nl : STD_LOGIC;
  SIGNAL or_4121_nl : STD_LOGIC;
  SIGNAL mux_1427_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL mux_1425_nl : STD_LOGIC;
  SIGNAL or_1539_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL or_1536_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL or_1533_nl : STD_LOGIC;
  SIGNAL mux_1421_nl : STD_LOGIC;
  SIGNAL or_1530_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL or_1573_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL or_1572_nl : STD_LOGIC;
  SIGNAL or_1571_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL or_1569_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL or_1567_nl : STD_LOGIC;
  SIGNAL mux_1443_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL or_1566_nl : STD_LOGIC;
  SIGNAL mux_1441_nl : STD_LOGIC;
  SIGNAL or_1564_nl : STD_LOGIC;
  SIGNAL or_1563_nl : STD_LOGIC;
  SIGNAL mux_1440_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL or_1562_nl : STD_LOGIC;
  SIGNAL or_1560_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL or_1558_nl : STD_LOGIC;
  SIGNAL or_1557_nl : STD_LOGIC;
  SIGNAL nand_57_nl : STD_LOGIC;
  SIGNAL mux_1436_nl : STD_LOGIC;
  SIGNAL nor_1182_nl : STD_LOGIC;
  SIGNAL nor_1183_nl : STD_LOGIC;
  SIGNAL mux_1465_nl : STD_LOGIC;
  SIGNAL nand_447_nl : STD_LOGIC;
  SIGNAL mux_1464_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL nor_1173_nl : STD_LOGIC;
  SIGNAL nor_1174_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL nor_1175_nl : STD_LOGIC;
  SIGNAL nor_1176_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL mux_1459_nl : STD_LOGIC;
  SIGNAL nor_1177_nl : STD_LOGIC;
  SIGNAL nor_1178_nl : STD_LOGIC;
  SIGNAL mux_1458_nl : STD_LOGIC;
  SIGNAL nor_1179_nl : STD_LOGIC;
  SIGNAL nor_1180_nl : STD_LOGIC;
  SIGNAL or_4120_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL or_1583_nl : STD_LOGIC;
  SIGNAL mux_1454_nl : STD_LOGIC;
  SIGNAL or_1580_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL or_1577_nl : STD_LOGIC;
  SIGNAL mux_1451_nl : STD_LOGIC;
  SIGNAL or_1574_nl : STD_LOGIC;
  SIGNAL mux_1480_nl : STD_LOGIC;
  SIGNAL mux_1479_nl : STD_LOGIC;
  SIGNAL or_1617_nl : STD_LOGIC;
  SIGNAL mux_1478_nl : STD_LOGIC;
  SIGNAL or_1616_nl : STD_LOGIC;
  SIGNAL or_1615_nl : STD_LOGIC;
  SIGNAL mux_1477_nl : STD_LOGIC;
  SIGNAL mux_1476_nl : STD_LOGIC;
  SIGNAL mux_1475_nl : STD_LOGIC;
  SIGNAL or_1613_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL or_1611_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL or_1610_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL or_1608_nl : STD_LOGIC;
  SIGNAL or_1607_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL mux_1469_nl : STD_LOGIC;
  SIGNAL mux_1468_nl : STD_LOGIC;
  SIGNAL or_1606_nl : STD_LOGIC;
  SIGNAL or_1604_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL or_1602_nl : STD_LOGIC;
  SIGNAL or_1601_nl : STD_LOGIC;
  SIGNAL nand_59_nl : STD_LOGIC;
  SIGNAL mux_1466_nl : STD_LOGIC;
  SIGNAL nor_1171_nl : STD_LOGIC;
  SIGNAL nor_1172_nl : STD_LOGIC;
  SIGNAL mux_1495_nl : STD_LOGIC;
  SIGNAL nand_446_nl : STD_LOGIC;
  SIGNAL mux_1494_nl : STD_LOGIC;
  SIGNAL mux_1493_nl : STD_LOGIC;
  SIGNAL mux_1492_nl : STD_LOGIC;
  SIGNAL nor_1162_nl : STD_LOGIC;
  SIGNAL nor_1163_nl : STD_LOGIC;
  SIGNAL mux_1491_nl : STD_LOGIC;
  SIGNAL nor_1164_nl : STD_LOGIC;
  SIGNAL nor_1165_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL mux_1489_nl : STD_LOGIC;
  SIGNAL nor_1166_nl : STD_LOGIC;
  SIGNAL nor_1167_nl : STD_LOGIC;
  SIGNAL mux_1488_nl : STD_LOGIC;
  SIGNAL nor_1168_nl : STD_LOGIC;
  SIGNAL nor_1169_nl : STD_LOGIC;
  SIGNAL or_4119_nl : STD_LOGIC;
  SIGNAL mux_1487_nl : STD_LOGIC;
  SIGNAL mux_1486_nl : STD_LOGIC;
  SIGNAL mux_1485_nl : STD_LOGIC;
  SIGNAL nand_326_nl : STD_LOGIC;
  SIGNAL mux_1484_nl : STD_LOGIC;
  SIGNAL or_1624_nl : STD_LOGIC;
  SIGNAL mux_1483_nl : STD_LOGIC;
  SIGNAL mux_1482_nl : STD_LOGIC;
  SIGNAL or_1621_nl : STD_LOGIC;
  SIGNAL mux_1481_nl : STD_LOGIC;
  SIGNAL or_1618_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL or_1661_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL or_1660_nl : STD_LOGIC;
  SIGNAL or_1659_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL mux_1506_nl : STD_LOGIC;
  SIGNAL mux_1505_nl : STD_LOGIC;
  SIGNAL nand_325_nl : STD_LOGIC;
  SIGNAL mux_1504_nl : STD_LOGIC;
  SIGNAL or_1655_nl : STD_LOGIC;
  SIGNAL mux_1503_nl : STD_LOGIC;
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL or_1654_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL or_1652_nl : STD_LOGIC;
  SIGNAL or_1651_nl : STD_LOGIC;
  SIGNAL mux_1500_nl : STD_LOGIC;
  SIGNAL mux_1499_nl : STD_LOGIC;
  SIGNAL mux_1498_nl : STD_LOGIC;
  SIGNAL or_1650_nl : STD_LOGIC;
  SIGNAL or_1648_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL or_1646_nl : STD_LOGIC;
  SIGNAL or_1645_nl : STD_LOGIC;
  SIGNAL nand_61_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL nor_1160_nl : STD_LOGIC;
  SIGNAL nor_1161_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL nand_445_nl : STD_LOGIC;
  SIGNAL mux_1524_nl : STD_LOGIC;
  SIGNAL mux_1523_nl : STD_LOGIC;
  SIGNAL mux_1522_nl : STD_LOGIC;
  SIGNAL nor_1151_nl : STD_LOGIC;
  SIGNAL nor_1152_nl : STD_LOGIC;
  SIGNAL mux_1521_nl : STD_LOGIC;
  SIGNAL nor_1153_nl : STD_LOGIC;
  SIGNAL nor_1154_nl : STD_LOGIC;
  SIGNAL mux_1520_nl : STD_LOGIC;
  SIGNAL mux_1519_nl : STD_LOGIC;
  SIGNAL nor_1155_nl : STD_LOGIC;
  SIGNAL nor_1156_nl : STD_LOGIC;
  SIGNAL mux_1518_nl : STD_LOGIC;
  SIGNAL nor_1157_nl : STD_LOGIC;
  SIGNAL nor_1158_nl : STD_LOGIC;
  SIGNAL or_4118_nl : STD_LOGIC;
  SIGNAL mux_1517_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL mux_1515_nl : STD_LOGIC;
  SIGNAL or_1671_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL or_1668_nl : STD_LOGIC;
  SIGNAL mux_1513_nl : STD_LOGIC;
  SIGNAL mux_1512_nl : STD_LOGIC;
  SIGNAL or_1665_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL or_1662_nl : STD_LOGIC;
  SIGNAL mux_1540_nl : STD_LOGIC;
  SIGNAL mux_1539_nl : STD_LOGIC;
  SIGNAL or_1705_nl : STD_LOGIC;
  SIGNAL mux_1538_nl : STD_LOGIC;
  SIGNAL or_1704_nl : STD_LOGIC;
  SIGNAL or_1703_nl : STD_LOGIC;
  SIGNAL mux_1537_nl : STD_LOGIC;
  SIGNAL mux_1536_nl : STD_LOGIC;
  SIGNAL mux_1535_nl : STD_LOGIC;
  SIGNAL or_1701_nl : STD_LOGIC;
  SIGNAL mux_1534_nl : STD_LOGIC;
  SIGNAL or_1699_nl : STD_LOGIC;
  SIGNAL mux_1533_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL or_1698_nl : STD_LOGIC;
  SIGNAL mux_1531_nl : STD_LOGIC;
  SIGNAL or_1696_nl : STD_LOGIC;
  SIGNAL or_1695_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL mux_1529_nl : STD_LOGIC;
  SIGNAL mux_1528_nl : STD_LOGIC;
  SIGNAL or_1694_nl : STD_LOGIC;
  SIGNAL or_1692_nl : STD_LOGIC;
  SIGNAL mux_1527_nl : STD_LOGIC;
  SIGNAL or_1690_nl : STD_LOGIC;
  SIGNAL or_1689_nl : STD_LOGIC;
  SIGNAL nand_63_nl : STD_LOGIC;
  SIGNAL mux_1526_nl : STD_LOGIC;
  SIGNAL nor_1149_nl : STD_LOGIC;
  SIGNAL nor_1150_nl : STD_LOGIC;
  SIGNAL mux_1555_nl : STD_LOGIC;
  SIGNAL nand_444_nl : STD_LOGIC;
  SIGNAL mux_1554_nl : STD_LOGIC;
  SIGNAL mux_1553_nl : STD_LOGIC;
  SIGNAL mux_1552_nl : STD_LOGIC;
  SIGNAL nor_1140_nl : STD_LOGIC;
  SIGNAL nor_1141_nl : STD_LOGIC;
  SIGNAL mux_1551_nl : STD_LOGIC;
  SIGNAL nor_1142_nl : STD_LOGIC;
  SIGNAL nor_1143_nl : STD_LOGIC;
  SIGNAL mux_1550_nl : STD_LOGIC;
  SIGNAL mux_1549_nl : STD_LOGIC;
  SIGNAL nor_1144_nl : STD_LOGIC;
  SIGNAL nor_1145_nl : STD_LOGIC;
  SIGNAL mux_1548_nl : STD_LOGIC;
  SIGNAL nor_1146_nl : STD_LOGIC;
  SIGNAL nor_1147_nl : STD_LOGIC;
  SIGNAL or_4117_nl : STD_LOGIC;
  SIGNAL mux_1547_nl : STD_LOGIC;
  SIGNAL mux_1546_nl : STD_LOGIC;
  SIGNAL mux_1545_nl : STD_LOGIC;
  SIGNAL or_1715_nl : STD_LOGIC;
  SIGNAL mux_1544_nl : STD_LOGIC;
  SIGNAL or_1712_nl : STD_LOGIC;
  SIGNAL mux_1543_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL or_1709_nl : STD_LOGIC;
  SIGNAL mux_1541_nl : STD_LOGIC;
  SIGNAL or_1706_nl : STD_LOGIC;
  SIGNAL mux_1570_nl : STD_LOGIC;
  SIGNAL mux_1569_nl : STD_LOGIC;
  SIGNAL or_1749_nl : STD_LOGIC;
  SIGNAL mux_1568_nl : STD_LOGIC;
  SIGNAL or_1748_nl : STD_LOGIC;
  SIGNAL or_1747_nl : STD_LOGIC;
  SIGNAL mux_1567_nl : STD_LOGIC;
  SIGNAL mux_1566_nl : STD_LOGIC;
  SIGNAL mux_1565_nl : STD_LOGIC;
  SIGNAL or_1745_nl : STD_LOGIC;
  SIGNAL mux_1564_nl : STD_LOGIC;
  SIGNAL or_1743_nl : STD_LOGIC;
  SIGNAL mux_1563_nl : STD_LOGIC;
  SIGNAL mux_1562_nl : STD_LOGIC;
  SIGNAL or_1742_nl : STD_LOGIC;
  SIGNAL mux_1561_nl : STD_LOGIC;
  SIGNAL or_1740_nl : STD_LOGIC;
  SIGNAL or_1739_nl : STD_LOGIC;
  SIGNAL mux_1560_nl : STD_LOGIC;
  SIGNAL mux_1559_nl : STD_LOGIC;
  SIGNAL mux_1558_nl : STD_LOGIC;
  SIGNAL or_1738_nl : STD_LOGIC;
  SIGNAL or_1736_nl : STD_LOGIC;
  SIGNAL mux_1557_nl : STD_LOGIC;
  SIGNAL or_1734_nl : STD_LOGIC;
  SIGNAL or_1733_nl : STD_LOGIC;
  SIGNAL nand_65_nl : STD_LOGIC;
  SIGNAL mux_1556_nl : STD_LOGIC;
  SIGNAL nor_1138_nl : STD_LOGIC;
  SIGNAL nor_1139_nl : STD_LOGIC;
  SIGNAL mux_1585_nl : STD_LOGIC;
  SIGNAL nand_443_nl : STD_LOGIC;
  SIGNAL mux_1584_nl : STD_LOGIC;
  SIGNAL mux_1583_nl : STD_LOGIC;
  SIGNAL mux_1582_nl : STD_LOGIC;
  SIGNAL nor_1129_nl : STD_LOGIC;
  SIGNAL nor_1130_nl : STD_LOGIC;
  SIGNAL mux_1581_nl : STD_LOGIC;
  SIGNAL nor_1131_nl : STD_LOGIC;
  SIGNAL nor_1132_nl : STD_LOGIC;
  SIGNAL mux_1580_nl : STD_LOGIC;
  SIGNAL mux_1579_nl : STD_LOGIC;
  SIGNAL nor_1133_nl : STD_LOGIC;
  SIGNAL nor_1134_nl : STD_LOGIC;
  SIGNAL mux_1578_nl : STD_LOGIC;
  SIGNAL nor_1135_nl : STD_LOGIC;
  SIGNAL nor_1136_nl : STD_LOGIC;
  SIGNAL or_4116_nl : STD_LOGIC;
  SIGNAL mux_1577_nl : STD_LOGIC;
  SIGNAL mux_1576_nl : STD_LOGIC;
  SIGNAL mux_1575_nl : STD_LOGIC;
  SIGNAL or_1759_nl : STD_LOGIC;
  SIGNAL mux_1574_nl : STD_LOGIC;
  SIGNAL or_1756_nl : STD_LOGIC;
  SIGNAL mux_1573_nl : STD_LOGIC;
  SIGNAL mux_1572_nl : STD_LOGIC;
  SIGNAL or_1753_nl : STD_LOGIC;
  SIGNAL mux_1571_nl : STD_LOGIC;
  SIGNAL or_1750_nl : STD_LOGIC;
  SIGNAL mux_1600_nl : STD_LOGIC;
  SIGNAL mux_1599_nl : STD_LOGIC;
  SIGNAL or_1793_nl : STD_LOGIC;
  SIGNAL mux_1598_nl : STD_LOGIC;
  SIGNAL or_1792_nl : STD_LOGIC;
  SIGNAL or_1791_nl : STD_LOGIC;
  SIGNAL mux_1597_nl : STD_LOGIC;
  SIGNAL mux_1596_nl : STD_LOGIC;
  SIGNAL mux_1595_nl : STD_LOGIC;
  SIGNAL or_1789_nl : STD_LOGIC;
  SIGNAL mux_1594_nl : STD_LOGIC;
  SIGNAL or_1787_nl : STD_LOGIC;
  SIGNAL mux_1593_nl : STD_LOGIC;
  SIGNAL mux_1592_nl : STD_LOGIC;
  SIGNAL or_1786_nl : STD_LOGIC;
  SIGNAL mux_1591_nl : STD_LOGIC;
  SIGNAL or_1784_nl : STD_LOGIC;
  SIGNAL or_1783_nl : STD_LOGIC;
  SIGNAL mux_1590_nl : STD_LOGIC;
  SIGNAL mux_1589_nl : STD_LOGIC;
  SIGNAL mux_1588_nl : STD_LOGIC;
  SIGNAL or_1782_nl : STD_LOGIC;
  SIGNAL or_1780_nl : STD_LOGIC;
  SIGNAL mux_1587_nl : STD_LOGIC;
  SIGNAL or_1778_nl : STD_LOGIC;
  SIGNAL or_1777_nl : STD_LOGIC;
  SIGNAL nand_67_nl : STD_LOGIC;
  SIGNAL mux_1586_nl : STD_LOGIC;
  SIGNAL nor_1127_nl : STD_LOGIC;
  SIGNAL nor_1128_nl : STD_LOGIC;
  SIGNAL mux_1615_nl : STD_LOGIC;
  SIGNAL nand_442_nl : STD_LOGIC;
  SIGNAL mux_1614_nl : STD_LOGIC;
  SIGNAL mux_1613_nl : STD_LOGIC;
  SIGNAL mux_1612_nl : STD_LOGIC;
  SIGNAL nor_1118_nl : STD_LOGIC;
  SIGNAL nor_1119_nl : STD_LOGIC;
  SIGNAL mux_1611_nl : STD_LOGIC;
  SIGNAL nor_1120_nl : STD_LOGIC;
  SIGNAL nor_1121_nl : STD_LOGIC;
  SIGNAL mux_1610_nl : STD_LOGIC;
  SIGNAL mux_1609_nl : STD_LOGIC;
  SIGNAL nor_1122_nl : STD_LOGIC;
  SIGNAL nor_1123_nl : STD_LOGIC;
  SIGNAL mux_1608_nl : STD_LOGIC;
  SIGNAL nor_1124_nl : STD_LOGIC;
  SIGNAL nor_1125_nl : STD_LOGIC;
  SIGNAL or_4115_nl : STD_LOGIC;
  SIGNAL mux_1607_nl : STD_LOGIC;
  SIGNAL mux_1606_nl : STD_LOGIC;
  SIGNAL mux_1605_nl : STD_LOGIC;
  SIGNAL nand_324_nl : STD_LOGIC;
  SIGNAL mux_1604_nl : STD_LOGIC;
  SIGNAL or_1800_nl : STD_LOGIC;
  SIGNAL mux_1603_nl : STD_LOGIC;
  SIGNAL mux_1602_nl : STD_LOGIC;
  SIGNAL or_1797_nl : STD_LOGIC;
  SIGNAL mux_1601_nl : STD_LOGIC;
  SIGNAL or_1794_nl : STD_LOGIC;
  SIGNAL mux_1630_nl : STD_LOGIC;
  SIGNAL mux_1629_nl : STD_LOGIC;
  SIGNAL or_1837_nl : STD_LOGIC;
  SIGNAL mux_1628_nl : STD_LOGIC;
  SIGNAL or_1836_nl : STD_LOGIC;
  SIGNAL or_1835_nl : STD_LOGIC;
  SIGNAL mux_1627_nl : STD_LOGIC;
  SIGNAL mux_1626_nl : STD_LOGIC;
  SIGNAL mux_1625_nl : STD_LOGIC;
  SIGNAL nand_323_nl : STD_LOGIC;
  SIGNAL mux_1624_nl : STD_LOGIC;
  SIGNAL or_1831_nl : STD_LOGIC;
  SIGNAL mux_1623_nl : STD_LOGIC;
  SIGNAL mux_1622_nl : STD_LOGIC;
  SIGNAL or_1830_nl : STD_LOGIC;
  SIGNAL mux_1621_nl : STD_LOGIC;
  SIGNAL or_1828_nl : STD_LOGIC;
  SIGNAL or_1827_nl : STD_LOGIC;
  SIGNAL mux_1620_nl : STD_LOGIC;
  SIGNAL mux_1619_nl : STD_LOGIC;
  SIGNAL mux_1618_nl : STD_LOGIC;
  SIGNAL or_1826_nl : STD_LOGIC;
  SIGNAL or_1824_nl : STD_LOGIC;
  SIGNAL mux_1617_nl : STD_LOGIC;
  SIGNAL or_1822_nl : STD_LOGIC;
  SIGNAL or_1821_nl : STD_LOGIC;
  SIGNAL nand_69_nl : STD_LOGIC;
  SIGNAL mux_1616_nl : STD_LOGIC;
  SIGNAL nor_1116_nl : STD_LOGIC;
  SIGNAL nor_1117_nl : STD_LOGIC;
  SIGNAL mux_1645_nl : STD_LOGIC;
  SIGNAL nand_441_nl : STD_LOGIC;
  SIGNAL mux_1644_nl : STD_LOGIC;
  SIGNAL mux_1643_nl : STD_LOGIC;
  SIGNAL mux_1642_nl : STD_LOGIC;
  SIGNAL nor_1107_nl : STD_LOGIC;
  SIGNAL nor_1108_nl : STD_LOGIC;
  SIGNAL mux_1641_nl : STD_LOGIC;
  SIGNAL nor_1109_nl : STD_LOGIC;
  SIGNAL nor_1110_nl : STD_LOGIC;
  SIGNAL mux_1640_nl : STD_LOGIC;
  SIGNAL mux_1639_nl : STD_LOGIC;
  SIGNAL nor_1111_nl : STD_LOGIC;
  SIGNAL nor_1112_nl : STD_LOGIC;
  SIGNAL mux_1638_nl : STD_LOGIC;
  SIGNAL nor_1113_nl : STD_LOGIC;
  SIGNAL nor_1114_nl : STD_LOGIC;
  SIGNAL or_4114_nl : STD_LOGIC;
  SIGNAL mux_1637_nl : STD_LOGIC;
  SIGNAL mux_1636_nl : STD_LOGIC;
  SIGNAL mux_1635_nl : STD_LOGIC;
  SIGNAL or_1847_nl : STD_LOGIC;
  SIGNAL mux_1634_nl : STD_LOGIC;
  SIGNAL or_1844_nl : STD_LOGIC;
  SIGNAL mux_1633_nl : STD_LOGIC;
  SIGNAL mux_1632_nl : STD_LOGIC;
  SIGNAL or_1841_nl : STD_LOGIC;
  SIGNAL mux_1631_nl : STD_LOGIC;
  SIGNAL or_1838_nl : STD_LOGIC;
  SIGNAL mux_1660_nl : STD_LOGIC;
  SIGNAL mux_1659_nl : STD_LOGIC;
  SIGNAL or_1881_nl : STD_LOGIC;
  SIGNAL mux_1658_nl : STD_LOGIC;
  SIGNAL or_1880_nl : STD_LOGIC;
  SIGNAL or_1879_nl : STD_LOGIC;
  SIGNAL mux_1657_nl : STD_LOGIC;
  SIGNAL mux_1656_nl : STD_LOGIC;
  SIGNAL mux_1655_nl : STD_LOGIC;
  SIGNAL or_1877_nl : STD_LOGIC;
  SIGNAL mux_1654_nl : STD_LOGIC;
  SIGNAL or_1875_nl : STD_LOGIC;
  SIGNAL mux_1653_nl : STD_LOGIC;
  SIGNAL mux_1652_nl : STD_LOGIC;
  SIGNAL or_1874_nl : STD_LOGIC;
  SIGNAL mux_1651_nl : STD_LOGIC;
  SIGNAL or_1872_nl : STD_LOGIC;
  SIGNAL or_1871_nl : STD_LOGIC;
  SIGNAL mux_1650_nl : STD_LOGIC;
  SIGNAL mux_1649_nl : STD_LOGIC;
  SIGNAL mux_1648_nl : STD_LOGIC;
  SIGNAL or_1870_nl : STD_LOGIC;
  SIGNAL or_1868_nl : STD_LOGIC;
  SIGNAL mux_1647_nl : STD_LOGIC;
  SIGNAL or_1866_nl : STD_LOGIC;
  SIGNAL or_1865_nl : STD_LOGIC;
  SIGNAL nand_71_nl : STD_LOGIC;
  SIGNAL mux_1646_nl : STD_LOGIC;
  SIGNAL nor_1105_nl : STD_LOGIC;
  SIGNAL nor_1106_nl : STD_LOGIC;
  SIGNAL mux_1675_nl : STD_LOGIC;
  SIGNAL nand_440_nl : STD_LOGIC;
  SIGNAL mux_1674_nl : STD_LOGIC;
  SIGNAL mux_1673_nl : STD_LOGIC;
  SIGNAL mux_1672_nl : STD_LOGIC;
  SIGNAL nor_1096_nl : STD_LOGIC;
  SIGNAL nor_1097_nl : STD_LOGIC;
  SIGNAL mux_1671_nl : STD_LOGIC;
  SIGNAL nor_1098_nl : STD_LOGIC;
  SIGNAL nor_1099_nl : STD_LOGIC;
  SIGNAL mux_1670_nl : STD_LOGIC;
  SIGNAL mux_1669_nl : STD_LOGIC;
  SIGNAL nor_1100_nl : STD_LOGIC;
  SIGNAL nor_1101_nl : STD_LOGIC;
  SIGNAL mux_1668_nl : STD_LOGIC;
  SIGNAL nor_1102_nl : STD_LOGIC;
  SIGNAL nor_1103_nl : STD_LOGIC;
  SIGNAL or_4113_nl : STD_LOGIC;
  SIGNAL mux_1667_nl : STD_LOGIC;
  SIGNAL mux_1666_nl : STD_LOGIC;
  SIGNAL mux_1665_nl : STD_LOGIC;
  SIGNAL nand_322_nl : STD_LOGIC;
  SIGNAL mux_1664_nl : STD_LOGIC;
  SIGNAL or_1888_nl : STD_LOGIC;
  SIGNAL mux_1663_nl : STD_LOGIC;
  SIGNAL mux_1662_nl : STD_LOGIC;
  SIGNAL or_1885_nl : STD_LOGIC;
  SIGNAL mux_1661_nl : STD_LOGIC;
  SIGNAL or_1882_nl : STD_LOGIC;
  SIGNAL mux_1690_nl : STD_LOGIC;
  SIGNAL mux_1689_nl : STD_LOGIC;
  SIGNAL or_1925_nl : STD_LOGIC;
  SIGNAL mux_1688_nl : STD_LOGIC;
  SIGNAL or_1924_nl : STD_LOGIC;
  SIGNAL or_1923_nl : STD_LOGIC;
  SIGNAL mux_1687_nl : STD_LOGIC;
  SIGNAL mux_1686_nl : STD_LOGIC;
  SIGNAL mux_1685_nl : STD_LOGIC;
  SIGNAL nand_321_nl : STD_LOGIC;
  SIGNAL mux_1684_nl : STD_LOGIC;
  SIGNAL or_1919_nl : STD_LOGIC;
  SIGNAL mux_1683_nl : STD_LOGIC;
  SIGNAL mux_1682_nl : STD_LOGIC;
  SIGNAL or_1918_nl : STD_LOGIC;
  SIGNAL mux_1681_nl : STD_LOGIC;
  SIGNAL or_1916_nl : STD_LOGIC;
  SIGNAL or_1915_nl : STD_LOGIC;
  SIGNAL mux_1680_nl : STD_LOGIC;
  SIGNAL mux_1679_nl : STD_LOGIC;
  SIGNAL mux_1678_nl : STD_LOGIC;
  SIGNAL or_1914_nl : STD_LOGIC;
  SIGNAL or_1912_nl : STD_LOGIC;
  SIGNAL mux_1677_nl : STD_LOGIC;
  SIGNAL or_1910_nl : STD_LOGIC;
  SIGNAL or_1909_nl : STD_LOGIC;
  SIGNAL nand_73_nl : STD_LOGIC;
  SIGNAL mux_1676_nl : STD_LOGIC;
  SIGNAL nor_1094_nl : STD_LOGIC;
  SIGNAL nor_1095_nl : STD_LOGIC;
  SIGNAL mux_1705_nl : STD_LOGIC;
  SIGNAL nand_439_nl : STD_LOGIC;
  SIGNAL mux_1704_nl : STD_LOGIC;
  SIGNAL mux_1703_nl : STD_LOGIC;
  SIGNAL mux_1702_nl : STD_LOGIC;
  SIGNAL nor_1086_nl : STD_LOGIC;
  SIGNAL and_602_nl : STD_LOGIC;
  SIGNAL mux_1701_nl : STD_LOGIC;
  SIGNAL nor_1087_nl : STD_LOGIC;
  SIGNAL nor_1088_nl : STD_LOGIC;
  SIGNAL mux_1700_nl : STD_LOGIC;
  SIGNAL mux_1699_nl : STD_LOGIC;
  SIGNAL nor_1089_nl : STD_LOGIC;
  SIGNAL nor_1090_nl : STD_LOGIC;
  SIGNAL mux_1698_nl : STD_LOGIC;
  SIGNAL nor_1091_nl : STD_LOGIC;
  SIGNAL nor_1092_nl : STD_LOGIC;
  SIGNAL or_4112_nl : STD_LOGIC;
  SIGNAL mux_1697_nl : STD_LOGIC;
  SIGNAL mux_1696_nl : STD_LOGIC;
  SIGNAL mux_1695_nl : STD_LOGIC;
  SIGNAL nand_320_nl : STD_LOGIC;
  SIGNAL mux_1694_nl : STD_LOGIC;
  SIGNAL or_1932_nl : STD_LOGIC;
  SIGNAL mux_1693_nl : STD_LOGIC;
  SIGNAL mux_1692_nl : STD_LOGIC;
  SIGNAL or_1929_nl : STD_LOGIC;
  SIGNAL mux_1691_nl : STD_LOGIC;
  SIGNAL or_1926_nl : STD_LOGIC;
  SIGNAL mux_1720_nl : STD_LOGIC;
  SIGNAL mux_1719_nl : STD_LOGIC;
  SIGNAL or_1969_nl : STD_LOGIC;
  SIGNAL mux_1718_nl : STD_LOGIC;
  SIGNAL or_1968_nl : STD_LOGIC;
  SIGNAL or_1967_nl : STD_LOGIC;
  SIGNAL mux_1717_nl : STD_LOGIC;
  SIGNAL mux_1716_nl : STD_LOGIC;
  SIGNAL mux_1715_nl : STD_LOGIC;
  SIGNAL nand_318_nl : STD_LOGIC;
  SIGNAL mux_1714_nl : STD_LOGIC;
  SIGNAL or_1963_nl : STD_LOGIC;
  SIGNAL mux_1713_nl : STD_LOGIC;
  SIGNAL mux_1712_nl : STD_LOGIC;
  SIGNAL or_1962_nl : STD_LOGIC;
  SIGNAL mux_1711_nl : STD_LOGIC;
  SIGNAL or_1960_nl : STD_LOGIC;
  SIGNAL or_1959_nl : STD_LOGIC;
  SIGNAL mux_1710_nl : STD_LOGIC;
  SIGNAL mux_1709_nl : STD_LOGIC;
  SIGNAL mux_1708_nl : STD_LOGIC;
  SIGNAL nand_319_nl : STD_LOGIC;
  SIGNAL or_1956_nl : STD_LOGIC;
  SIGNAL mux_1707_nl : STD_LOGIC;
  SIGNAL or_1954_nl : STD_LOGIC;
  SIGNAL or_1953_nl : STD_LOGIC;
  SIGNAL nand_75_nl : STD_LOGIC;
  SIGNAL mux_1706_nl : STD_LOGIC;
  SIGNAL nor_1084_nl : STD_LOGIC;
  SIGNAL nor_1085_nl : STD_LOGIC;
  SIGNAL mux_1735_nl : STD_LOGIC;
  SIGNAL nand_438_nl : STD_LOGIC;
  SIGNAL mux_1734_nl : STD_LOGIC;
  SIGNAL mux_1733_nl : STD_LOGIC;
  SIGNAL mux_1732_nl : STD_LOGIC;
  SIGNAL nor_1077_nl : STD_LOGIC;
  SIGNAL nor_1078_nl : STD_LOGIC;
  SIGNAL mux_1731_nl : STD_LOGIC;
  SIGNAL and_599_nl : STD_LOGIC;
  SIGNAL and_600_nl : STD_LOGIC;
  SIGNAL mux_1730_nl : STD_LOGIC;
  SIGNAL mux_1729_nl : STD_LOGIC;
  SIGNAL and_811_nl : STD_LOGIC;
  SIGNAL and_818_nl : STD_LOGIC;
  SIGNAL mux_1728_nl : STD_LOGIC;
  SIGNAL nor_1081_nl : STD_LOGIC;
  SIGNAL nor_1082_nl : STD_LOGIC;
  SIGNAL or_4111_nl : STD_LOGIC;
  SIGNAL mux_1727_nl : STD_LOGIC;
  SIGNAL mux_1726_nl : STD_LOGIC;
  SIGNAL mux_1725_nl : STD_LOGIC;
  SIGNAL nand_313_nl : STD_LOGIC;
  SIGNAL mux_1724_nl : STD_LOGIC;
  SIGNAL nand_314_nl : STD_LOGIC;
  SIGNAL mux_1723_nl : STD_LOGIC;
  SIGNAL mux_1722_nl : STD_LOGIC;
  SIGNAL nand_478_nl : STD_LOGIC;
  SIGNAL mux_1721_nl : STD_LOGIC;
  SIGNAL or_1970_nl : STD_LOGIC;
  SIGNAL mux_1750_nl : STD_LOGIC;
  SIGNAL mux_1749_nl : STD_LOGIC;
  SIGNAL or_2012_nl : STD_LOGIC;
  SIGNAL mux_1748_nl : STD_LOGIC;
  SIGNAL or_2011_nl : STD_LOGIC;
  SIGNAL or_2010_nl : STD_LOGIC;
  SIGNAL mux_1747_nl : STD_LOGIC;
  SIGNAL mux_1746_nl : STD_LOGIC;
  SIGNAL mux_1745_nl : STD_LOGIC;
  SIGNAL nand_302_nl : STD_LOGIC;
  SIGNAL mux_1744_nl : STD_LOGIC;
  SIGNAL nand_303_nl : STD_LOGIC;
  SIGNAL mux_1743_nl : STD_LOGIC;
  SIGNAL mux_1742_nl : STD_LOGIC;
  SIGNAL nand_404_nl : STD_LOGIC;
  SIGNAL mux_1741_nl : STD_LOGIC;
  SIGNAL or_2003_nl : STD_LOGIC;
  SIGNAL or_2002_nl : STD_LOGIC;
  SIGNAL mux_1740_nl : STD_LOGIC;
  SIGNAL mux_1739_nl : STD_LOGIC;
  SIGNAL mux_1738_nl : STD_LOGIC;
  SIGNAL or_2001_nl : STD_LOGIC;
  SIGNAL or_1999_nl : STD_LOGIC;
  SIGNAL mux_1737_nl : STD_LOGIC;
  SIGNAL nand_307_nl : STD_LOGIC;
  SIGNAL nand_308_nl : STD_LOGIC;
  SIGNAL nand_77_nl : STD_LOGIC;
  SIGNAL mux_1736_nl : STD_LOGIC;
  SIGNAL nor_1075_nl : STD_LOGIC;
  SIGNAL nor_1076_nl : STD_LOGIC;
  SIGNAL mux_1765_nl : STD_LOGIC;
  SIGNAL nand_437_nl : STD_LOGIC;
  SIGNAL mux_1764_nl : STD_LOGIC;
  SIGNAL mux_1763_nl : STD_LOGIC;
  SIGNAL mux_1762_nl : STD_LOGIC;
  SIGNAL nor_1066_nl : STD_LOGIC;
  SIGNAL nor_1067_nl : STD_LOGIC;
  SIGNAL mux_1761_nl : STD_LOGIC;
  SIGNAL nor_1068_nl : STD_LOGIC;
  SIGNAL nor_1069_nl : STD_LOGIC;
  SIGNAL mux_1760_nl : STD_LOGIC;
  SIGNAL mux_1759_nl : STD_LOGIC;
  SIGNAL nor_1070_nl : STD_LOGIC;
  SIGNAL nor_1071_nl : STD_LOGIC;
  SIGNAL mux_1758_nl : STD_LOGIC;
  SIGNAL nor_1072_nl : STD_LOGIC;
  SIGNAL nor_1073_nl : STD_LOGIC;
  SIGNAL or_4110_nl : STD_LOGIC;
  SIGNAL mux_1757_nl : STD_LOGIC;
  SIGNAL mux_1756_nl : STD_LOGIC;
  SIGNAL mux_1755_nl : STD_LOGIC;
  SIGNAL or_2022_nl : STD_LOGIC;
  SIGNAL mux_1754_nl : STD_LOGIC;
  SIGNAL or_2019_nl : STD_LOGIC;
  SIGNAL mux_1753_nl : STD_LOGIC;
  SIGNAL mux_1752_nl : STD_LOGIC;
  SIGNAL or_2016_nl : STD_LOGIC;
  SIGNAL mux_1751_nl : STD_LOGIC;
  SIGNAL or_2013_nl : STD_LOGIC;
  SIGNAL mux_1780_nl : STD_LOGIC;
  SIGNAL mux_1779_nl : STD_LOGIC;
  SIGNAL or_2056_nl : STD_LOGIC;
  SIGNAL mux_1778_nl : STD_LOGIC;
  SIGNAL or_2055_nl : STD_LOGIC;
  SIGNAL or_2054_nl : STD_LOGIC;
  SIGNAL mux_1777_nl : STD_LOGIC;
  SIGNAL mux_1776_nl : STD_LOGIC;
  SIGNAL mux_1775_nl : STD_LOGIC;
  SIGNAL or_2052_nl : STD_LOGIC;
  SIGNAL mux_1774_nl : STD_LOGIC;
  SIGNAL or_2050_nl : STD_LOGIC;
  SIGNAL mux_1773_nl : STD_LOGIC;
  SIGNAL mux_1772_nl : STD_LOGIC;
  SIGNAL or_2049_nl : STD_LOGIC;
  SIGNAL mux_1771_nl : STD_LOGIC;
  SIGNAL or_2047_nl : STD_LOGIC;
  SIGNAL or_2046_nl : STD_LOGIC;
  SIGNAL mux_1770_nl : STD_LOGIC;
  SIGNAL mux_1769_nl : STD_LOGIC;
  SIGNAL mux_1768_nl : STD_LOGIC;
  SIGNAL or_2045_nl : STD_LOGIC;
  SIGNAL or_2043_nl : STD_LOGIC;
  SIGNAL mux_1767_nl : STD_LOGIC;
  SIGNAL or_2041_nl : STD_LOGIC;
  SIGNAL or_2040_nl : STD_LOGIC;
  SIGNAL nand_79_nl : STD_LOGIC;
  SIGNAL mux_1766_nl : STD_LOGIC;
  SIGNAL nor_1064_nl : STD_LOGIC;
  SIGNAL nor_1065_nl : STD_LOGIC;
  SIGNAL mux_1795_nl : STD_LOGIC;
  SIGNAL nand_436_nl : STD_LOGIC;
  SIGNAL mux_1794_nl : STD_LOGIC;
  SIGNAL mux_1793_nl : STD_LOGIC;
  SIGNAL mux_1792_nl : STD_LOGIC;
  SIGNAL nor_1055_nl : STD_LOGIC;
  SIGNAL nor_1056_nl : STD_LOGIC;
  SIGNAL mux_1791_nl : STD_LOGIC;
  SIGNAL nor_1057_nl : STD_LOGIC;
  SIGNAL nor_1058_nl : STD_LOGIC;
  SIGNAL mux_1790_nl : STD_LOGIC;
  SIGNAL mux_1789_nl : STD_LOGIC;
  SIGNAL nor_1059_nl : STD_LOGIC;
  SIGNAL nor_1060_nl : STD_LOGIC;
  SIGNAL mux_1788_nl : STD_LOGIC;
  SIGNAL nor_1061_nl : STD_LOGIC;
  SIGNAL nor_1062_nl : STD_LOGIC;
  SIGNAL or_4109_nl : STD_LOGIC;
  SIGNAL mux_1787_nl : STD_LOGIC;
  SIGNAL mux_1786_nl : STD_LOGIC;
  SIGNAL mux_1785_nl : STD_LOGIC;
  SIGNAL or_2066_nl : STD_LOGIC;
  SIGNAL mux_1784_nl : STD_LOGIC;
  SIGNAL or_2063_nl : STD_LOGIC;
  SIGNAL mux_1783_nl : STD_LOGIC;
  SIGNAL mux_1782_nl : STD_LOGIC;
  SIGNAL or_2060_nl : STD_LOGIC;
  SIGNAL mux_1781_nl : STD_LOGIC;
  SIGNAL or_2057_nl : STD_LOGIC;
  SIGNAL mux_1810_nl : STD_LOGIC;
  SIGNAL mux_1809_nl : STD_LOGIC;
  SIGNAL or_2100_nl : STD_LOGIC;
  SIGNAL mux_1808_nl : STD_LOGIC;
  SIGNAL or_2099_nl : STD_LOGIC;
  SIGNAL or_2098_nl : STD_LOGIC;
  SIGNAL mux_1807_nl : STD_LOGIC;
  SIGNAL mux_1806_nl : STD_LOGIC;
  SIGNAL mux_1805_nl : STD_LOGIC;
  SIGNAL or_2096_nl : STD_LOGIC;
  SIGNAL mux_1804_nl : STD_LOGIC;
  SIGNAL or_2094_nl : STD_LOGIC;
  SIGNAL mux_1803_nl : STD_LOGIC;
  SIGNAL mux_1802_nl : STD_LOGIC;
  SIGNAL or_2093_nl : STD_LOGIC;
  SIGNAL mux_1801_nl : STD_LOGIC;
  SIGNAL or_2091_nl : STD_LOGIC;
  SIGNAL or_2090_nl : STD_LOGIC;
  SIGNAL mux_1800_nl : STD_LOGIC;
  SIGNAL mux_1799_nl : STD_LOGIC;
  SIGNAL mux_1798_nl : STD_LOGIC;
  SIGNAL or_2089_nl : STD_LOGIC;
  SIGNAL or_2087_nl : STD_LOGIC;
  SIGNAL mux_1797_nl : STD_LOGIC;
  SIGNAL or_2085_nl : STD_LOGIC;
  SIGNAL or_2084_nl : STD_LOGIC;
  SIGNAL nand_81_nl : STD_LOGIC;
  SIGNAL mux_1796_nl : STD_LOGIC;
  SIGNAL nor_1053_nl : STD_LOGIC;
  SIGNAL nor_1054_nl : STD_LOGIC;
  SIGNAL mux_1825_nl : STD_LOGIC;
  SIGNAL nand_435_nl : STD_LOGIC;
  SIGNAL mux_1824_nl : STD_LOGIC;
  SIGNAL mux_1823_nl : STD_LOGIC;
  SIGNAL mux_1822_nl : STD_LOGIC;
  SIGNAL nor_1044_nl : STD_LOGIC;
  SIGNAL nor_1045_nl : STD_LOGIC;
  SIGNAL mux_1821_nl : STD_LOGIC;
  SIGNAL nor_1046_nl : STD_LOGIC;
  SIGNAL nor_1047_nl : STD_LOGIC;
  SIGNAL mux_1820_nl : STD_LOGIC;
  SIGNAL mux_1819_nl : STD_LOGIC;
  SIGNAL nor_1048_nl : STD_LOGIC;
  SIGNAL nor_1049_nl : STD_LOGIC;
  SIGNAL mux_1818_nl : STD_LOGIC;
  SIGNAL nor_1050_nl : STD_LOGIC;
  SIGNAL nor_1051_nl : STD_LOGIC;
  SIGNAL or_4108_nl : STD_LOGIC;
  SIGNAL mux_1817_nl : STD_LOGIC;
  SIGNAL mux_1816_nl : STD_LOGIC;
  SIGNAL mux_1815_nl : STD_LOGIC;
  SIGNAL or_2110_nl : STD_LOGIC;
  SIGNAL mux_1814_nl : STD_LOGIC;
  SIGNAL or_2107_nl : STD_LOGIC;
  SIGNAL mux_1813_nl : STD_LOGIC;
  SIGNAL mux_1812_nl : STD_LOGIC;
  SIGNAL or_2104_nl : STD_LOGIC;
  SIGNAL mux_1811_nl : STD_LOGIC;
  SIGNAL or_2101_nl : STD_LOGIC;
  SIGNAL mux_1840_nl : STD_LOGIC;
  SIGNAL mux_1839_nl : STD_LOGIC;
  SIGNAL or_2144_nl : STD_LOGIC;
  SIGNAL mux_1838_nl : STD_LOGIC;
  SIGNAL or_2143_nl : STD_LOGIC;
  SIGNAL or_2142_nl : STD_LOGIC;
  SIGNAL mux_1837_nl : STD_LOGIC;
  SIGNAL mux_1836_nl : STD_LOGIC;
  SIGNAL mux_1835_nl : STD_LOGIC;
  SIGNAL or_2140_nl : STD_LOGIC;
  SIGNAL mux_1834_nl : STD_LOGIC;
  SIGNAL or_2138_nl : STD_LOGIC;
  SIGNAL mux_1833_nl : STD_LOGIC;
  SIGNAL mux_1832_nl : STD_LOGIC;
  SIGNAL or_2137_nl : STD_LOGIC;
  SIGNAL mux_1831_nl : STD_LOGIC;
  SIGNAL or_2135_nl : STD_LOGIC;
  SIGNAL or_2134_nl : STD_LOGIC;
  SIGNAL mux_1830_nl : STD_LOGIC;
  SIGNAL mux_1829_nl : STD_LOGIC;
  SIGNAL mux_1828_nl : STD_LOGIC;
  SIGNAL or_2133_nl : STD_LOGIC;
  SIGNAL or_2131_nl : STD_LOGIC;
  SIGNAL mux_1827_nl : STD_LOGIC;
  SIGNAL or_2129_nl : STD_LOGIC;
  SIGNAL or_2128_nl : STD_LOGIC;
  SIGNAL nand_83_nl : STD_LOGIC;
  SIGNAL mux_1826_nl : STD_LOGIC;
  SIGNAL nor_1042_nl : STD_LOGIC;
  SIGNAL nor_1043_nl : STD_LOGIC;
  SIGNAL mux_1855_nl : STD_LOGIC;
  SIGNAL nand_434_nl : STD_LOGIC;
  SIGNAL mux_1854_nl : STD_LOGIC;
  SIGNAL mux_1853_nl : STD_LOGIC;
  SIGNAL mux_1852_nl : STD_LOGIC;
  SIGNAL nor_1033_nl : STD_LOGIC;
  SIGNAL nor_1034_nl : STD_LOGIC;
  SIGNAL mux_1851_nl : STD_LOGIC;
  SIGNAL nor_1035_nl : STD_LOGIC;
  SIGNAL nor_1036_nl : STD_LOGIC;
  SIGNAL mux_1850_nl : STD_LOGIC;
  SIGNAL mux_1849_nl : STD_LOGIC;
  SIGNAL nor_1037_nl : STD_LOGIC;
  SIGNAL nor_1038_nl : STD_LOGIC;
  SIGNAL mux_1848_nl : STD_LOGIC;
  SIGNAL nor_1039_nl : STD_LOGIC;
  SIGNAL nor_1040_nl : STD_LOGIC;
  SIGNAL or_4107_nl : STD_LOGIC;
  SIGNAL mux_1847_nl : STD_LOGIC;
  SIGNAL mux_1846_nl : STD_LOGIC;
  SIGNAL mux_1845_nl : STD_LOGIC;
  SIGNAL or_2154_nl : STD_LOGIC;
  SIGNAL mux_1844_nl : STD_LOGIC;
  SIGNAL or_2151_nl : STD_LOGIC;
  SIGNAL mux_1843_nl : STD_LOGIC;
  SIGNAL mux_1842_nl : STD_LOGIC;
  SIGNAL or_2148_nl : STD_LOGIC;
  SIGNAL mux_1841_nl : STD_LOGIC;
  SIGNAL or_2145_nl : STD_LOGIC;
  SIGNAL mux_1870_nl : STD_LOGIC;
  SIGNAL mux_1869_nl : STD_LOGIC;
  SIGNAL or_2188_nl : STD_LOGIC;
  SIGNAL mux_1868_nl : STD_LOGIC;
  SIGNAL or_2187_nl : STD_LOGIC;
  SIGNAL or_2186_nl : STD_LOGIC;
  SIGNAL mux_1867_nl : STD_LOGIC;
  SIGNAL mux_1866_nl : STD_LOGIC;
  SIGNAL mux_1865_nl : STD_LOGIC;
  SIGNAL or_2184_nl : STD_LOGIC;
  SIGNAL mux_1864_nl : STD_LOGIC;
  SIGNAL or_2182_nl : STD_LOGIC;
  SIGNAL mux_1863_nl : STD_LOGIC;
  SIGNAL mux_1862_nl : STD_LOGIC;
  SIGNAL or_2181_nl : STD_LOGIC;
  SIGNAL mux_1861_nl : STD_LOGIC;
  SIGNAL or_2179_nl : STD_LOGIC;
  SIGNAL or_2178_nl : STD_LOGIC;
  SIGNAL mux_1860_nl : STD_LOGIC;
  SIGNAL mux_1859_nl : STD_LOGIC;
  SIGNAL mux_1858_nl : STD_LOGIC;
  SIGNAL or_2177_nl : STD_LOGIC;
  SIGNAL or_2175_nl : STD_LOGIC;
  SIGNAL mux_1857_nl : STD_LOGIC;
  SIGNAL or_2173_nl : STD_LOGIC;
  SIGNAL or_2172_nl : STD_LOGIC;
  SIGNAL nand_85_nl : STD_LOGIC;
  SIGNAL mux_1856_nl : STD_LOGIC;
  SIGNAL nor_1031_nl : STD_LOGIC;
  SIGNAL nor_1032_nl : STD_LOGIC;
  SIGNAL mux_1885_nl : STD_LOGIC;
  SIGNAL nand_433_nl : STD_LOGIC;
  SIGNAL mux_1884_nl : STD_LOGIC;
  SIGNAL mux_1883_nl : STD_LOGIC;
  SIGNAL mux_1882_nl : STD_LOGIC;
  SIGNAL nor_1022_nl : STD_LOGIC;
  SIGNAL nor_1023_nl : STD_LOGIC;
  SIGNAL mux_1881_nl : STD_LOGIC;
  SIGNAL nor_1024_nl : STD_LOGIC;
  SIGNAL nor_1025_nl : STD_LOGIC;
  SIGNAL mux_1880_nl : STD_LOGIC;
  SIGNAL mux_1879_nl : STD_LOGIC;
  SIGNAL nor_1026_nl : STD_LOGIC;
  SIGNAL nor_1027_nl : STD_LOGIC;
  SIGNAL mux_1878_nl : STD_LOGIC;
  SIGNAL nor_1028_nl : STD_LOGIC;
  SIGNAL nor_1029_nl : STD_LOGIC;
  SIGNAL or_4106_nl : STD_LOGIC;
  SIGNAL mux_1877_nl : STD_LOGIC;
  SIGNAL mux_1876_nl : STD_LOGIC;
  SIGNAL mux_1875_nl : STD_LOGIC;
  SIGNAL or_2198_nl : STD_LOGIC;
  SIGNAL mux_1874_nl : STD_LOGIC;
  SIGNAL or_2195_nl : STD_LOGIC;
  SIGNAL mux_1873_nl : STD_LOGIC;
  SIGNAL mux_1872_nl : STD_LOGIC;
  SIGNAL or_2192_nl : STD_LOGIC;
  SIGNAL mux_1871_nl : STD_LOGIC;
  SIGNAL or_2189_nl : STD_LOGIC;
  SIGNAL mux_1900_nl : STD_LOGIC;
  SIGNAL mux_1899_nl : STD_LOGIC;
  SIGNAL or_2232_nl : STD_LOGIC;
  SIGNAL mux_1898_nl : STD_LOGIC;
  SIGNAL or_2231_nl : STD_LOGIC;
  SIGNAL or_2230_nl : STD_LOGIC;
  SIGNAL mux_1897_nl : STD_LOGIC;
  SIGNAL mux_1896_nl : STD_LOGIC;
  SIGNAL mux_1895_nl : STD_LOGIC;
  SIGNAL or_2228_nl : STD_LOGIC;
  SIGNAL mux_1894_nl : STD_LOGIC;
  SIGNAL or_2226_nl : STD_LOGIC;
  SIGNAL mux_1893_nl : STD_LOGIC;
  SIGNAL mux_1892_nl : STD_LOGIC;
  SIGNAL or_2225_nl : STD_LOGIC;
  SIGNAL mux_1891_nl : STD_LOGIC;
  SIGNAL or_2223_nl : STD_LOGIC;
  SIGNAL or_2222_nl : STD_LOGIC;
  SIGNAL mux_1890_nl : STD_LOGIC;
  SIGNAL mux_1889_nl : STD_LOGIC;
  SIGNAL mux_1888_nl : STD_LOGIC;
  SIGNAL or_2221_nl : STD_LOGIC;
  SIGNAL or_2219_nl : STD_LOGIC;
  SIGNAL mux_1887_nl : STD_LOGIC;
  SIGNAL or_2217_nl : STD_LOGIC;
  SIGNAL or_2216_nl : STD_LOGIC;
  SIGNAL nand_87_nl : STD_LOGIC;
  SIGNAL mux_1886_nl : STD_LOGIC;
  SIGNAL nor_1020_nl : STD_LOGIC;
  SIGNAL nor_1021_nl : STD_LOGIC;
  SIGNAL mux_1915_nl : STD_LOGIC;
  SIGNAL nand_432_nl : STD_LOGIC;
  SIGNAL mux_1914_nl : STD_LOGIC;
  SIGNAL mux_1913_nl : STD_LOGIC;
  SIGNAL mux_1912_nl : STD_LOGIC;
  SIGNAL nor_1011_nl : STD_LOGIC;
  SIGNAL nor_1012_nl : STD_LOGIC;
  SIGNAL mux_1911_nl : STD_LOGIC;
  SIGNAL nor_1013_nl : STD_LOGIC;
  SIGNAL nor_1014_nl : STD_LOGIC;
  SIGNAL mux_1910_nl : STD_LOGIC;
  SIGNAL mux_1909_nl : STD_LOGIC;
  SIGNAL nor_1015_nl : STD_LOGIC;
  SIGNAL nor_1016_nl : STD_LOGIC;
  SIGNAL mux_1908_nl : STD_LOGIC;
  SIGNAL nor_1017_nl : STD_LOGIC;
  SIGNAL nor_1018_nl : STD_LOGIC;
  SIGNAL or_4105_nl : STD_LOGIC;
  SIGNAL mux_1907_nl : STD_LOGIC;
  SIGNAL mux_1906_nl : STD_LOGIC;
  SIGNAL mux_1905_nl : STD_LOGIC;
  SIGNAL or_2242_nl : STD_LOGIC;
  SIGNAL mux_1904_nl : STD_LOGIC;
  SIGNAL or_2239_nl : STD_LOGIC;
  SIGNAL mux_1903_nl : STD_LOGIC;
  SIGNAL mux_1902_nl : STD_LOGIC;
  SIGNAL or_2236_nl : STD_LOGIC;
  SIGNAL mux_1901_nl : STD_LOGIC;
  SIGNAL or_2233_nl : STD_LOGIC;
  SIGNAL mux_1930_nl : STD_LOGIC;
  SIGNAL mux_1929_nl : STD_LOGIC;
  SIGNAL or_2276_nl : STD_LOGIC;
  SIGNAL mux_1928_nl : STD_LOGIC;
  SIGNAL or_2275_nl : STD_LOGIC;
  SIGNAL or_2274_nl : STD_LOGIC;
  SIGNAL mux_1927_nl : STD_LOGIC;
  SIGNAL mux_1926_nl : STD_LOGIC;
  SIGNAL mux_1925_nl : STD_LOGIC;
  SIGNAL or_2272_nl : STD_LOGIC;
  SIGNAL mux_1924_nl : STD_LOGIC;
  SIGNAL or_2270_nl : STD_LOGIC;
  SIGNAL mux_1923_nl : STD_LOGIC;
  SIGNAL mux_1922_nl : STD_LOGIC;
  SIGNAL or_2269_nl : STD_LOGIC;
  SIGNAL mux_1921_nl : STD_LOGIC;
  SIGNAL or_2267_nl : STD_LOGIC;
  SIGNAL or_2266_nl : STD_LOGIC;
  SIGNAL mux_1920_nl : STD_LOGIC;
  SIGNAL mux_1919_nl : STD_LOGIC;
  SIGNAL mux_1918_nl : STD_LOGIC;
  SIGNAL or_2265_nl : STD_LOGIC;
  SIGNAL or_2263_nl : STD_LOGIC;
  SIGNAL mux_1917_nl : STD_LOGIC;
  SIGNAL or_2261_nl : STD_LOGIC;
  SIGNAL or_2260_nl : STD_LOGIC;
  SIGNAL nand_89_nl : STD_LOGIC;
  SIGNAL mux_1916_nl : STD_LOGIC;
  SIGNAL nor_1009_nl : STD_LOGIC;
  SIGNAL nor_1010_nl : STD_LOGIC;
  SIGNAL mux_1945_nl : STD_LOGIC;
  SIGNAL nand_431_nl : STD_LOGIC;
  SIGNAL mux_1944_nl : STD_LOGIC;
  SIGNAL mux_1943_nl : STD_LOGIC;
  SIGNAL mux_1942_nl : STD_LOGIC;
  SIGNAL nor_1000_nl : STD_LOGIC;
  SIGNAL nor_1001_nl : STD_LOGIC;
  SIGNAL mux_1941_nl : STD_LOGIC;
  SIGNAL nor_1002_nl : STD_LOGIC;
  SIGNAL nor_1003_nl : STD_LOGIC;
  SIGNAL mux_1940_nl : STD_LOGIC;
  SIGNAL mux_1939_nl : STD_LOGIC;
  SIGNAL nor_1004_nl : STD_LOGIC;
  SIGNAL nor_1005_nl : STD_LOGIC;
  SIGNAL mux_1938_nl : STD_LOGIC;
  SIGNAL nor_1006_nl : STD_LOGIC;
  SIGNAL nor_1007_nl : STD_LOGIC;
  SIGNAL or_4104_nl : STD_LOGIC;
  SIGNAL mux_1937_nl : STD_LOGIC;
  SIGNAL mux_1936_nl : STD_LOGIC;
  SIGNAL mux_1935_nl : STD_LOGIC;
  SIGNAL or_2286_nl : STD_LOGIC;
  SIGNAL mux_1934_nl : STD_LOGIC;
  SIGNAL or_2283_nl : STD_LOGIC;
  SIGNAL mux_1933_nl : STD_LOGIC;
  SIGNAL mux_1932_nl : STD_LOGIC;
  SIGNAL or_2280_nl : STD_LOGIC;
  SIGNAL mux_1931_nl : STD_LOGIC;
  SIGNAL or_2277_nl : STD_LOGIC;
  SIGNAL mux_1960_nl : STD_LOGIC;
  SIGNAL mux_1959_nl : STD_LOGIC;
  SIGNAL or_2320_nl : STD_LOGIC;
  SIGNAL mux_1958_nl : STD_LOGIC;
  SIGNAL or_2319_nl : STD_LOGIC;
  SIGNAL or_2318_nl : STD_LOGIC;
  SIGNAL mux_1957_nl : STD_LOGIC;
  SIGNAL mux_1956_nl : STD_LOGIC;
  SIGNAL mux_1955_nl : STD_LOGIC;
  SIGNAL or_2316_nl : STD_LOGIC;
  SIGNAL mux_1954_nl : STD_LOGIC;
  SIGNAL or_2314_nl : STD_LOGIC;
  SIGNAL mux_1953_nl : STD_LOGIC;
  SIGNAL mux_1952_nl : STD_LOGIC;
  SIGNAL or_2313_nl : STD_LOGIC;
  SIGNAL mux_1951_nl : STD_LOGIC;
  SIGNAL or_2311_nl : STD_LOGIC;
  SIGNAL or_2310_nl : STD_LOGIC;
  SIGNAL mux_1950_nl : STD_LOGIC;
  SIGNAL mux_1949_nl : STD_LOGIC;
  SIGNAL mux_1948_nl : STD_LOGIC;
  SIGNAL or_2309_nl : STD_LOGIC;
  SIGNAL or_2307_nl : STD_LOGIC;
  SIGNAL mux_1947_nl : STD_LOGIC;
  SIGNAL or_2305_nl : STD_LOGIC;
  SIGNAL or_2304_nl : STD_LOGIC;
  SIGNAL nand_91_nl : STD_LOGIC;
  SIGNAL mux_1946_nl : STD_LOGIC;
  SIGNAL nor_998_nl : STD_LOGIC;
  SIGNAL nor_999_nl : STD_LOGIC;
  SIGNAL mux_1975_nl : STD_LOGIC;
  SIGNAL nand_430_nl : STD_LOGIC;
  SIGNAL mux_1974_nl : STD_LOGIC;
  SIGNAL mux_1973_nl : STD_LOGIC;
  SIGNAL mux_1972_nl : STD_LOGIC;
  SIGNAL and_590_nl : STD_LOGIC;
  SIGNAL nor_990_nl : STD_LOGIC;
  SIGNAL mux_1971_nl : STD_LOGIC;
  SIGNAL nor_991_nl : STD_LOGIC;
  SIGNAL nor_992_nl : STD_LOGIC;
  SIGNAL mux_1970_nl : STD_LOGIC;
  SIGNAL mux_1969_nl : STD_LOGIC;
  SIGNAL nor_993_nl : STD_LOGIC;
  SIGNAL nor_994_nl : STD_LOGIC;
  SIGNAL mux_1968_nl : STD_LOGIC;
  SIGNAL nor_995_nl : STD_LOGIC;
  SIGNAL nor_996_nl : STD_LOGIC;
  SIGNAL or_4103_nl : STD_LOGIC;
  SIGNAL mux_1967_nl : STD_LOGIC;
  SIGNAL mux_1966_nl : STD_LOGIC;
  SIGNAL mux_1965_nl : STD_LOGIC;
  SIGNAL or_2330_nl : STD_LOGIC;
  SIGNAL mux_1964_nl : STD_LOGIC;
  SIGNAL or_2327_nl : STD_LOGIC;
  SIGNAL mux_1963_nl : STD_LOGIC;
  SIGNAL mux_1962_nl : STD_LOGIC;
  SIGNAL or_2324_nl : STD_LOGIC;
  SIGNAL mux_1961_nl : STD_LOGIC;
  SIGNAL or_2321_nl : STD_LOGIC;
  SIGNAL mux_1990_nl : STD_LOGIC;
  SIGNAL mux_1989_nl : STD_LOGIC;
  SIGNAL or_2364_nl : STD_LOGIC;
  SIGNAL mux_1988_nl : STD_LOGIC;
  SIGNAL or_2363_nl : STD_LOGIC;
  SIGNAL or_2362_nl : STD_LOGIC;
  SIGNAL mux_1987_nl : STD_LOGIC;
  SIGNAL mux_1986_nl : STD_LOGIC;
  SIGNAL mux_1985_nl : STD_LOGIC;
  SIGNAL or_2360_nl : STD_LOGIC;
  SIGNAL mux_1984_nl : STD_LOGIC;
  SIGNAL or_2358_nl : STD_LOGIC;
  SIGNAL mux_1983_nl : STD_LOGIC;
  SIGNAL mux_1982_nl : STD_LOGIC;
  SIGNAL or_2357_nl : STD_LOGIC;
  SIGNAL mux_1981_nl : STD_LOGIC;
  SIGNAL or_2355_nl : STD_LOGIC;
  SIGNAL or_2354_nl : STD_LOGIC;
  SIGNAL mux_1980_nl : STD_LOGIC;
  SIGNAL mux_1979_nl : STD_LOGIC;
  SIGNAL mux_1978_nl : STD_LOGIC;
  SIGNAL or_2353_nl : STD_LOGIC;
  SIGNAL nand_296_nl : STD_LOGIC;
  SIGNAL mux_1977_nl : STD_LOGIC;
  SIGNAL or_2349_nl : STD_LOGIC;
  SIGNAL or_2348_nl : STD_LOGIC;
  SIGNAL nand_93_nl : STD_LOGIC;
  SIGNAL mux_1976_nl : STD_LOGIC;
  SIGNAL nor_988_nl : STD_LOGIC;
  SIGNAL nor_989_nl : STD_LOGIC;
  SIGNAL mux_2005_nl : STD_LOGIC;
  SIGNAL nand_429_nl : STD_LOGIC;
  SIGNAL mux_2004_nl : STD_LOGIC;
  SIGNAL mux_2003_nl : STD_LOGIC;
  SIGNAL mux_2002_nl : STD_LOGIC;
  SIGNAL nor_979_nl : STD_LOGIC;
  SIGNAL nor_980_nl : STD_LOGIC;
  SIGNAL mux_2001_nl : STD_LOGIC;
  SIGNAL nor_981_nl : STD_LOGIC;
  SIGNAL nor_982_nl : STD_LOGIC;
  SIGNAL mux_2000_nl : STD_LOGIC;
  SIGNAL mux_1999_nl : STD_LOGIC;
  SIGNAL nor_983_nl : STD_LOGIC;
  SIGNAL nor_984_nl : STD_LOGIC;
  SIGNAL mux_1998_nl : STD_LOGIC;
  SIGNAL nor_985_nl : STD_LOGIC;
  SIGNAL nor_986_nl : STD_LOGIC;
  SIGNAL or_4102_nl : STD_LOGIC;
  SIGNAL mux_1997_nl : STD_LOGIC;
  SIGNAL mux_1996_nl : STD_LOGIC;
  SIGNAL mux_1995_nl : STD_LOGIC;
  SIGNAL or_2374_nl : STD_LOGIC;
  SIGNAL mux_1994_nl : STD_LOGIC;
  SIGNAL or_2371_nl : STD_LOGIC;
  SIGNAL mux_1993_nl : STD_LOGIC;
  SIGNAL mux_1992_nl : STD_LOGIC;
  SIGNAL or_2368_nl : STD_LOGIC;
  SIGNAL mux_1991_nl : STD_LOGIC;
  SIGNAL or_2365_nl : STD_LOGIC;
  SIGNAL mux_2020_nl : STD_LOGIC;
  SIGNAL mux_2019_nl : STD_LOGIC;
  SIGNAL or_2408_nl : STD_LOGIC;
  SIGNAL mux_2018_nl : STD_LOGIC;
  SIGNAL or_2407_nl : STD_LOGIC;
  SIGNAL or_2406_nl : STD_LOGIC;
  SIGNAL mux_2017_nl : STD_LOGIC;
  SIGNAL mux_2016_nl : STD_LOGIC;
  SIGNAL mux_2015_nl : STD_LOGIC;
  SIGNAL or_2404_nl : STD_LOGIC;
  SIGNAL mux_2014_nl : STD_LOGIC;
  SIGNAL or_2402_nl : STD_LOGIC;
  SIGNAL mux_2013_nl : STD_LOGIC;
  SIGNAL mux_2012_nl : STD_LOGIC;
  SIGNAL or_2401_nl : STD_LOGIC;
  SIGNAL mux_2011_nl : STD_LOGIC;
  SIGNAL or_2399_nl : STD_LOGIC;
  SIGNAL or_2398_nl : STD_LOGIC;
  SIGNAL mux_2010_nl : STD_LOGIC;
  SIGNAL mux_2009_nl : STD_LOGIC;
  SIGNAL mux_2008_nl : STD_LOGIC;
  SIGNAL or_2397_nl : STD_LOGIC;
  SIGNAL or_2395_nl : STD_LOGIC;
  SIGNAL mux_2007_nl : STD_LOGIC;
  SIGNAL or_2393_nl : STD_LOGIC;
  SIGNAL or_2392_nl : STD_LOGIC;
  SIGNAL nand_95_nl : STD_LOGIC;
  SIGNAL mux_2006_nl : STD_LOGIC;
  SIGNAL nor_977_nl : STD_LOGIC;
  SIGNAL nor_978_nl : STD_LOGIC;
  SIGNAL mux_2035_nl : STD_LOGIC;
  SIGNAL nand_428_nl : STD_LOGIC;
  SIGNAL mux_2034_nl : STD_LOGIC;
  SIGNAL mux_2033_nl : STD_LOGIC;
  SIGNAL mux_2032_nl : STD_LOGIC;
  SIGNAL nor_968_nl : STD_LOGIC;
  SIGNAL nor_969_nl : STD_LOGIC;
  SIGNAL mux_2031_nl : STD_LOGIC;
  SIGNAL nor_970_nl : STD_LOGIC;
  SIGNAL nor_971_nl : STD_LOGIC;
  SIGNAL mux_2030_nl : STD_LOGIC;
  SIGNAL mux_2029_nl : STD_LOGIC;
  SIGNAL nor_972_nl : STD_LOGIC;
  SIGNAL nor_973_nl : STD_LOGIC;
  SIGNAL mux_2028_nl : STD_LOGIC;
  SIGNAL nor_974_nl : STD_LOGIC;
  SIGNAL nor_975_nl : STD_LOGIC;
  SIGNAL or_4101_nl : STD_LOGIC;
  SIGNAL mux_2027_nl : STD_LOGIC;
  SIGNAL mux_2026_nl : STD_LOGIC;
  SIGNAL mux_2025_nl : STD_LOGIC;
  SIGNAL or_2418_nl : STD_LOGIC;
  SIGNAL mux_2024_nl : STD_LOGIC;
  SIGNAL or_2415_nl : STD_LOGIC;
  SIGNAL mux_2023_nl : STD_LOGIC;
  SIGNAL mux_2022_nl : STD_LOGIC;
  SIGNAL or_2412_nl : STD_LOGIC;
  SIGNAL mux_2021_nl : STD_LOGIC;
  SIGNAL or_2409_nl : STD_LOGIC;
  SIGNAL mux_2050_nl : STD_LOGIC;
  SIGNAL mux_2049_nl : STD_LOGIC;
  SIGNAL or_2452_nl : STD_LOGIC;
  SIGNAL mux_2048_nl : STD_LOGIC;
  SIGNAL or_2451_nl : STD_LOGIC;
  SIGNAL or_2450_nl : STD_LOGIC;
  SIGNAL mux_2047_nl : STD_LOGIC;
  SIGNAL mux_2046_nl : STD_LOGIC;
  SIGNAL mux_2045_nl : STD_LOGIC;
  SIGNAL or_2448_nl : STD_LOGIC;
  SIGNAL mux_2044_nl : STD_LOGIC;
  SIGNAL or_2446_nl : STD_LOGIC;
  SIGNAL mux_2043_nl : STD_LOGIC;
  SIGNAL mux_2042_nl : STD_LOGIC;
  SIGNAL or_2445_nl : STD_LOGIC;
  SIGNAL mux_2041_nl : STD_LOGIC;
  SIGNAL or_2443_nl : STD_LOGIC;
  SIGNAL or_2442_nl : STD_LOGIC;
  SIGNAL mux_2040_nl : STD_LOGIC;
  SIGNAL mux_2039_nl : STD_LOGIC;
  SIGNAL mux_2038_nl : STD_LOGIC;
  SIGNAL or_2441_nl : STD_LOGIC;
  SIGNAL or_2439_nl : STD_LOGIC;
  SIGNAL mux_2037_nl : STD_LOGIC;
  SIGNAL or_2437_nl : STD_LOGIC;
  SIGNAL or_2436_nl : STD_LOGIC;
  SIGNAL nand_97_nl : STD_LOGIC;
  SIGNAL mux_2036_nl : STD_LOGIC;
  SIGNAL nor_966_nl : STD_LOGIC;
  SIGNAL nor_967_nl : STD_LOGIC;
  SIGNAL mux_2065_nl : STD_LOGIC;
  SIGNAL nand_427_nl : STD_LOGIC;
  SIGNAL mux_2064_nl : STD_LOGIC;
  SIGNAL mux_2063_nl : STD_LOGIC;
  SIGNAL mux_2062_nl : STD_LOGIC;
  SIGNAL nor_957_nl : STD_LOGIC;
  SIGNAL nor_958_nl : STD_LOGIC;
  SIGNAL mux_2061_nl : STD_LOGIC;
  SIGNAL nor_959_nl : STD_LOGIC;
  SIGNAL nor_960_nl : STD_LOGIC;
  SIGNAL mux_2060_nl : STD_LOGIC;
  SIGNAL mux_2059_nl : STD_LOGIC;
  SIGNAL nor_961_nl : STD_LOGIC;
  SIGNAL nor_962_nl : STD_LOGIC;
  SIGNAL mux_2058_nl : STD_LOGIC;
  SIGNAL nor_963_nl : STD_LOGIC;
  SIGNAL nor_964_nl : STD_LOGIC;
  SIGNAL or_4100_nl : STD_LOGIC;
  SIGNAL mux_2057_nl : STD_LOGIC;
  SIGNAL mux_2056_nl : STD_LOGIC;
  SIGNAL mux_2055_nl : STD_LOGIC;
  SIGNAL or_2462_nl : STD_LOGIC;
  SIGNAL mux_2054_nl : STD_LOGIC;
  SIGNAL or_2459_nl : STD_LOGIC;
  SIGNAL mux_2053_nl : STD_LOGIC;
  SIGNAL mux_2052_nl : STD_LOGIC;
  SIGNAL or_2456_nl : STD_LOGIC;
  SIGNAL mux_2051_nl : STD_LOGIC;
  SIGNAL or_2453_nl : STD_LOGIC;
  SIGNAL mux_2080_nl : STD_LOGIC;
  SIGNAL mux_2079_nl : STD_LOGIC;
  SIGNAL or_2496_nl : STD_LOGIC;
  SIGNAL mux_2078_nl : STD_LOGIC;
  SIGNAL or_2495_nl : STD_LOGIC;
  SIGNAL or_2494_nl : STD_LOGIC;
  SIGNAL mux_2077_nl : STD_LOGIC;
  SIGNAL mux_2076_nl : STD_LOGIC;
  SIGNAL mux_2075_nl : STD_LOGIC;
  SIGNAL or_2492_nl : STD_LOGIC;
  SIGNAL mux_2074_nl : STD_LOGIC;
  SIGNAL or_2490_nl : STD_LOGIC;
  SIGNAL mux_2073_nl : STD_LOGIC;
  SIGNAL mux_2072_nl : STD_LOGIC;
  SIGNAL or_2489_nl : STD_LOGIC;
  SIGNAL mux_2071_nl : STD_LOGIC;
  SIGNAL or_2487_nl : STD_LOGIC;
  SIGNAL or_2486_nl : STD_LOGIC;
  SIGNAL mux_2070_nl : STD_LOGIC;
  SIGNAL mux_2069_nl : STD_LOGIC;
  SIGNAL mux_2068_nl : STD_LOGIC;
  SIGNAL or_2485_nl : STD_LOGIC;
  SIGNAL or_2483_nl : STD_LOGIC;
  SIGNAL mux_2067_nl : STD_LOGIC;
  SIGNAL or_2481_nl : STD_LOGIC;
  SIGNAL or_2480_nl : STD_LOGIC;
  SIGNAL nand_99_nl : STD_LOGIC;
  SIGNAL mux_2066_nl : STD_LOGIC;
  SIGNAL nor_955_nl : STD_LOGIC;
  SIGNAL nor_956_nl : STD_LOGIC;
  SIGNAL mux_2095_nl : STD_LOGIC;
  SIGNAL nand_426_nl : STD_LOGIC;
  SIGNAL mux_2094_nl : STD_LOGIC;
  SIGNAL mux_2093_nl : STD_LOGIC;
  SIGNAL mux_2092_nl : STD_LOGIC;
  SIGNAL and_585_nl : STD_LOGIC;
  SIGNAL nor_947_nl : STD_LOGIC;
  SIGNAL mux_2091_nl : STD_LOGIC;
  SIGNAL nor_948_nl : STD_LOGIC;
  SIGNAL nor_949_nl : STD_LOGIC;
  SIGNAL mux_2090_nl : STD_LOGIC;
  SIGNAL mux_2089_nl : STD_LOGIC;
  SIGNAL nor_950_nl : STD_LOGIC;
  SIGNAL nor_951_nl : STD_LOGIC;
  SIGNAL mux_2088_nl : STD_LOGIC;
  SIGNAL nor_952_nl : STD_LOGIC;
  SIGNAL nor_953_nl : STD_LOGIC;
  SIGNAL or_4099_nl : STD_LOGIC;
  SIGNAL mux_2087_nl : STD_LOGIC;
  SIGNAL mux_2086_nl : STD_LOGIC;
  SIGNAL mux_2085_nl : STD_LOGIC;
  SIGNAL or_2506_nl : STD_LOGIC;
  SIGNAL mux_2084_nl : STD_LOGIC;
  SIGNAL or_2503_nl : STD_LOGIC;
  SIGNAL mux_2083_nl : STD_LOGIC;
  SIGNAL mux_2082_nl : STD_LOGIC;
  SIGNAL or_2500_nl : STD_LOGIC;
  SIGNAL mux_2081_nl : STD_LOGIC;
  SIGNAL or_2497_nl : STD_LOGIC;
  SIGNAL mux_2110_nl : STD_LOGIC;
  SIGNAL mux_2109_nl : STD_LOGIC;
  SIGNAL or_2540_nl : STD_LOGIC;
  SIGNAL mux_2108_nl : STD_LOGIC;
  SIGNAL or_2539_nl : STD_LOGIC;
  SIGNAL or_2538_nl : STD_LOGIC;
  SIGNAL mux_2107_nl : STD_LOGIC;
  SIGNAL mux_2106_nl : STD_LOGIC;
  SIGNAL mux_2105_nl : STD_LOGIC;
  SIGNAL or_2536_nl : STD_LOGIC;
  SIGNAL mux_2104_nl : STD_LOGIC;
  SIGNAL or_2534_nl : STD_LOGIC;
  SIGNAL mux_2103_nl : STD_LOGIC;
  SIGNAL mux_2102_nl : STD_LOGIC;
  SIGNAL or_2533_nl : STD_LOGIC;
  SIGNAL mux_2101_nl : STD_LOGIC;
  SIGNAL or_2531_nl : STD_LOGIC;
  SIGNAL or_2530_nl : STD_LOGIC;
  SIGNAL mux_2100_nl : STD_LOGIC;
  SIGNAL mux_2099_nl : STD_LOGIC;
  SIGNAL mux_2098_nl : STD_LOGIC;
  SIGNAL or_2529_nl : STD_LOGIC;
  SIGNAL nand_295_nl : STD_LOGIC;
  SIGNAL mux_2097_nl : STD_LOGIC;
  SIGNAL or_2525_nl : STD_LOGIC;
  SIGNAL or_2524_nl : STD_LOGIC;
  SIGNAL nand_101_nl : STD_LOGIC;
  SIGNAL mux_2096_nl : STD_LOGIC;
  SIGNAL nor_945_nl : STD_LOGIC;
  SIGNAL nor_946_nl : STD_LOGIC;
  SIGNAL mux_2125_nl : STD_LOGIC;
  SIGNAL nand_425_nl : STD_LOGIC;
  SIGNAL mux_2124_nl : STD_LOGIC;
  SIGNAL mux_2123_nl : STD_LOGIC;
  SIGNAL mux_2122_nl : STD_LOGIC;
  SIGNAL nor_936_nl : STD_LOGIC;
  SIGNAL nor_937_nl : STD_LOGIC;
  SIGNAL mux_2121_nl : STD_LOGIC;
  SIGNAL nor_938_nl : STD_LOGIC;
  SIGNAL nor_939_nl : STD_LOGIC;
  SIGNAL mux_2120_nl : STD_LOGIC;
  SIGNAL mux_2119_nl : STD_LOGIC;
  SIGNAL nor_940_nl : STD_LOGIC;
  SIGNAL nor_941_nl : STD_LOGIC;
  SIGNAL mux_2118_nl : STD_LOGIC;
  SIGNAL nor_942_nl : STD_LOGIC;
  SIGNAL nor_943_nl : STD_LOGIC;
  SIGNAL or_4098_nl : STD_LOGIC;
  SIGNAL mux_2117_nl : STD_LOGIC;
  SIGNAL mux_2116_nl : STD_LOGIC;
  SIGNAL mux_2115_nl : STD_LOGIC;
  SIGNAL or_2550_nl : STD_LOGIC;
  SIGNAL mux_2114_nl : STD_LOGIC;
  SIGNAL or_2547_nl : STD_LOGIC;
  SIGNAL mux_2113_nl : STD_LOGIC;
  SIGNAL mux_2112_nl : STD_LOGIC;
  SIGNAL or_2544_nl : STD_LOGIC;
  SIGNAL mux_2111_nl : STD_LOGIC;
  SIGNAL or_2541_nl : STD_LOGIC;
  SIGNAL mux_2140_nl : STD_LOGIC;
  SIGNAL mux_2139_nl : STD_LOGIC;
  SIGNAL or_2584_nl : STD_LOGIC;
  SIGNAL mux_2138_nl : STD_LOGIC;
  SIGNAL or_2583_nl : STD_LOGIC;
  SIGNAL or_2582_nl : STD_LOGIC;
  SIGNAL mux_2137_nl : STD_LOGIC;
  SIGNAL mux_2136_nl : STD_LOGIC;
  SIGNAL mux_2135_nl : STD_LOGIC;
  SIGNAL or_2580_nl : STD_LOGIC;
  SIGNAL mux_2134_nl : STD_LOGIC;
  SIGNAL or_2578_nl : STD_LOGIC;
  SIGNAL mux_2133_nl : STD_LOGIC;
  SIGNAL mux_2132_nl : STD_LOGIC;
  SIGNAL or_2577_nl : STD_LOGIC;
  SIGNAL mux_2131_nl : STD_LOGIC;
  SIGNAL or_2575_nl : STD_LOGIC;
  SIGNAL or_2574_nl : STD_LOGIC;
  SIGNAL mux_2130_nl : STD_LOGIC;
  SIGNAL mux_2129_nl : STD_LOGIC;
  SIGNAL mux_2128_nl : STD_LOGIC;
  SIGNAL or_2573_nl : STD_LOGIC;
  SIGNAL or_2571_nl : STD_LOGIC;
  SIGNAL mux_2127_nl : STD_LOGIC;
  SIGNAL or_2569_nl : STD_LOGIC;
  SIGNAL or_2568_nl : STD_LOGIC;
  SIGNAL nand_103_nl : STD_LOGIC;
  SIGNAL mux_2126_nl : STD_LOGIC;
  SIGNAL nor_934_nl : STD_LOGIC;
  SIGNAL nor_935_nl : STD_LOGIC;
  SIGNAL mux_2155_nl : STD_LOGIC;
  SIGNAL nand_424_nl : STD_LOGIC;
  SIGNAL mux_2154_nl : STD_LOGIC;
  SIGNAL mux_2153_nl : STD_LOGIC;
  SIGNAL mux_2152_nl : STD_LOGIC;
  SIGNAL and_582_nl : STD_LOGIC;
  SIGNAL nor_926_nl : STD_LOGIC;
  SIGNAL mux_2151_nl : STD_LOGIC;
  SIGNAL nor_927_nl : STD_LOGIC;
  SIGNAL nor_928_nl : STD_LOGIC;
  SIGNAL mux_2150_nl : STD_LOGIC;
  SIGNAL mux_2149_nl : STD_LOGIC;
  SIGNAL nor_929_nl : STD_LOGIC;
  SIGNAL nor_930_nl : STD_LOGIC;
  SIGNAL mux_2148_nl : STD_LOGIC;
  SIGNAL nor_931_nl : STD_LOGIC;
  SIGNAL nor_932_nl : STD_LOGIC;
  SIGNAL or_4097_nl : STD_LOGIC;
  SIGNAL mux_2147_nl : STD_LOGIC;
  SIGNAL mux_2146_nl : STD_LOGIC;
  SIGNAL mux_2145_nl : STD_LOGIC;
  SIGNAL or_2594_nl : STD_LOGIC;
  SIGNAL mux_2144_nl : STD_LOGIC;
  SIGNAL or_2591_nl : STD_LOGIC;
  SIGNAL mux_2143_nl : STD_LOGIC;
  SIGNAL mux_2142_nl : STD_LOGIC;
  SIGNAL or_2588_nl : STD_LOGIC;
  SIGNAL mux_2141_nl : STD_LOGIC;
  SIGNAL or_2585_nl : STD_LOGIC;
  SIGNAL mux_2170_nl : STD_LOGIC;
  SIGNAL mux_2169_nl : STD_LOGIC;
  SIGNAL or_2628_nl : STD_LOGIC;
  SIGNAL mux_2168_nl : STD_LOGIC;
  SIGNAL or_2627_nl : STD_LOGIC;
  SIGNAL or_2626_nl : STD_LOGIC;
  SIGNAL mux_2167_nl : STD_LOGIC;
  SIGNAL mux_2166_nl : STD_LOGIC;
  SIGNAL mux_2165_nl : STD_LOGIC;
  SIGNAL or_2624_nl : STD_LOGIC;
  SIGNAL mux_2164_nl : STD_LOGIC;
  SIGNAL or_2622_nl : STD_LOGIC;
  SIGNAL mux_2163_nl : STD_LOGIC;
  SIGNAL mux_2162_nl : STD_LOGIC;
  SIGNAL or_2621_nl : STD_LOGIC;
  SIGNAL mux_2161_nl : STD_LOGIC;
  SIGNAL or_2619_nl : STD_LOGIC;
  SIGNAL or_2618_nl : STD_LOGIC;
  SIGNAL mux_2160_nl : STD_LOGIC;
  SIGNAL mux_2159_nl : STD_LOGIC;
  SIGNAL mux_2158_nl : STD_LOGIC;
  SIGNAL or_2617_nl : STD_LOGIC;
  SIGNAL nand_294_nl : STD_LOGIC;
  SIGNAL mux_2157_nl : STD_LOGIC;
  SIGNAL or_2613_nl : STD_LOGIC;
  SIGNAL or_2612_nl : STD_LOGIC;
  SIGNAL nand_105_nl : STD_LOGIC;
  SIGNAL mux_2156_nl : STD_LOGIC;
  SIGNAL nor_924_nl : STD_LOGIC;
  SIGNAL nor_925_nl : STD_LOGIC;
  SIGNAL mux_2185_nl : STD_LOGIC;
  SIGNAL nand_423_nl : STD_LOGIC;
  SIGNAL mux_2184_nl : STD_LOGIC;
  SIGNAL mux_2183_nl : STD_LOGIC;
  SIGNAL mux_2182_nl : STD_LOGIC;
  SIGNAL and_579_nl : STD_LOGIC;
  SIGNAL and_580_nl : STD_LOGIC;
  SIGNAL mux_2181_nl : STD_LOGIC;
  SIGNAL nor_917_nl : STD_LOGIC;
  SIGNAL nor_918_nl : STD_LOGIC;
  SIGNAL mux_2180_nl : STD_LOGIC;
  SIGNAL mux_2179_nl : STD_LOGIC;
  SIGNAL nor_919_nl : STD_LOGIC;
  SIGNAL nor_920_nl : STD_LOGIC;
  SIGNAL mux_2178_nl : STD_LOGIC;
  SIGNAL nor_921_nl : STD_LOGIC;
  SIGNAL nor_922_nl : STD_LOGIC;
  SIGNAL or_4096_nl : STD_LOGIC;
  SIGNAL mux_2177_nl : STD_LOGIC;
  SIGNAL mux_2176_nl : STD_LOGIC;
  SIGNAL mux_2175_nl : STD_LOGIC;
  SIGNAL or_2638_nl : STD_LOGIC;
  SIGNAL mux_2174_nl : STD_LOGIC;
  SIGNAL or_2635_nl : STD_LOGIC;
  SIGNAL mux_2173_nl : STD_LOGIC;
  SIGNAL mux_2172_nl : STD_LOGIC;
  SIGNAL or_2632_nl : STD_LOGIC;
  SIGNAL mux_2171_nl : STD_LOGIC;
  SIGNAL or_2629_nl : STD_LOGIC;
  SIGNAL mux_2200_nl : STD_LOGIC;
  SIGNAL mux_2199_nl : STD_LOGIC;
  SIGNAL or_2672_nl : STD_LOGIC;
  SIGNAL mux_2198_nl : STD_LOGIC;
  SIGNAL or_2671_nl : STD_LOGIC;
  SIGNAL or_2670_nl : STD_LOGIC;
  SIGNAL mux_2197_nl : STD_LOGIC;
  SIGNAL mux_2196_nl : STD_LOGIC;
  SIGNAL mux_2195_nl : STD_LOGIC;
  SIGNAL or_2668_nl : STD_LOGIC;
  SIGNAL mux_2194_nl : STD_LOGIC;
  SIGNAL or_2666_nl : STD_LOGIC;
  SIGNAL mux_2193_nl : STD_LOGIC;
  SIGNAL mux_2192_nl : STD_LOGIC;
  SIGNAL or_2665_nl : STD_LOGIC;
  SIGNAL mux_2191_nl : STD_LOGIC;
  SIGNAL or_2663_nl : STD_LOGIC;
  SIGNAL or_2662_nl : STD_LOGIC;
  SIGNAL mux_2190_nl : STD_LOGIC;
  SIGNAL mux_2189_nl : STD_LOGIC;
  SIGNAL mux_2188_nl : STD_LOGIC;
  SIGNAL nand_292_nl : STD_LOGIC;
  SIGNAL nand_293_nl : STD_LOGIC;
  SIGNAL mux_2187_nl : STD_LOGIC;
  SIGNAL or_2657_nl : STD_LOGIC;
  SIGNAL or_2656_nl : STD_LOGIC;
  SIGNAL nand_107_nl : STD_LOGIC;
  SIGNAL mux_2186_nl : STD_LOGIC;
  SIGNAL nor_915_nl : STD_LOGIC;
  SIGNAL nor_916_nl : STD_LOGIC;
  SIGNAL mux_2215_nl : STD_LOGIC;
  SIGNAL nand_422_nl : STD_LOGIC;
  SIGNAL mux_2214_nl : STD_LOGIC;
  SIGNAL mux_2213_nl : STD_LOGIC;
  SIGNAL mux_2212_nl : STD_LOGIC;
  SIGNAL and_575_nl : STD_LOGIC;
  SIGNAL nor_909_nl : STD_LOGIC;
  SIGNAL mux_2211_nl : STD_LOGIC;
  SIGNAL and_576_nl : STD_LOGIC;
  SIGNAL and_577_nl : STD_LOGIC;
  SIGNAL mux_2210_nl : STD_LOGIC;
  SIGNAL mux_2209_nl : STD_LOGIC;
  SIGNAL and_812_nl : STD_LOGIC;
  SIGNAL and_819_nl : STD_LOGIC;
  SIGNAL mux_2208_nl : STD_LOGIC;
  SIGNAL nor_912_nl : STD_LOGIC;
  SIGNAL nor_913_nl : STD_LOGIC;
  SIGNAL or_4095_nl : STD_LOGIC;
  SIGNAL mux_2207_nl : STD_LOGIC;
  SIGNAL mux_2206_nl : STD_LOGIC;
  SIGNAL mux_2205_nl : STD_LOGIC;
  SIGNAL or_2682_nl : STD_LOGIC;
  SIGNAL mux_2204_nl : STD_LOGIC;
  SIGNAL nand_287_nl : STD_LOGIC;
  SIGNAL mux_2203_nl : STD_LOGIC;
  SIGNAL mux_2202_nl : STD_LOGIC;
  SIGNAL nand_477_nl : STD_LOGIC;
  SIGNAL mux_2201_nl : STD_LOGIC;
  SIGNAL or_2673_nl : STD_LOGIC;
  SIGNAL mux_2230_nl : STD_LOGIC;
  SIGNAL mux_2229_nl : STD_LOGIC;
  SIGNAL or_2715_nl : STD_LOGIC;
  SIGNAL mux_2228_nl : STD_LOGIC;
  SIGNAL or_2714_nl : STD_LOGIC;
  SIGNAL or_2713_nl : STD_LOGIC;
  SIGNAL mux_2227_nl : STD_LOGIC;
  SIGNAL mux_2226_nl : STD_LOGIC;
  SIGNAL mux_2225_nl : STD_LOGIC;
  SIGNAL or_2711_nl : STD_LOGIC;
  SIGNAL mux_2224_nl : STD_LOGIC;
  SIGNAL nand_278_nl : STD_LOGIC;
  SIGNAL mux_2223_nl : STD_LOGIC;
  SIGNAL mux_2222_nl : STD_LOGIC;
  SIGNAL nand_402_nl : STD_LOGIC;
  SIGNAL mux_2221_nl : STD_LOGIC;
  SIGNAL or_2706_nl : STD_LOGIC;
  SIGNAL or_2705_nl : STD_LOGIC;
  SIGNAL mux_2220_nl : STD_LOGIC;
  SIGNAL mux_2219_nl : STD_LOGIC;
  SIGNAL mux_2218_nl : STD_LOGIC;
  SIGNAL or_2704_nl : STD_LOGIC;
  SIGNAL nand_281_nl : STD_LOGIC;
  SIGNAL mux_2217_nl : STD_LOGIC;
  SIGNAL nand_282_nl : STD_LOGIC;
  SIGNAL nand_283_nl : STD_LOGIC;
  SIGNAL nand_109_nl : STD_LOGIC;
  SIGNAL mux_2216_nl : STD_LOGIC;
  SIGNAL nor_907_nl : STD_LOGIC;
  SIGNAL nor_908_nl : STD_LOGIC;
  SIGNAL mux_2245_nl : STD_LOGIC;
  SIGNAL nand_421_nl : STD_LOGIC;
  SIGNAL mux_2244_nl : STD_LOGIC;
  SIGNAL mux_2243_nl : STD_LOGIC;
  SIGNAL mux_2242_nl : STD_LOGIC;
  SIGNAL nor_898_nl : STD_LOGIC;
  SIGNAL nor_899_nl : STD_LOGIC;
  SIGNAL mux_2241_nl : STD_LOGIC;
  SIGNAL nor_900_nl : STD_LOGIC;
  SIGNAL nor_901_nl : STD_LOGIC;
  SIGNAL mux_2240_nl : STD_LOGIC;
  SIGNAL mux_2239_nl : STD_LOGIC;
  SIGNAL nor_902_nl : STD_LOGIC;
  SIGNAL nor_903_nl : STD_LOGIC;
  SIGNAL mux_2238_nl : STD_LOGIC;
  SIGNAL nor_904_nl : STD_LOGIC;
  SIGNAL nor_905_nl : STD_LOGIC;
  SIGNAL or_4094_nl : STD_LOGIC;
  SIGNAL mux_2237_nl : STD_LOGIC;
  SIGNAL mux_2236_nl : STD_LOGIC;
  SIGNAL mux_2235_nl : STD_LOGIC;
  SIGNAL or_2725_nl : STD_LOGIC;
  SIGNAL mux_2234_nl : STD_LOGIC;
  SIGNAL or_2722_nl : STD_LOGIC;
  SIGNAL mux_2233_nl : STD_LOGIC;
  SIGNAL mux_2232_nl : STD_LOGIC;
  SIGNAL or_2719_nl : STD_LOGIC;
  SIGNAL mux_2231_nl : STD_LOGIC;
  SIGNAL or_2716_nl : STD_LOGIC;
  SIGNAL mux_2260_nl : STD_LOGIC;
  SIGNAL mux_2259_nl : STD_LOGIC;
  SIGNAL or_2759_nl : STD_LOGIC;
  SIGNAL mux_2258_nl : STD_LOGIC;
  SIGNAL or_2758_nl : STD_LOGIC;
  SIGNAL or_2757_nl : STD_LOGIC;
  SIGNAL mux_2257_nl : STD_LOGIC;
  SIGNAL mux_2256_nl : STD_LOGIC;
  SIGNAL mux_2255_nl : STD_LOGIC;
  SIGNAL or_2755_nl : STD_LOGIC;
  SIGNAL mux_2254_nl : STD_LOGIC;
  SIGNAL or_2753_nl : STD_LOGIC;
  SIGNAL mux_2253_nl : STD_LOGIC;
  SIGNAL mux_2252_nl : STD_LOGIC;
  SIGNAL or_2752_nl : STD_LOGIC;
  SIGNAL mux_2251_nl : STD_LOGIC;
  SIGNAL or_2750_nl : STD_LOGIC;
  SIGNAL or_2749_nl : STD_LOGIC;
  SIGNAL mux_2250_nl : STD_LOGIC;
  SIGNAL mux_2249_nl : STD_LOGIC;
  SIGNAL mux_2248_nl : STD_LOGIC;
  SIGNAL or_2748_nl : STD_LOGIC;
  SIGNAL or_2746_nl : STD_LOGIC;
  SIGNAL mux_2247_nl : STD_LOGIC;
  SIGNAL or_2744_nl : STD_LOGIC;
  SIGNAL or_2743_nl : STD_LOGIC;
  SIGNAL nand_111_nl : STD_LOGIC;
  SIGNAL mux_2246_nl : STD_LOGIC;
  SIGNAL nor_896_nl : STD_LOGIC;
  SIGNAL nor_897_nl : STD_LOGIC;
  SIGNAL mux_2275_nl : STD_LOGIC;
  SIGNAL nand_420_nl : STD_LOGIC;
  SIGNAL mux_2274_nl : STD_LOGIC;
  SIGNAL mux_2273_nl : STD_LOGIC;
  SIGNAL mux_2272_nl : STD_LOGIC;
  SIGNAL nor_887_nl : STD_LOGIC;
  SIGNAL nor_888_nl : STD_LOGIC;
  SIGNAL mux_2271_nl : STD_LOGIC;
  SIGNAL nor_889_nl : STD_LOGIC;
  SIGNAL nor_890_nl : STD_LOGIC;
  SIGNAL mux_2270_nl : STD_LOGIC;
  SIGNAL mux_2269_nl : STD_LOGIC;
  SIGNAL nor_891_nl : STD_LOGIC;
  SIGNAL nor_892_nl : STD_LOGIC;
  SIGNAL mux_2268_nl : STD_LOGIC;
  SIGNAL nor_893_nl : STD_LOGIC;
  SIGNAL nor_894_nl : STD_LOGIC;
  SIGNAL or_4093_nl : STD_LOGIC;
  SIGNAL mux_2267_nl : STD_LOGIC;
  SIGNAL mux_2266_nl : STD_LOGIC;
  SIGNAL mux_2265_nl : STD_LOGIC;
  SIGNAL or_2769_nl : STD_LOGIC;
  SIGNAL mux_2264_nl : STD_LOGIC;
  SIGNAL or_2766_nl : STD_LOGIC;
  SIGNAL mux_2263_nl : STD_LOGIC;
  SIGNAL mux_2262_nl : STD_LOGIC;
  SIGNAL or_2763_nl : STD_LOGIC;
  SIGNAL mux_2261_nl : STD_LOGIC;
  SIGNAL or_2760_nl : STD_LOGIC;
  SIGNAL mux_2290_nl : STD_LOGIC;
  SIGNAL mux_2289_nl : STD_LOGIC;
  SIGNAL or_2803_nl : STD_LOGIC;
  SIGNAL mux_2288_nl : STD_LOGIC;
  SIGNAL or_2802_nl : STD_LOGIC;
  SIGNAL or_2801_nl : STD_LOGIC;
  SIGNAL mux_2287_nl : STD_LOGIC;
  SIGNAL mux_2286_nl : STD_LOGIC;
  SIGNAL mux_2285_nl : STD_LOGIC;
  SIGNAL or_2799_nl : STD_LOGIC;
  SIGNAL mux_2284_nl : STD_LOGIC;
  SIGNAL or_2797_nl : STD_LOGIC;
  SIGNAL mux_2283_nl : STD_LOGIC;
  SIGNAL mux_2282_nl : STD_LOGIC;
  SIGNAL or_2796_nl : STD_LOGIC;
  SIGNAL mux_2281_nl : STD_LOGIC;
  SIGNAL or_2794_nl : STD_LOGIC;
  SIGNAL or_2793_nl : STD_LOGIC;
  SIGNAL mux_2280_nl : STD_LOGIC;
  SIGNAL mux_2279_nl : STD_LOGIC;
  SIGNAL mux_2278_nl : STD_LOGIC;
  SIGNAL or_2792_nl : STD_LOGIC;
  SIGNAL or_2790_nl : STD_LOGIC;
  SIGNAL mux_2277_nl : STD_LOGIC;
  SIGNAL or_2788_nl : STD_LOGIC;
  SIGNAL or_2787_nl : STD_LOGIC;
  SIGNAL nand_113_nl : STD_LOGIC;
  SIGNAL mux_2276_nl : STD_LOGIC;
  SIGNAL nor_885_nl : STD_LOGIC;
  SIGNAL nor_886_nl : STD_LOGIC;
  SIGNAL mux_2305_nl : STD_LOGIC;
  SIGNAL nand_419_nl : STD_LOGIC;
  SIGNAL mux_2304_nl : STD_LOGIC;
  SIGNAL mux_2303_nl : STD_LOGIC;
  SIGNAL mux_2302_nl : STD_LOGIC;
  SIGNAL nor_876_nl : STD_LOGIC;
  SIGNAL nor_877_nl : STD_LOGIC;
  SIGNAL mux_2301_nl : STD_LOGIC;
  SIGNAL nor_878_nl : STD_LOGIC;
  SIGNAL nor_879_nl : STD_LOGIC;
  SIGNAL mux_2300_nl : STD_LOGIC;
  SIGNAL mux_2299_nl : STD_LOGIC;
  SIGNAL nor_880_nl : STD_LOGIC;
  SIGNAL nor_881_nl : STD_LOGIC;
  SIGNAL mux_2298_nl : STD_LOGIC;
  SIGNAL nor_882_nl : STD_LOGIC;
  SIGNAL nor_883_nl : STD_LOGIC;
  SIGNAL or_4092_nl : STD_LOGIC;
  SIGNAL mux_2297_nl : STD_LOGIC;
  SIGNAL mux_2296_nl : STD_LOGIC;
  SIGNAL mux_2295_nl : STD_LOGIC;
  SIGNAL or_2813_nl : STD_LOGIC;
  SIGNAL mux_2294_nl : STD_LOGIC;
  SIGNAL or_2810_nl : STD_LOGIC;
  SIGNAL mux_2293_nl : STD_LOGIC;
  SIGNAL mux_2292_nl : STD_LOGIC;
  SIGNAL or_2807_nl : STD_LOGIC;
  SIGNAL mux_2291_nl : STD_LOGIC;
  SIGNAL or_2804_nl : STD_LOGIC;
  SIGNAL mux_2320_nl : STD_LOGIC;
  SIGNAL mux_2319_nl : STD_LOGIC;
  SIGNAL or_2847_nl : STD_LOGIC;
  SIGNAL mux_2318_nl : STD_LOGIC;
  SIGNAL or_2846_nl : STD_LOGIC;
  SIGNAL or_2845_nl : STD_LOGIC;
  SIGNAL mux_2317_nl : STD_LOGIC;
  SIGNAL mux_2316_nl : STD_LOGIC;
  SIGNAL mux_2315_nl : STD_LOGIC;
  SIGNAL or_2843_nl : STD_LOGIC;
  SIGNAL mux_2314_nl : STD_LOGIC;
  SIGNAL or_2841_nl : STD_LOGIC;
  SIGNAL mux_2313_nl : STD_LOGIC;
  SIGNAL mux_2312_nl : STD_LOGIC;
  SIGNAL or_2840_nl : STD_LOGIC;
  SIGNAL mux_2311_nl : STD_LOGIC;
  SIGNAL or_2838_nl : STD_LOGIC;
  SIGNAL or_2837_nl : STD_LOGIC;
  SIGNAL mux_2310_nl : STD_LOGIC;
  SIGNAL mux_2309_nl : STD_LOGIC;
  SIGNAL mux_2308_nl : STD_LOGIC;
  SIGNAL or_2836_nl : STD_LOGIC;
  SIGNAL or_2834_nl : STD_LOGIC;
  SIGNAL mux_2307_nl : STD_LOGIC;
  SIGNAL or_2832_nl : STD_LOGIC;
  SIGNAL or_2831_nl : STD_LOGIC;
  SIGNAL nand_115_nl : STD_LOGIC;
  SIGNAL mux_2306_nl : STD_LOGIC;
  SIGNAL nor_874_nl : STD_LOGIC;
  SIGNAL nor_875_nl : STD_LOGIC;
  SIGNAL mux_2335_nl : STD_LOGIC;
  SIGNAL nand_418_nl : STD_LOGIC;
  SIGNAL mux_2334_nl : STD_LOGIC;
  SIGNAL mux_2333_nl : STD_LOGIC;
  SIGNAL mux_2332_nl : STD_LOGIC;
  SIGNAL nor_865_nl : STD_LOGIC;
  SIGNAL nor_866_nl : STD_LOGIC;
  SIGNAL mux_2331_nl : STD_LOGIC;
  SIGNAL nor_867_nl : STD_LOGIC;
  SIGNAL nor_868_nl : STD_LOGIC;
  SIGNAL mux_2330_nl : STD_LOGIC;
  SIGNAL mux_2329_nl : STD_LOGIC;
  SIGNAL nor_869_nl : STD_LOGIC;
  SIGNAL nor_870_nl : STD_LOGIC;
  SIGNAL mux_2328_nl : STD_LOGIC;
  SIGNAL nor_871_nl : STD_LOGIC;
  SIGNAL nor_872_nl : STD_LOGIC;
  SIGNAL or_4091_nl : STD_LOGIC;
  SIGNAL mux_2327_nl : STD_LOGIC;
  SIGNAL mux_2326_nl : STD_LOGIC;
  SIGNAL mux_2325_nl : STD_LOGIC;
  SIGNAL or_2857_nl : STD_LOGIC;
  SIGNAL mux_2324_nl : STD_LOGIC;
  SIGNAL or_2854_nl : STD_LOGIC;
  SIGNAL mux_2323_nl : STD_LOGIC;
  SIGNAL mux_2322_nl : STD_LOGIC;
  SIGNAL or_2851_nl : STD_LOGIC;
  SIGNAL mux_2321_nl : STD_LOGIC;
  SIGNAL or_2848_nl : STD_LOGIC;
  SIGNAL mux_2350_nl : STD_LOGIC;
  SIGNAL mux_2349_nl : STD_LOGIC;
  SIGNAL or_2891_nl : STD_LOGIC;
  SIGNAL mux_2348_nl : STD_LOGIC;
  SIGNAL or_2890_nl : STD_LOGIC;
  SIGNAL or_2889_nl : STD_LOGIC;
  SIGNAL mux_2347_nl : STD_LOGIC;
  SIGNAL mux_2346_nl : STD_LOGIC;
  SIGNAL mux_2345_nl : STD_LOGIC;
  SIGNAL or_2887_nl : STD_LOGIC;
  SIGNAL mux_2344_nl : STD_LOGIC;
  SIGNAL or_2885_nl : STD_LOGIC;
  SIGNAL mux_2343_nl : STD_LOGIC;
  SIGNAL mux_2342_nl : STD_LOGIC;
  SIGNAL or_2884_nl : STD_LOGIC;
  SIGNAL mux_2341_nl : STD_LOGIC;
  SIGNAL or_2882_nl : STD_LOGIC;
  SIGNAL or_2881_nl : STD_LOGIC;
  SIGNAL mux_2340_nl : STD_LOGIC;
  SIGNAL mux_2339_nl : STD_LOGIC;
  SIGNAL mux_2338_nl : STD_LOGIC;
  SIGNAL or_2880_nl : STD_LOGIC;
  SIGNAL or_2878_nl : STD_LOGIC;
  SIGNAL mux_2337_nl : STD_LOGIC;
  SIGNAL or_2876_nl : STD_LOGIC;
  SIGNAL or_2875_nl : STD_LOGIC;
  SIGNAL nand_117_nl : STD_LOGIC;
  SIGNAL mux_2336_nl : STD_LOGIC;
  SIGNAL nor_863_nl : STD_LOGIC;
  SIGNAL nor_864_nl : STD_LOGIC;
  SIGNAL mux_2365_nl : STD_LOGIC;
  SIGNAL nand_417_nl : STD_LOGIC;
  SIGNAL mux_2364_nl : STD_LOGIC;
  SIGNAL mux_2363_nl : STD_LOGIC;
  SIGNAL mux_2362_nl : STD_LOGIC;
  SIGNAL nor_854_nl : STD_LOGIC;
  SIGNAL nor_855_nl : STD_LOGIC;
  SIGNAL mux_2361_nl : STD_LOGIC;
  SIGNAL nor_856_nl : STD_LOGIC;
  SIGNAL nor_857_nl : STD_LOGIC;
  SIGNAL mux_2360_nl : STD_LOGIC;
  SIGNAL mux_2359_nl : STD_LOGIC;
  SIGNAL nor_858_nl : STD_LOGIC;
  SIGNAL nor_859_nl : STD_LOGIC;
  SIGNAL mux_2358_nl : STD_LOGIC;
  SIGNAL nor_860_nl : STD_LOGIC;
  SIGNAL nor_861_nl : STD_LOGIC;
  SIGNAL or_4090_nl : STD_LOGIC;
  SIGNAL mux_2357_nl : STD_LOGIC;
  SIGNAL mux_2356_nl : STD_LOGIC;
  SIGNAL mux_2355_nl : STD_LOGIC;
  SIGNAL or_2901_nl : STD_LOGIC;
  SIGNAL mux_2354_nl : STD_LOGIC;
  SIGNAL or_2898_nl : STD_LOGIC;
  SIGNAL mux_2353_nl : STD_LOGIC;
  SIGNAL mux_2352_nl : STD_LOGIC;
  SIGNAL or_2895_nl : STD_LOGIC;
  SIGNAL mux_2351_nl : STD_LOGIC;
  SIGNAL or_2892_nl : STD_LOGIC;
  SIGNAL mux_2380_nl : STD_LOGIC;
  SIGNAL mux_2379_nl : STD_LOGIC;
  SIGNAL or_2935_nl : STD_LOGIC;
  SIGNAL mux_2378_nl : STD_LOGIC;
  SIGNAL or_2934_nl : STD_LOGIC;
  SIGNAL or_2933_nl : STD_LOGIC;
  SIGNAL mux_2377_nl : STD_LOGIC;
  SIGNAL mux_2376_nl : STD_LOGIC;
  SIGNAL mux_2375_nl : STD_LOGIC;
  SIGNAL or_2931_nl : STD_LOGIC;
  SIGNAL mux_2374_nl : STD_LOGIC;
  SIGNAL or_2929_nl : STD_LOGIC;
  SIGNAL mux_2373_nl : STD_LOGIC;
  SIGNAL mux_2372_nl : STD_LOGIC;
  SIGNAL or_2928_nl : STD_LOGIC;
  SIGNAL mux_2371_nl : STD_LOGIC;
  SIGNAL or_2926_nl : STD_LOGIC;
  SIGNAL or_2925_nl : STD_LOGIC;
  SIGNAL mux_2370_nl : STD_LOGIC;
  SIGNAL mux_2369_nl : STD_LOGIC;
  SIGNAL mux_2368_nl : STD_LOGIC;
  SIGNAL or_2924_nl : STD_LOGIC;
  SIGNAL or_2922_nl : STD_LOGIC;
  SIGNAL mux_2367_nl : STD_LOGIC;
  SIGNAL or_2920_nl : STD_LOGIC;
  SIGNAL or_2919_nl : STD_LOGIC;
  SIGNAL nand_119_nl : STD_LOGIC;
  SIGNAL mux_2366_nl : STD_LOGIC;
  SIGNAL nor_852_nl : STD_LOGIC;
  SIGNAL nor_853_nl : STD_LOGIC;
  SIGNAL mux_2395_nl : STD_LOGIC;
  SIGNAL nand_416_nl : STD_LOGIC;
  SIGNAL mux_2394_nl : STD_LOGIC;
  SIGNAL mux_2393_nl : STD_LOGIC;
  SIGNAL mux_2392_nl : STD_LOGIC;
  SIGNAL nor_843_nl : STD_LOGIC;
  SIGNAL nor_844_nl : STD_LOGIC;
  SIGNAL mux_2391_nl : STD_LOGIC;
  SIGNAL nor_845_nl : STD_LOGIC;
  SIGNAL nor_846_nl : STD_LOGIC;
  SIGNAL mux_2390_nl : STD_LOGIC;
  SIGNAL mux_2389_nl : STD_LOGIC;
  SIGNAL nor_847_nl : STD_LOGIC;
  SIGNAL nor_848_nl : STD_LOGIC;
  SIGNAL mux_2388_nl : STD_LOGIC;
  SIGNAL nor_849_nl : STD_LOGIC;
  SIGNAL nor_850_nl : STD_LOGIC;
  SIGNAL or_4089_nl : STD_LOGIC;
  SIGNAL mux_2387_nl : STD_LOGIC;
  SIGNAL mux_2386_nl : STD_LOGIC;
  SIGNAL mux_2385_nl : STD_LOGIC;
  SIGNAL or_2945_nl : STD_LOGIC;
  SIGNAL mux_2384_nl : STD_LOGIC;
  SIGNAL or_2942_nl : STD_LOGIC;
  SIGNAL mux_2383_nl : STD_LOGIC;
  SIGNAL mux_2382_nl : STD_LOGIC;
  SIGNAL or_2939_nl : STD_LOGIC;
  SIGNAL mux_2381_nl : STD_LOGIC;
  SIGNAL or_2936_nl : STD_LOGIC;
  SIGNAL mux_2410_nl : STD_LOGIC;
  SIGNAL mux_2409_nl : STD_LOGIC;
  SIGNAL or_2979_nl : STD_LOGIC;
  SIGNAL mux_2408_nl : STD_LOGIC;
  SIGNAL or_2978_nl : STD_LOGIC;
  SIGNAL or_2977_nl : STD_LOGIC;
  SIGNAL mux_2407_nl : STD_LOGIC;
  SIGNAL mux_2406_nl : STD_LOGIC;
  SIGNAL mux_2405_nl : STD_LOGIC;
  SIGNAL or_2975_nl : STD_LOGIC;
  SIGNAL mux_2404_nl : STD_LOGIC;
  SIGNAL or_2973_nl : STD_LOGIC;
  SIGNAL mux_2403_nl : STD_LOGIC;
  SIGNAL mux_2402_nl : STD_LOGIC;
  SIGNAL or_2972_nl : STD_LOGIC;
  SIGNAL mux_2401_nl : STD_LOGIC;
  SIGNAL or_2970_nl : STD_LOGIC;
  SIGNAL or_2969_nl : STD_LOGIC;
  SIGNAL mux_2400_nl : STD_LOGIC;
  SIGNAL mux_2399_nl : STD_LOGIC;
  SIGNAL mux_2398_nl : STD_LOGIC;
  SIGNAL or_2968_nl : STD_LOGIC;
  SIGNAL or_2966_nl : STD_LOGIC;
  SIGNAL mux_2397_nl : STD_LOGIC;
  SIGNAL or_2964_nl : STD_LOGIC;
  SIGNAL or_2963_nl : STD_LOGIC;
  SIGNAL nand_121_nl : STD_LOGIC;
  SIGNAL mux_2396_nl : STD_LOGIC;
  SIGNAL nor_841_nl : STD_LOGIC;
  SIGNAL nor_842_nl : STD_LOGIC;
  SIGNAL mux_2425_nl : STD_LOGIC;
  SIGNAL nand_415_nl : STD_LOGIC;
  SIGNAL mux_2424_nl : STD_LOGIC;
  SIGNAL mux_2423_nl : STD_LOGIC;
  SIGNAL mux_2422_nl : STD_LOGIC;
  SIGNAL nor_833_nl : STD_LOGIC;
  SIGNAL and_567_nl : STD_LOGIC;
  SIGNAL mux_2421_nl : STD_LOGIC;
  SIGNAL nor_834_nl : STD_LOGIC;
  SIGNAL nor_835_nl : STD_LOGIC;
  SIGNAL mux_2420_nl : STD_LOGIC;
  SIGNAL mux_2419_nl : STD_LOGIC;
  SIGNAL nor_836_nl : STD_LOGIC;
  SIGNAL nor_837_nl : STD_LOGIC;
  SIGNAL mux_2418_nl : STD_LOGIC;
  SIGNAL nor_838_nl : STD_LOGIC;
  SIGNAL nor_839_nl : STD_LOGIC;
  SIGNAL or_4088_nl : STD_LOGIC;
  SIGNAL mux_2417_nl : STD_LOGIC;
  SIGNAL mux_2416_nl : STD_LOGIC;
  SIGNAL mux_2415_nl : STD_LOGIC;
  SIGNAL or_2989_nl : STD_LOGIC;
  SIGNAL mux_2414_nl : STD_LOGIC;
  SIGNAL or_2986_nl : STD_LOGIC;
  SIGNAL mux_2413_nl : STD_LOGIC;
  SIGNAL mux_2412_nl : STD_LOGIC;
  SIGNAL or_2983_nl : STD_LOGIC;
  SIGNAL mux_2411_nl : STD_LOGIC;
  SIGNAL or_2980_nl : STD_LOGIC;
  SIGNAL mux_2440_nl : STD_LOGIC;
  SIGNAL mux_2439_nl : STD_LOGIC;
  SIGNAL or_3023_nl : STD_LOGIC;
  SIGNAL mux_2438_nl : STD_LOGIC;
  SIGNAL or_3022_nl : STD_LOGIC;
  SIGNAL or_3021_nl : STD_LOGIC;
  SIGNAL mux_2437_nl : STD_LOGIC;
  SIGNAL mux_2436_nl : STD_LOGIC;
  SIGNAL mux_2435_nl : STD_LOGIC;
  SIGNAL or_3019_nl : STD_LOGIC;
  SIGNAL mux_2434_nl : STD_LOGIC;
  SIGNAL or_3017_nl : STD_LOGIC;
  SIGNAL mux_2433_nl : STD_LOGIC;
  SIGNAL mux_2432_nl : STD_LOGIC;
  SIGNAL or_3016_nl : STD_LOGIC;
  SIGNAL mux_2431_nl : STD_LOGIC;
  SIGNAL or_3014_nl : STD_LOGIC;
  SIGNAL or_3013_nl : STD_LOGIC;
  SIGNAL mux_2430_nl : STD_LOGIC;
  SIGNAL mux_2429_nl : STD_LOGIC;
  SIGNAL mux_2428_nl : STD_LOGIC;
  SIGNAL nand_271_nl : STD_LOGIC;
  SIGNAL or_3010_nl : STD_LOGIC;
  SIGNAL mux_2427_nl : STD_LOGIC;
  SIGNAL or_3008_nl : STD_LOGIC;
  SIGNAL or_3007_nl : STD_LOGIC;
  SIGNAL nand_123_nl : STD_LOGIC;
  SIGNAL mux_2426_nl : STD_LOGIC;
  SIGNAL nor_831_nl : STD_LOGIC;
  SIGNAL nor_832_nl : STD_LOGIC;
  SIGNAL mux_2455_nl : STD_LOGIC;
  SIGNAL nand_414_nl : STD_LOGIC;
  SIGNAL mux_2454_nl : STD_LOGIC;
  SIGNAL mux_2453_nl : STD_LOGIC;
  SIGNAL mux_2452_nl : STD_LOGIC;
  SIGNAL nor_824_nl : STD_LOGIC;
  SIGNAL nor_825_nl : STD_LOGIC;
  SIGNAL mux_2451_nl : STD_LOGIC;
  SIGNAL and_564_nl : STD_LOGIC;
  SIGNAL and_565_nl : STD_LOGIC;
  SIGNAL mux_2450_nl : STD_LOGIC;
  SIGNAL mux_2449_nl : STD_LOGIC;
  SIGNAL and_813_nl : STD_LOGIC;
  SIGNAL and_820_nl : STD_LOGIC;
  SIGNAL mux_2448_nl : STD_LOGIC;
  SIGNAL nor_828_nl : STD_LOGIC;
  SIGNAL nor_829_nl : STD_LOGIC;
  SIGNAL or_4087_nl : STD_LOGIC;
  SIGNAL mux_2447_nl : STD_LOGIC;
  SIGNAL mux_2446_nl : STD_LOGIC;
  SIGNAL mux_2445_nl : STD_LOGIC;
  SIGNAL or_3033_nl : STD_LOGIC;
  SIGNAL mux_2444_nl : STD_LOGIC;
  SIGNAL nand_267_nl : STD_LOGIC;
  SIGNAL mux_2443_nl : STD_LOGIC;
  SIGNAL mux_2442_nl : STD_LOGIC;
  SIGNAL nand_476_nl : STD_LOGIC;
  SIGNAL mux_2441_nl : STD_LOGIC;
  SIGNAL or_3024_nl : STD_LOGIC;
  SIGNAL mux_2470_nl : STD_LOGIC;
  SIGNAL mux_2469_nl : STD_LOGIC;
  SIGNAL or_3067_nl : STD_LOGIC;
  SIGNAL mux_2468_nl : STD_LOGIC;
  SIGNAL or_3066_nl : STD_LOGIC;
  SIGNAL or_3065_nl : STD_LOGIC;
  SIGNAL mux_2467_nl : STD_LOGIC;
  SIGNAL mux_2466_nl : STD_LOGIC;
  SIGNAL mux_2465_nl : STD_LOGIC;
  SIGNAL or_3063_nl : STD_LOGIC;
  SIGNAL mux_2464_nl : STD_LOGIC;
  SIGNAL nand_258_nl : STD_LOGIC;
  SIGNAL mux_2463_nl : STD_LOGIC;
  SIGNAL mux_2462_nl : STD_LOGIC;
  SIGNAL nand_400_nl : STD_LOGIC;
  SIGNAL mux_2461_nl : STD_LOGIC;
  SIGNAL or_3058_nl : STD_LOGIC;
  SIGNAL or_3057_nl : STD_LOGIC;
  SIGNAL mux_2460_nl : STD_LOGIC;
  SIGNAL mux_2459_nl : STD_LOGIC;
  SIGNAL mux_2458_nl : STD_LOGIC;
  SIGNAL or_3056_nl : STD_LOGIC;
  SIGNAL or_3054_nl : STD_LOGIC;
  SIGNAL mux_2457_nl : STD_LOGIC;
  SIGNAL nand_261_nl : STD_LOGIC;
  SIGNAL nand_262_nl : STD_LOGIC;
  SIGNAL nand_125_nl : STD_LOGIC;
  SIGNAL mux_2456_nl : STD_LOGIC;
  SIGNAL nor_822_nl : STD_LOGIC;
  SIGNAL nor_823_nl : STD_LOGIC;
  SIGNAL mux_2485_nl : STD_LOGIC;
  SIGNAL nand_413_nl : STD_LOGIC;
  SIGNAL mux_2484_nl : STD_LOGIC;
  SIGNAL mux_2483_nl : STD_LOGIC;
  SIGNAL mux_2482_nl : STD_LOGIC;
  SIGNAL nor_813_nl : STD_LOGIC;
  SIGNAL nor_814_nl : STD_LOGIC;
  SIGNAL mux_2481_nl : STD_LOGIC;
  SIGNAL nor_815_nl : STD_LOGIC;
  SIGNAL nor_816_nl : STD_LOGIC;
  SIGNAL mux_2480_nl : STD_LOGIC;
  SIGNAL mux_2479_nl : STD_LOGIC;
  SIGNAL nor_817_nl : STD_LOGIC;
  SIGNAL nor_818_nl : STD_LOGIC;
  SIGNAL mux_2478_nl : STD_LOGIC;
  SIGNAL nor_819_nl : STD_LOGIC;
  SIGNAL nor_820_nl : STD_LOGIC;
  SIGNAL or_4086_nl : STD_LOGIC;
  SIGNAL mux_2477_nl : STD_LOGIC;
  SIGNAL mux_2476_nl : STD_LOGIC;
  SIGNAL mux_2475_nl : STD_LOGIC;
  SIGNAL or_3077_nl : STD_LOGIC;
  SIGNAL mux_2474_nl : STD_LOGIC;
  SIGNAL or_3074_nl : STD_LOGIC;
  SIGNAL mux_2473_nl : STD_LOGIC;
  SIGNAL mux_2472_nl : STD_LOGIC;
  SIGNAL or_3071_nl : STD_LOGIC;
  SIGNAL mux_2471_nl : STD_LOGIC;
  SIGNAL or_3068_nl : STD_LOGIC;
  SIGNAL mux_2500_nl : STD_LOGIC;
  SIGNAL mux_2499_nl : STD_LOGIC;
  SIGNAL or_3111_nl : STD_LOGIC;
  SIGNAL mux_2498_nl : STD_LOGIC;
  SIGNAL or_3110_nl : STD_LOGIC;
  SIGNAL or_3109_nl : STD_LOGIC;
  SIGNAL mux_2497_nl : STD_LOGIC;
  SIGNAL mux_2496_nl : STD_LOGIC;
  SIGNAL mux_2495_nl : STD_LOGIC;
  SIGNAL or_3107_nl : STD_LOGIC;
  SIGNAL mux_2494_nl : STD_LOGIC;
  SIGNAL or_3105_nl : STD_LOGIC;
  SIGNAL mux_2493_nl : STD_LOGIC;
  SIGNAL mux_2492_nl : STD_LOGIC;
  SIGNAL or_3104_nl : STD_LOGIC;
  SIGNAL mux_2491_nl : STD_LOGIC;
  SIGNAL or_3102_nl : STD_LOGIC;
  SIGNAL or_3101_nl : STD_LOGIC;
  SIGNAL mux_2490_nl : STD_LOGIC;
  SIGNAL mux_2489_nl : STD_LOGIC;
  SIGNAL mux_2488_nl : STD_LOGIC;
  SIGNAL or_3100_nl : STD_LOGIC;
  SIGNAL or_3098_nl : STD_LOGIC;
  SIGNAL mux_2487_nl : STD_LOGIC;
  SIGNAL or_3096_nl : STD_LOGIC;
  SIGNAL or_3095_nl : STD_LOGIC;
  SIGNAL nand_127_nl : STD_LOGIC;
  SIGNAL mux_2486_nl : STD_LOGIC;
  SIGNAL nor_811_nl : STD_LOGIC;
  SIGNAL nor_812_nl : STD_LOGIC;
  SIGNAL mux_2515_nl : STD_LOGIC;
  SIGNAL nand_412_nl : STD_LOGIC;
  SIGNAL mux_2514_nl : STD_LOGIC;
  SIGNAL mux_2513_nl : STD_LOGIC;
  SIGNAL mux_2512_nl : STD_LOGIC;
  SIGNAL nor_802_nl : STD_LOGIC;
  SIGNAL nor_803_nl : STD_LOGIC;
  SIGNAL mux_2511_nl : STD_LOGIC;
  SIGNAL nor_804_nl : STD_LOGIC;
  SIGNAL nor_805_nl : STD_LOGIC;
  SIGNAL mux_2510_nl : STD_LOGIC;
  SIGNAL mux_2509_nl : STD_LOGIC;
  SIGNAL nor_806_nl : STD_LOGIC;
  SIGNAL nor_807_nl : STD_LOGIC;
  SIGNAL mux_2508_nl : STD_LOGIC;
  SIGNAL nor_808_nl : STD_LOGIC;
  SIGNAL nor_809_nl : STD_LOGIC;
  SIGNAL or_4085_nl : STD_LOGIC;
  SIGNAL mux_2507_nl : STD_LOGIC;
  SIGNAL mux_2506_nl : STD_LOGIC;
  SIGNAL mux_2505_nl : STD_LOGIC;
  SIGNAL or_3121_nl : STD_LOGIC;
  SIGNAL mux_2504_nl : STD_LOGIC;
  SIGNAL or_3118_nl : STD_LOGIC;
  SIGNAL mux_2503_nl : STD_LOGIC;
  SIGNAL mux_2502_nl : STD_LOGIC;
  SIGNAL or_3115_nl : STD_LOGIC;
  SIGNAL mux_2501_nl : STD_LOGIC;
  SIGNAL or_3112_nl : STD_LOGIC;
  SIGNAL mux_2530_nl : STD_LOGIC;
  SIGNAL mux_2529_nl : STD_LOGIC;
  SIGNAL or_3155_nl : STD_LOGIC;
  SIGNAL mux_2528_nl : STD_LOGIC;
  SIGNAL or_3154_nl : STD_LOGIC;
  SIGNAL or_3153_nl : STD_LOGIC;
  SIGNAL mux_2527_nl : STD_LOGIC;
  SIGNAL mux_2526_nl : STD_LOGIC;
  SIGNAL mux_2525_nl : STD_LOGIC;
  SIGNAL or_3151_nl : STD_LOGIC;
  SIGNAL mux_2524_nl : STD_LOGIC;
  SIGNAL or_3149_nl : STD_LOGIC;
  SIGNAL mux_2523_nl : STD_LOGIC;
  SIGNAL mux_2522_nl : STD_LOGIC;
  SIGNAL or_3148_nl : STD_LOGIC;
  SIGNAL mux_2521_nl : STD_LOGIC;
  SIGNAL or_3146_nl : STD_LOGIC;
  SIGNAL or_3145_nl : STD_LOGIC;
  SIGNAL mux_2520_nl : STD_LOGIC;
  SIGNAL mux_2519_nl : STD_LOGIC;
  SIGNAL mux_2518_nl : STD_LOGIC;
  SIGNAL or_3144_nl : STD_LOGIC;
  SIGNAL or_3142_nl : STD_LOGIC;
  SIGNAL mux_2517_nl : STD_LOGIC;
  SIGNAL or_3140_nl : STD_LOGIC;
  SIGNAL or_3139_nl : STD_LOGIC;
  SIGNAL nand_129_nl : STD_LOGIC;
  SIGNAL mux_2516_nl : STD_LOGIC;
  SIGNAL nor_800_nl : STD_LOGIC;
  SIGNAL nor_801_nl : STD_LOGIC;
  SIGNAL mux_2545_nl : STD_LOGIC;
  SIGNAL nand_411_nl : STD_LOGIC;
  SIGNAL mux_2544_nl : STD_LOGIC;
  SIGNAL mux_2543_nl : STD_LOGIC;
  SIGNAL mux_2542_nl : STD_LOGIC;
  SIGNAL nor_792_nl : STD_LOGIC;
  SIGNAL and_560_nl : STD_LOGIC;
  SIGNAL mux_2541_nl : STD_LOGIC;
  SIGNAL nor_793_nl : STD_LOGIC;
  SIGNAL nor_794_nl : STD_LOGIC;
  SIGNAL mux_2540_nl : STD_LOGIC;
  SIGNAL mux_2539_nl : STD_LOGIC;
  SIGNAL nor_795_nl : STD_LOGIC;
  SIGNAL nor_796_nl : STD_LOGIC;
  SIGNAL mux_2538_nl : STD_LOGIC;
  SIGNAL nor_797_nl : STD_LOGIC;
  SIGNAL nor_798_nl : STD_LOGIC;
  SIGNAL or_4084_nl : STD_LOGIC;
  SIGNAL mux_2537_nl : STD_LOGIC;
  SIGNAL mux_2536_nl : STD_LOGIC;
  SIGNAL mux_2535_nl : STD_LOGIC;
  SIGNAL or_3165_nl : STD_LOGIC;
  SIGNAL mux_2534_nl : STD_LOGIC;
  SIGNAL or_3162_nl : STD_LOGIC;
  SIGNAL mux_2533_nl : STD_LOGIC;
  SIGNAL mux_2532_nl : STD_LOGIC;
  SIGNAL or_3159_nl : STD_LOGIC;
  SIGNAL mux_2531_nl : STD_LOGIC;
  SIGNAL or_3156_nl : STD_LOGIC;
  SIGNAL mux_2560_nl : STD_LOGIC;
  SIGNAL mux_2559_nl : STD_LOGIC;
  SIGNAL or_3199_nl : STD_LOGIC;
  SIGNAL mux_2558_nl : STD_LOGIC;
  SIGNAL or_3198_nl : STD_LOGIC;
  SIGNAL or_3197_nl : STD_LOGIC;
  SIGNAL mux_2557_nl : STD_LOGIC;
  SIGNAL mux_2556_nl : STD_LOGIC;
  SIGNAL mux_2555_nl : STD_LOGIC;
  SIGNAL or_3195_nl : STD_LOGIC;
  SIGNAL mux_2554_nl : STD_LOGIC;
  SIGNAL or_3193_nl : STD_LOGIC;
  SIGNAL mux_2553_nl : STD_LOGIC;
  SIGNAL mux_2552_nl : STD_LOGIC;
  SIGNAL or_3192_nl : STD_LOGIC;
  SIGNAL mux_2551_nl : STD_LOGIC;
  SIGNAL or_3190_nl : STD_LOGIC;
  SIGNAL or_3189_nl : STD_LOGIC;
  SIGNAL mux_2550_nl : STD_LOGIC;
  SIGNAL mux_2549_nl : STD_LOGIC;
  SIGNAL mux_2548_nl : STD_LOGIC;
  SIGNAL nand_252_nl : STD_LOGIC;
  SIGNAL or_3186_nl : STD_LOGIC;
  SIGNAL mux_2547_nl : STD_LOGIC;
  SIGNAL or_3184_nl : STD_LOGIC;
  SIGNAL or_3183_nl : STD_LOGIC;
  SIGNAL nand_131_nl : STD_LOGIC;
  SIGNAL mux_2546_nl : STD_LOGIC;
  SIGNAL nor_790_nl : STD_LOGIC;
  SIGNAL nor_791_nl : STD_LOGIC;
  SIGNAL mux_2575_nl : STD_LOGIC;
  SIGNAL nand_410_nl : STD_LOGIC;
  SIGNAL mux_2574_nl : STD_LOGIC;
  SIGNAL mux_2573_nl : STD_LOGIC;
  SIGNAL mux_2572_nl : STD_LOGIC;
  SIGNAL nor_783_nl : STD_LOGIC;
  SIGNAL nor_784_nl : STD_LOGIC;
  SIGNAL mux_2571_nl : STD_LOGIC;
  SIGNAL and_557_nl : STD_LOGIC;
  SIGNAL and_558_nl : STD_LOGIC;
  SIGNAL mux_2570_nl : STD_LOGIC;
  SIGNAL mux_2569_nl : STD_LOGIC;
  SIGNAL and_814_nl : STD_LOGIC;
  SIGNAL and_821_nl : STD_LOGIC;
  SIGNAL mux_2568_nl : STD_LOGIC;
  SIGNAL nor_787_nl : STD_LOGIC;
  SIGNAL nor_788_nl : STD_LOGIC;
  SIGNAL or_4083_nl : STD_LOGIC;
  SIGNAL mux_2567_nl : STD_LOGIC;
  SIGNAL mux_2566_nl : STD_LOGIC;
  SIGNAL mux_2565_nl : STD_LOGIC;
  SIGNAL or_3208_nl : STD_LOGIC;
  SIGNAL mux_2564_nl : STD_LOGIC;
  SIGNAL nand_247_nl : STD_LOGIC;
  SIGNAL mux_2563_nl : STD_LOGIC;
  SIGNAL mux_2562_nl : STD_LOGIC;
  SIGNAL nand_475_nl : STD_LOGIC;
  SIGNAL mux_2561_nl : STD_LOGIC;
  SIGNAL or_3200_nl : STD_LOGIC;
  SIGNAL mux_2590_nl : STD_LOGIC;
  SIGNAL mux_2589_nl : STD_LOGIC;
  SIGNAL or_3242_nl : STD_LOGIC;
  SIGNAL mux_2588_nl : STD_LOGIC;
  SIGNAL or_3241_nl : STD_LOGIC;
  SIGNAL or_3240_nl : STD_LOGIC;
  SIGNAL mux_2587_nl : STD_LOGIC;
  SIGNAL mux_2586_nl : STD_LOGIC;
  SIGNAL mux_2585_nl : STD_LOGIC;
  SIGNAL or_3238_nl : STD_LOGIC;
  SIGNAL mux_2584_nl : STD_LOGIC;
  SIGNAL nand_238_nl : STD_LOGIC;
  SIGNAL mux_2583_nl : STD_LOGIC;
  SIGNAL mux_2582_nl : STD_LOGIC;
  SIGNAL nand_398_nl : STD_LOGIC;
  SIGNAL mux_2581_nl : STD_LOGIC;
  SIGNAL or_3233_nl : STD_LOGIC;
  SIGNAL or_3232_nl : STD_LOGIC;
  SIGNAL mux_2580_nl : STD_LOGIC;
  SIGNAL mux_2579_nl : STD_LOGIC;
  SIGNAL mux_2578_nl : STD_LOGIC;
  SIGNAL or_3231_nl : STD_LOGIC;
  SIGNAL or_3229_nl : STD_LOGIC;
  SIGNAL mux_2577_nl : STD_LOGIC;
  SIGNAL nand_242_nl : STD_LOGIC;
  SIGNAL nand_243_nl : STD_LOGIC;
  SIGNAL nand_133_nl : STD_LOGIC;
  SIGNAL mux_2576_nl : STD_LOGIC;
  SIGNAL nor_781_nl : STD_LOGIC;
  SIGNAL nor_782_nl : STD_LOGIC;
  SIGNAL mux_2605_nl : STD_LOGIC;
  SIGNAL nand_409_nl : STD_LOGIC;
  SIGNAL mux_2604_nl : STD_LOGIC;
  SIGNAL mux_2603_nl : STD_LOGIC;
  SIGNAL mux_2602_nl : STD_LOGIC;
  SIGNAL nor_773_nl : STD_LOGIC;
  SIGNAL and_555_nl : STD_LOGIC;
  SIGNAL mux_2601_nl : STD_LOGIC;
  SIGNAL nor_774_nl : STD_LOGIC;
  SIGNAL nor_775_nl : STD_LOGIC;
  SIGNAL mux_2600_nl : STD_LOGIC;
  SIGNAL mux_2599_nl : STD_LOGIC;
  SIGNAL nor_776_nl : STD_LOGIC;
  SIGNAL nor_777_nl : STD_LOGIC;
  SIGNAL mux_2598_nl : STD_LOGIC;
  SIGNAL nor_778_nl : STD_LOGIC;
  SIGNAL nor_779_nl : STD_LOGIC;
  SIGNAL or_4082_nl : STD_LOGIC;
  SIGNAL mux_2597_nl : STD_LOGIC;
  SIGNAL mux_2596_nl : STD_LOGIC;
  SIGNAL mux_2595_nl : STD_LOGIC;
  SIGNAL or_3252_nl : STD_LOGIC;
  SIGNAL mux_2594_nl : STD_LOGIC;
  SIGNAL or_3249_nl : STD_LOGIC;
  SIGNAL mux_2593_nl : STD_LOGIC;
  SIGNAL mux_2592_nl : STD_LOGIC;
  SIGNAL or_3246_nl : STD_LOGIC;
  SIGNAL mux_2591_nl : STD_LOGIC;
  SIGNAL or_3243_nl : STD_LOGIC;
  SIGNAL mux_2620_nl : STD_LOGIC;
  SIGNAL mux_2619_nl : STD_LOGIC;
  SIGNAL or_3286_nl : STD_LOGIC;
  SIGNAL mux_2618_nl : STD_LOGIC;
  SIGNAL or_3285_nl : STD_LOGIC;
  SIGNAL or_3284_nl : STD_LOGIC;
  SIGNAL mux_2617_nl : STD_LOGIC;
  SIGNAL mux_2616_nl : STD_LOGIC;
  SIGNAL mux_2615_nl : STD_LOGIC;
  SIGNAL or_3282_nl : STD_LOGIC;
  SIGNAL mux_2614_nl : STD_LOGIC;
  SIGNAL or_3280_nl : STD_LOGIC;
  SIGNAL mux_2613_nl : STD_LOGIC;
  SIGNAL mux_2612_nl : STD_LOGIC;
  SIGNAL or_3279_nl : STD_LOGIC;
  SIGNAL mux_2611_nl : STD_LOGIC;
  SIGNAL or_3277_nl : STD_LOGIC;
  SIGNAL or_3276_nl : STD_LOGIC;
  SIGNAL mux_2610_nl : STD_LOGIC;
  SIGNAL mux_2609_nl : STD_LOGIC;
  SIGNAL mux_2608_nl : STD_LOGIC;
  SIGNAL nand_237_nl : STD_LOGIC;
  SIGNAL or_3273_nl : STD_LOGIC;
  SIGNAL mux_2607_nl : STD_LOGIC;
  SIGNAL or_3271_nl : STD_LOGIC;
  SIGNAL or_3270_nl : STD_LOGIC;
  SIGNAL nand_135_nl : STD_LOGIC;
  SIGNAL mux_2606_nl : STD_LOGIC;
  SIGNAL nor_771_nl : STD_LOGIC;
  SIGNAL nor_772_nl : STD_LOGIC;
  SIGNAL mux_2635_nl : STD_LOGIC;
  SIGNAL nand_408_nl : STD_LOGIC;
  SIGNAL mux_2634_nl : STD_LOGIC;
  SIGNAL mux_2633_nl : STD_LOGIC;
  SIGNAL mux_2632_nl : STD_LOGIC;
  SIGNAL nor_764_nl : STD_LOGIC;
  SIGNAL nor_765_nl : STD_LOGIC;
  SIGNAL mux_2631_nl : STD_LOGIC;
  SIGNAL and_552_nl : STD_LOGIC;
  SIGNAL and_553_nl : STD_LOGIC;
  SIGNAL mux_2630_nl : STD_LOGIC;
  SIGNAL mux_2629_nl : STD_LOGIC;
  SIGNAL and_815_nl : STD_LOGIC;
  SIGNAL and_822_nl : STD_LOGIC;
  SIGNAL mux_2628_nl : STD_LOGIC;
  SIGNAL nor_768_nl : STD_LOGIC;
  SIGNAL nor_769_nl : STD_LOGIC;
  SIGNAL or_4081_nl : STD_LOGIC;
  SIGNAL mux_2627_nl : STD_LOGIC;
  SIGNAL mux_2626_nl : STD_LOGIC;
  SIGNAL mux_2625_nl : STD_LOGIC;
  SIGNAL or_3296_nl : STD_LOGIC;
  SIGNAL mux_2624_nl : STD_LOGIC;
  SIGNAL nand_232_nl : STD_LOGIC;
  SIGNAL mux_2623_nl : STD_LOGIC;
  SIGNAL mux_2622_nl : STD_LOGIC;
  SIGNAL nand_474_nl : STD_LOGIC;
  SIGNAL mux_2621_nl : STD_LOGIC;
  SIGNAL or_3287_nl : STD_LOGIC;
  SIGNAL mux_2650_nl : STD_LOGIC;
  SIGNAL mux_2649_nl : STD_LOGIC;
  SIGNAL or_3329_nl : STD_LOGIC;
  SIGNAL mux_2648_nl : STD_LOGIC;
  SIGNAL or_3328_nl : STD_LOGIC;
  SIGNAL or_3327_nl : STD_LOGIC;
  SIGNAL mux_2647_nl : STD_LOGIC;
  SIGNAL mux_2646_nl : STD_LOGIC;
  SIGNAL mux_2645_nl : STD_LOGIC;
  SIGNAL or_3325_nl : STD_LOGIC;
  SIGNAL mux_2644_nl : STD_LOGIC;
  SIGNAL nand_223_nl : STD_LOGIC;
  SIGNAL mux_2643_nl : STD_LOGIC;
  SIGNAL mux_2642_nl : STD_LOGIC;
  SIGNAL nand_396_nl : STD_LOGIC;
  SIGNAL mux_2641_nl : STD_LOGIC;
  SIGNAL or_3320_nl : STD_LOGIC;
  SIGNAL or_3319_nl : STD_LOGIC;
  SIGNAL mux_2640_nl : STD_LOGIC;
  SIGNAL mux_2639_nl : STD_LOGIC;
  SIGNAL mux_2638_nl : STD_LOGIC;
  SIGNAL or_3318_nl : STD_LOGIC;
  SIGNAL or_3316_nl : STD_LOGIC;
  SIGNAL mux_2637_nl : STD_LOGIC;
  SIGNAL nand_227_nl : STD_LOGIC;
  SIGNAL nand_228_nl : STD_LOGIC;
  SIGNAL nand_137_nl : STD_LOGIC;
  SIGNAL mux_2636_nl : STD_LOGIC;
  SIGNAL nor_762_nl : STD_LOGIC;
  SIGNAL nor_763_nl : STD_LOGIC;
  SIGNAL mux_2665_nl : STD_LOGIC;
  SIGNAL nand_407_nl : STD_LOGIC;
  SIGNAL mux_2664_nl : STD_LOGIC;
  SIGNAL mux_2663_nl : STD_LOGIC;
  SIGNAL mux_2662_nl : STD_LOGIC;
  SIGNAL nor_756_nl : STD_LOGIC;
  SIGNAL and_548_nl : STD_LOGIC;
  SIGNAL mux_2661_nl : STD_LOGIC;
  SIGNAL and_549_nl : STD_LOGIC;
  SIGNAL and_550_nl : STD_LOGIC;
  SIGNAL mux_2660_nl : STD_LOGIC;
  SIGNAL mux_2659_nl : STD_LOGIC;
  SIGNAL and_816_nl : STD_LOGIC;
  SIGNAL and_823_nl : STD_LOGIC;
  SIGNAL mux_2658_nl : STD_LOGIC;
  SIGNAL nor_759_nl : STD_LOGIC;
  SIGNAL nor_760_nl : STD_LOGIC;
  SIGNAL or_4080_nl : STD_LOGIC;
  SIGNAL mux_2657_nl : STD_LOGIC;
  SIGNAL mux_2656_nl : STD_LOGIC;
  SIGNAL mux_2655_nl : STD_LOGIC;
  SIGNAL or_3339_nl : STD_LOGIC;
  SIGNAL mux_2654_nl : STD_LOGIC;
  SIGNAL nand_218_nl : STD_LOGIC;
  SIGNAL mux_2653_nl : STD_LOGIC;
  SIGNAL mux_2652_nl : STD_LOGIC;
  SIGNAL nand_473_nl : STD_LOGIC;
  SIGNAL mux_2651_nl : STD_LOGIC;
  SIGNAL or_3330_nl : STD_LOGIC;
  SIGNAL mux_2680_nl : STD_LOGIC;
  SIGNAL mux_2679_nl : STD_LOGIC;
  SIGNAL or_3372_nl : STD_LOGIC;
  SIGNAL mux_2678_nl : STD_LOGIC;
  SIGNAL or_3371_nl : STD_LOGIC;
  SIGNAL or_3370_nl : STD_LOGIC;
  SIGNAL mux_2677_nl : STD_LOGIC;
  SIGNAL mux_2676_nl : STD_LOGIC;
  SIGNAL mux_2675_nl : STD_LOGIC;
  SIGNAL or_3368_nl : STD_LOGIC;
  SIGNAL mux_2674_nl : STD_LOGIC;
  SIGNAL nand_210_nl : STD_LOGIC;
  SIGNAL mux_2673_nl : STD_LOGIC;
  SIGNAL mux_2672_nl : STD_LOGIC;
  SIGNAL nand_394_nl : STD_LOGIC;
  SIGNAL mux_2671_nl : STD_LOGIC;
  SIGNAL or_3363_nl : STD_LOGIC;
  SIGNAL or_3362_nl : STD_LOGIC;
  SIGNAL mux_2670_nl : STD_LOGIC;
  SIGNAL mux_2669_nl : STD_LOGIC;
  SIGNAL mux_2668_nl : STD_LOGIC;
  SIGNAL nand_212_nl : STD_LOGIC;
  SIGNAL or_3359_nl : STD_LOGIC;
  SIGNAL mux_2667_nl : STD_LOGIC;
  SIGNAL nand_213_nl : STD_LOGIC;
  SIGNAL nand_214_nl : STD_LOGIC;
  SIGNAL nand_139_nl : STD_LOGIC;
  SIGNAL mux_2666_nl : STD_LOGIC;
  SIGNAL nor_754_nl : STD_LOGIC;
  SIGNAL nor_755_nl : STD_LOGIC;
  SIGNAL mux_2695_nl : STD_LOGIC;
  SIGNAL nand_406_nl : STD_LOGIC;
  SIGNAL mux_2694_nl : STD_LOGIC;
  SIGNAL mux_2693_nl : STD_LOGIC;
  SIGNAL mux_2692_nl : STD_LOGIC;
  SIGNAL and_539_nl : STD_LOGIC;
  SIGNAL and_540_nl : STD_LOGIC;
  SIGNAL mux_2691_nl : STD_LOGIC;
  SIGNAL and_541_nl : STD_LOGIC;
  SIGNAL and_542_nl : STD_LOGIC;
  SIGNAL mux_2690_nl : STD_LOGIC;
  SIGNAL mux_2689_nl : STD_LOGIC;
  SIGNAL and_817_nl : STD_LOGIC;
  SIGNAL and_824_nl : STD_LOGIC;
  SIGNAL mux_2688_nl : STD_LOGIC;
  SIGNAL and_543_nl : STD_LOGIC;
  SIGNAL and_544_nl : STD_LOGIC;
  SIGNAL or_4079_nl : STD_LOGIC;
  SIGNAL mux_2687_nl : STD_LOGIC;
  SIGNAL mux_2686_nl : STD_LOGIC;
  SIGNAL mux_2685_nl : STD_LOGIC;
  SIGNAL mux_2684_nl : STD_LOGIC;
  SIGNAL nand_203_nl : STD_LOGIC;
  SIGNAL mux_2683_nl : STD_LOGIC;
  SIGNAL mux_2682_nl : STD_LOGIC;
  SIGNAL nand_nl : STD_LOGIC;
  SIGNAL mux_2681_nl : STD_LOGIC;
  SIGNAL nand_205_nl : STD_LOGIC;
  SIGNAL mux_2710_nl : STD_LOGIC;
  SIGNAL mux_2709_nl : STD_LOGIC;
  SIGNAL or_3405_nl : STD_LOGIC;
  SIGNAL mux_2708_nl : STD_LOGIC;
  SIGNAL nand_192_nl : STD_LOGIC;
  SIGNAL nand_193_nl : STD_LOGIC;
  SIGNAL mux_2707_nl : STD_LOGIC;
  SIGNAL mux_2706_nl : STD_LOGIC;
  SIGNAL mux_2705_nl : STD_LOGIC;
  SIGNAL and_535_nl : STD_LOGIC;
  SIGNAL mux_2704_nl : STD_LOGIC;
  SIGNAL nand_194_nl : STD_LOGIC;
  SIGNAL mux_2703_nl : STD_LOGIC;
  SIGNAL mux_2702_nl : STD_LOGIC;
  SIGNAL nand_392_nl : STD_LOGIC;
  SIGNAL mux_2701_nl : STD_LOGIC;
  SIGNAL nand_196_nl : STD_LOGIC;
  SIGNAL or_3396_nl : STD_LOGIC;
  SIGNAL mux_2700_nl : STD_LOGIC;
  SIGNAL mux_2699_nl : STD_LOGIC;
  SIGNAL mux_2698_nl : STD_LOGIC;
  SIGNAL or_4002_nl : STD_LOGIC;
  SIGNAL nand_198_nl : STD_LOGIC;
  SIGNAL mux_2697_nl : STD_LOGIC;
  SIGNAL nand_199_nl : STD_LOGIC;
  SIGNAL nand_200_nl : STD_LOGIC;
  SIGNAL nand_141_nl : STD_LOGIC;
  SIGNAL mux_2696_nl : STD_LOGIC;
  SIGNAL and_536_nl : STD_LOGIC;
  SIGNAL and_537_nl : STD_LOGIC;
  SIGNAL mux_2717_nl : STD_LOGIC;
  SIGNAL mux_2716_nl : STD_LOGIC;
  SIGNAL mux_2715_nl : STD_LOGIC;
  SIGNAL nor_743_nl : STD_LOGIC;
  SIGNAL nor_744_nl : STD_LOGIC;
  SIGNAL mux_2714_nl : STD_LOGIC;
  SIGNAL nor_745_nl : STD_LOGIC;
  SIGNAL mux_2713_nl : STD_LOGIC;
  SIGNAL mux_2712_nl : STD_LOGIC;
  SIGNAL nor_747_nl : STD_LOGIC;
  SIGNAL mux_2711_nl : STD_LOGIC;
  SIGNAL nor_749_nl : STD_LOGIC;
  SIGNAL nor_750_nl : STD_LOGIC;
  SIGNAL mux_2720_nl : STD_LOGIC;
  SIGNAL mux_2719_nl : STD_LOGIC;
  SIGNAL nor_739_nl : STD_LOGIC;
  SIGNAL mux_2718_nl : STD_LOGIC;
  SIGNAL nor_742_nl : STD_LOGIC;
  SIGNAL mux_2725_nl : STD_LOGIC;
  SIGNAL mux_2724_nl : STD_LOGIC;
  SIGNAL nor_733_nl : STD_LOGIC;
  SIGNAL mux_2723_nl : STD_LOGIC;
  SIGNAL mux_2722_nl : STD_LOGIC;
  SIGNAL nor_736_nl : STD_LOGIC;
  SIGNAL mux_2721_nl : STD_LOGIC;
  SIGNAL mux_2728_nl : STD_LOGIC;
  SIGNAL mux_2727_nl : STD_LOGIC;
  SIGNAL nor_729_nl : STD_LOGIC;
  SIGNAL mux_2726_nl : STD_LOGIC;
  SIGNAL nor_732_nl : STD_LOGIC;
  SIGNAL mux_2734_nl : STD_LOGIC;
  SIGNAL mux_2733_nl : STD_LOGIC;
  SIGNAL mux_2732_nl : STD_LOGIC;
  SIGNAL nor_722_nl : STD_LOGIC;
  SIGNAL nor_723_nl : STD_LOGIC;
  SIGNAL mux_2731_nl : STD_LOGIC;
  SIGNAL nor_724_nl : STD_LOGIC;
  SIGNAL nor_725_nl : STD_LOGIC;
  SIGNAL mux_2730_nl : STD_LOGIC;
  SIGNAL nor_726_nl : STD_LOGIC;
  SIGNAL mux_2729_nl : STD_LOGIC;
  SIGNAL nor_727_nl : STD_LOGIC;
  SIGNAL nor_728_nl : STD_LOGIC;
  SIGNAL mux_2737_nl : STD_LOGIC;
  SIGNAL mux_2736_nl : STD_LOGIC;
  SIGNAL nor_718_nl : STD_LOGIC;
  SIGNAL mux_2735_nl : STD_LOGIC;
  SIGNAL nor_721_nl : STD_LOGIC;
  SIGNAL mux_2742_nl : STD_LOGIC;
  SIGNAL mux_2741_nl : STD_LOGIC;
  SIGNAL nor_712_nl : STD_LOGIC;
  SIGNAL mux_2740_nl : STD_LOGIC;
  SIGNAL mux_2739_nl : STD_LOGIC;
  SIGNAL nor_715_nl : STD_LOGIC;
  SIGNAL mux_2738_nl : STD_LOGIC;
  SIGNAL mux_2745_nl : STD_LOGIC;
  SIGNAL mux_2744_nl : STD_LOGIC;
  SIGNAL nor_708_nl : STD_LOGIC;
  SIGNAL mux_2743_nl : STD_LOGIC;
  SIGNAL nor_711_nl : STD_LOGIC;
  SIGNAL mux_2752_nl : STD_LOGIC;
  SIGNAL mux_2751_nl : STD_LOGIC;
  SIGNAL mux_2750_nl : STD_LOGIC;
  SIGNAL nor_700_nl : STD_LOGIC;
  SIGNAL nor_701_nl : STD_LOGIC;
  SIGNAL mux_2749_nl : STD_LOGIC;
  SIGNAL nor_702_nl : STD_LOGIC;
  SIGNAL mux_2748_nl : STD_LOGIC;
  SIGNAL mux_2747_nl : STD_LOGIC;
  SIGNAL nor_704_nl : STD_LOGIC;
  SIGNAL mux_2746_nl : STD_LOGIC;
  SIGNAL nor_706_nl : STD_LOGIC;
  SIGNAL nor_707_nl : STD_LOGIC;
  SIGNAL mux_2755_nl : STD_LOGIC;
  SIGNAL mux_2754_nl : STD_LOGIC;
  SIGNAL nor_696_nl : STD_LOGIC;
  SIGNAL mux_2753_nl : STD_LOGIC;
  SIGNAL nor_699_nl : STD_LOGIC;
  SIGNAL mux_2760_nl : STD_LOGIC;
  SIGNAL mux_2759_nl : STD_LOGIC;
  SIGNAL nor_690_nl : STD_LOGIC;
  SIGNAL mux_2758_nl : STD_LOGIC;
  SIGNAL mux_2757_nl : STD_LOGIC;
  SIGNAL nor_693_nl : STD_LOGIC;
  SIGNAL mux_2756_nl : STD_LOGIC;
  SIGNAL mux_2763_nl : STD_LOGIC;
  SIGNAL mux_2762_nl : STD_LOGIC;
  SIGNAL nor_686_nl : STD_LOGIC;
  SIGNAL mux_2761_nl : STD_LOGIC;
  SIGNAL nor_689_nl : STD_LOGIC;
  SIGNAL mux_2769_nl : STD_LOGIC;
  SIGNAL mux_2768_nl : STD_LOGIC;
  SIGNAL mux_2767_nl : STD_LOGIC;
  SIGNAL nor_679_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL mux_2766_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL nor_682_nl : STD_LOGIC;
  SIGNAL mux_2765_nl : STD_LOGIC;
  SIGNAL nor_683_nl : STD_LOGIC;
  SIGNAL mux_2764_nl : STD_LOGIC;
  SIGNAL nor_684_nl : STD_LOGIC;
  SIGNAL nor_685_nl : STD_LOGIC;
  SIGNAL mux_2772_nl : STD_LOGIC;
  SIGNAL mux_2771_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL mux_2770_nl : STD_LOGIC;
  SIGNAL nor_678_nl : STD_LOGIC;
  SIGNAL mux_2777_nl : STD_LOGIC;
  SIGNAL mux_2776_nl : STD_LOGIC;
  SIGNAL nor_669_nl : STD_LOGIC;
  SIGNAL mux_2775_nl : STD_LOGIC;
  SIGNAL mux_2774_nl : STD_LOGIC;
  SIGNAL nor_672_nl : STD_LOGIC;
  SIGNAL mux_2773_nl : STD_LOGIC;
  SIGNAL mux_2780_nl : STD_LOGIC;
  SIGNAL mux_2779_nl : STD_LOGIC;
  SIGNAL nor_665_nl : STD_LOGIC;
  SIGNAL mux_2778_nl : STD_LOGIC;
  SIGNAL nor_668_nl : STD_LOGIC;
  SIGNAL mux_2787_nl : STD_LOGIC;
  SIGNAL mux_2786_nl : STD_LOGIC;
  SIGNAL mux_2785_nl : STD_LOGIC;
  SIGNAL nor_657_nl : STD_LOGIC;
  SIGNAL nor_658_nl : STD_LOGIC;
  SIGNAL mux_2784_nl : STD_LOGIC;
  SIGNAL nor_659_nl : STD_LOGIC;
  SIGNAL mux_2783_nl : STD_LOGIC;
  SIGNAL mux_2782_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL mux_2781_nl : STD_LOGIC;
  SIGNAL nor_663_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL mux_2790_nl : STD_LOGIC;
  SIGNAL mux_2789_nl : STD_LOGIC;
  SIGNAL nor_653_nl : STD_LOGIC;
  SIGNAL mux_2788_nl : STD_LOGIC;
  SIGNAL nor_656_nl : STD_LOGIC;
  SIGNAL mux_2795_nl : STD_LOGIC;
  SIGNAL mux_2794_nl : STD_LOGIC;
  SIGNAL nor_647_nl : STD_LOGIC;
  SIGNAL mux_2793_nl : STD_LOGIC;
  SIGNAL mux_2792_nl : STD_LOGIC;
  SIGNAL nor_650_nl : STD_LOGIC;
  SIGNAL mux_2791_nl : STD_LOGIC;
  SIGNAL mux_2798_nl : STD_LOGIC;
  SIGNAL mux_2797_nl : STD_LOGIC;
  SIGNAL nor_643_nl : STD_LOGIC;
  SIGNAL mux_2796_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL mux_2804_nl : STD_LOGIC;
  SIGNAL mux_2803_nl : STD_LOGIC;
  SIGNAL mux_2802_nl : STD_LOGIC;
  SIGNAL nor_636_nl : STD_LOGIC;
  SIGNAL nor_637_nl : STD_LOGIC;
  SIGNAL mux_2801_nl : STD_LOGIC;
  SIGNAL nor_638_nl : STD_LOGIC;
  SIGNAL nor_639_nl : STD_LOGIC;
  SIGNAL mux_2800_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL mux_2799_nl : STD_LOGIC;
  SIGNAL nor_641_nl : STD_LOGIC;
  SIGNAL nor_642_nl : STD_LOGIC;
  SIGNAL mux_2807_nl : STD_LOGIC;
  SIGNAL mux_2806_nl : STD_LOGIC;
  SIGNAL nor_632_nl : STD_LOGIC;
  SIGNAL mux_2805_nl : STD_LOGIC;
  SIGNAL nor_635_nl : STD_LOGIC;
  SIGNAL mux_2812_nl : STD_LOGIC;
  SIGNAL mux_2811_nl : STD_LOGIC;
  SIGNAL nor_626_nl : STD_LOGIC;
  SIGNAL mux_2810_nl : STD_LOGIC;
  SIGNAL mux_2809_nl : STD_LOGIC;
  SIGNAL nor_629_nl : STD_LOGIC;
  SIGNAL mux_2808_nl : STD_LOGIC;
  SIGNAL mux_2815_nl : STD_LOGIC;
  SIGNAL mux_2814_nl : STD_LOGIC;
  SIGNAL nor_622_nl : STD_LOGIC;
  SIGNAL mux_2813_nl : STD_LOGIC;
  SIGNAL nor_625_nl : STD_LOGIC;
  SIGNAL mux_2822_nl : STD_LOGIC;
  SIGNAL mux_2821_nl : STD_LOGIC;
  SIGNAL mux_2820_nl : STD_LOGIC;
  SIGNAL nor_614_nl : STD_LOGIC;
  SIGNAL nor_615_nl : STD_LOGIC;
  SIGNAL mux_2819_nl : STD_LOGIC;
  SIGNAL nor_616_nl : STD_LOGIC;
  SIGNAL mux_2818_nl : STD_LOGIC;
  SIGNAL mux_2817_nl : STD_LOGIC;
  SIGNAL nor_618_nl : STD_LOGIC;
  SIGNAL mux_2816_nl : STD_LOGIC;
  SIGNAL nor_620_nl : STD_LOGIC;
  SIGNAL nor_621_nl : STD_LOGIC;
  SIGNAL mux_2825_nl : STD_LOGIC;
  SIGNAL mux_2824_nl : STD_LOGIC;
  SIGNAL nor_610_nl : STD_LOGIC;
  SIGNAL mux_2823_nl : STD_LOGIC;
  SIGNAL nor_613_nl : STD_LOGIC;
  SIGNAL mux_2830_nl : STD_LOGIC;
  SIGNAL mux_2829_nl : STD_LOGIC;
  SIGNAL nor_604_nl : STD_LOGIC;
  SIGNAL mux_2828_nl : STD_LOGIC;
  SIGNAL mux_2827_nl : STD_LOGIC;
  SIGNAL nor_607_nl : STD_LOGIC;
  SIGNAL mux_2826_nl : STD_LOGIC;
  SIGNAL mux_2833_nl : STD_LOGIC;
  SIGNAL mux_2832_nl : STD_LOGIC;
  SIGNAL nor_600_nl : STD_LOGIC;
  SIGNAL mux_2831_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL mux_2839_nl : STD_LOGIC;
  SIGNAL mux_2838_nl : STD_LOGIC;
  SIGNAL mux_2837_nl : STD_LOGIC;
  SIGNAL nor_593_nl : STD_LOGIC;
  SIGNAL nor_594_nl : STD_LOGIC;
  SIGNAL mux_2836_nl : STD_LOGIC;
  SIGNAL nor_595_nl : STD_LOGIC;
  SIGNAL nor_596_nl : STD_LOGIC;
  SIGNAL mux_2835_nl : STD_LOGIC;
  SIGNAL nor_597_nl : STD_LOGIC;
  SIGNAL mux_2834_nl : STD_LOGIC;
  SIGNAL nor_598_nl : STD_LOGIC;
  SIGNAL nor_599_nl : STD_LOGIC;
  SIGNAL mux_2842_nl : STD_LOGIC;
  SIGNAL mux_2841_nl : STD_LOGIC;
  SIGNAL nor_589_nl : STD_LOGIC;
  SIGNAL mux_2840_nl : STD_LOGIC;
  SIGNAL nor_592_nl : STD_LOGIC;
  SIGNAL mux_2847_nl : STD_LOGIC;
  SIGNAL mux_2846_nl : STD_LOGIC;
  SIGNAL nor_583_nl : STD_LOGIC;
  SIGNAL mux_2845_nl : STD_LOGIC;
  SIGNAL mux_2844_nl : STD_LOGIC;
  SIGNAL nor_586_nl : STD_LOGIC;
  SIGNAL mux_2843_nl : STD_LOGIC;
  SIGNAL mux_2850_nl : STD_LOGIC;
  SIGNAL mux_2849_nl : STD_LOGIC;
  SIGNAL nor_581_nl : STD_LOGIC;
  SIGNAL mux_2848_nl : STD_LOGIC;
  SIGNAL nor_582_nl : STD_LOGIC;
  SIGNAL mux_2857_nl : STD_LOGIC;
  SIGNAL mux_2856_nl : STD_LOGIC;
  SIGNAL mux_2855_nl : STD_LOGIC;
  SIGNAL nor_573_nl : STD_LOGIC;
  SIGNAL nor_574_nl : STD_LOGIC;
  SIGNAL mux_2854_nl : STD_LOGIC;
  SIGNAL nor_575_nl : STD_LOGIC;
  SIGNAL mux_2853_nl : STD_LOGIC;
  SIGNAL mux_2852_nl : STD_LOGIC;
  SIGNAL nor_577_nl : STD_LOGIC;
  SIGNAL mux_2851_nl : STD_LOGIC;
  SIGNAL nor_579_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL mux_2860_nl : STD_LOGIC;
  SIGNAL mux_2859_nl : STD_LOGIC;
  SIGNAL nor_569_nl : STD_LOGIC;
  SIGNAL mux_2858_nl : STD_LOGIC;
  SIGNAL nor_572_nl : STD_LOGIC;
  SIGNAL mux_2865_nl : STD_LOGIC;
  SIGNAL mux_2864_nl : STD_LOGIC;
  SIGNAL nor_563_nl : STD_LOGIC;
  SIGNAL mux_2863_nl : STD_LOGIC;
  SIGNAL mux_2862_nl : STD_LOGIC;
  SIGNAL nor_566_nl : STD_LOGIC;
  SIGNAL mux_2861_nl : STD_LOGIC;
  SIGNAL mux_2868_nl : STD_LOGIC;
  SIGNAL mux_2867_nl : STD_LOGIC;
  SIGNAL nor_559_nl : STD_LOGIC;
  SIGNAL mux_2866_nl : STD_LOGIC;
  SIGNAL nor_562_nl : STD_LOGIC;
  SIGNAL mux_2874_nl : STD_LOGIC;
  SIGNAL mux_2873_nl : STD_LOGIC;
  SIGNAL mux_2872_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL nor_553_nl : STD_LOGIC;
  SIGNAL mux_2871_nl : STD_LOGIC;
  SIGNAL nor_554_nl : STD_LOGIC;
  SIGNAL nor_555_nl : STD_LOGIC;
  SIGNAL mux_2870_nl : STD_LOGIC;
  SIGNAL nor_556_nl : STD_LOGIC;
  SIGNAL mux_2869_nl : STD_LOGIC;
  SIGNAL nor_557_nl : STD_LOGIC;
  SIGNAL nor_558_nl : STD_LOGIC;
  SIGNAL mux_2877_nl : STD_LOGIC;
  SIGNAL mux_2876_nl : STD_LOGIC;
  SIGNAL nor_548_nl : STD_LOGIC;
  SIGNAL mux_2875_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL mux_2882_nl : STD_LOGIC;
  SIGNAL mux_2881_nl : STD_LOGIC;
  SIGNAL nor_542_nl : STD_LOGIC;
  SIGNAL mux_2880_nl : STD_LOGIC;
  SIGNAL mux_2879_nl : STD_LOGIC;
  SIGNAL nor_545_nl : STD_LOGIC;
  SIGNAL mux_2878_nl : STD_LOGIC;
  SIGNAL mux_2885_nl : STD_LOGIC;
  SIGNAL mux_2884_nl : STD_LOGIC;
  SIGNAL nor_538_nl : STD_LOGIC;
  SIGNAL mux_2883_nl : STD_LOGIC;
  SIGNAL nor_541_nl : STD_LOGIC;
  SIGNAL mux_2892_nl : STD_LOGIC;
  SIGNAL mux_2891_nl : STD_LOGIC;
  SIGNAL mux_2890_nl : STD_LOGIC;
  SIGNAL nor_530_nl : STD_LOGIC;
  SIGNAL nor_531_nl : STD_LOGIC;
  SIGNAL mux_2889_nl : STD_LOGIC;
  SIGNAL nor_532_nl : STD_LOGIC;
  SIGNAL mux_2888_nl : STD_LOGIC;
  SIGNAL mux_2887_nl : STD_LOGIC;
  SIGNAL nor_534_nl : STD_LOGIC;
  SIGNAL mux_2886_nl : STD_LOGIC;
  SIGNAL nor_536_nl : STD_LOGIC;
  SIGNAL nor_537_nl : STD_LOGIC;
  SIGNAL mux_2895_nl : STD_LOGIC;
  SIGNAL mux_2894_nl : STD_LOGIC;
  SIGNAL nor_526_nl : STD_LOGIC;
  SIGNAL mux_2893_nl : STD_LOGIC;
  SIGNAL nor_529_nl : STD_LOGIC;
  SIGNAL mux_2900_nl : STD_LOGIC;
  SIGNAL mux_2899_nl : STD_LOGIC;
  SIGNAL nor_520_nl : STD_LOGIC;
  SIGNAL mux_2898_nl : STD_LOGIC;
  SIGNAL mux_2897_nl : STD_LOGIC;
  SIGNAL nor_523_nl : STD_LOGIC;
  SIGNAL mux_2896_nl : STD_LOGIC;
  SIGNAL mux_2903_nl : STD_LOGIC;
  SIGNAL mux_2902_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL mux_2901_nl : STD_LOGIC;
  SIGNAL nor_519_nl : STD_LOGIC;
  SIGNAL mux_2909_nl : STD_LOGIC;
  SIGNAL mux_2908_nl : STD_LOGIC;
  SIGNAL mux_2907_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL mux_2906_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL nor_512_nl : STD_LOGIC;
  SIGNAL mux_2905_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL mux_2904_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL mux_2912_nl : STD_LOGIC;
  SIGNAL mux_2911_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL mux_2910_nl : STD_LOGIC;
  SIGNAL nor_508_nl : STD_LOGIC;
  SIGNAL mux_2917_nl : STD_LOGIC;
  SIGNAL mux_2916_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL mux_2915_nl : STD_LOGIC;
  SIGNAL mux_2914_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL mux_2913_nl : STD_LOGIC;
  SIGNAL mux_2920_nl : STD_LOGIC;
  SIGNAL mux_2919_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL mux_2918_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL mux_2927_nl : STD_LOGIC;
  SIGNAL mux_2926_nl : STD_LOGIC;
  SIGNAL mux_2925_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL mux_2924_nl : STD_LOGIC;
  SIGNAL nor_491_nl : STD_LOGIC;
  SIGNAL mux_2923_nl : STD_LOGIC;
  SIGNAL mux_2922_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL mux_2921_nl : STD_LOGIC;
  SIGNAL nor_495_nl : STD_LOGIC;
  SIGNAL nor_496_nl : STD_LOGIC;
  SIGNAL mux_2930_nl : STD_LOGIC;
  SIGNAL mux_2929_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL mux_2928_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL mux_2935_nl : STD_LOGIC;
  SIGNAL mux_2934_nl : STD_LOGIC;
  SIGNAL nor_479_nl : STD_LOGIC;
  SIGNAL mux_2933_nl : STD_LOGIC;
  SIGNAL mux_2932_nl : STD_LOGIC;
  SIGNAL nor_482_nl : STD_LOGIC;
  SIGNAL mux_2931_nl : STD_LOGIC;
  SIGNAL mux_2938_nl : STD_LOGIC;
  SIGNAL mux_2937_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL mux_2936_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL mux_2944_nl : STD_LOGIC;
  SIGNAL mux_2943_nl : STD_LOGIC;
  SIGNAL mux_2942_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL mux_2941_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL nor_471_nl : STD_LOGIC;
  SIGNAL mux_2940_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL mux_2939_nl : STD_LOGIC;
  SIGNAL nor_473_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL mux_2947_nl : STD_LOGIC;
  SIGNAL mux_2946_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL mux_2945_nl : STD_LOGIC;
  SIGNAL nor_467_nl : STD_LOGIC;
  SIGNAL mux_2952_nl : STD_LOGIC;
  SIGNAL mux_2951_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL mux_2950_nl : STD_LOGIC;
  SIGNAL mux_2949_nl : STD_LOGIC;
  SIGNAL nor_461_nl : STD_LOGIC;
  SIGNAL mux_2948_nl : STD_LOGIC;
  SIGNAL mux_2955_nl : STD_LOGIC;
  SIGNAL mux_2954_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL mux_2953_nl : STD_LOGIC;
  SIGNAL nor_457_nl : STD_LOGIC;
  SIGNAL mux_2962_nl : STD_LOGIC;
  SIGNAL mux_2961_nl : STD_LOGIC;
  SIGNAL mux_2960_nl : STD_LOGIC;
  SIGNAL nor_449_nl : STD_LOGIC;
  SIGNAL nor_450_nl : STD_LOGIC;
  SIGNAL mux_2959_nl : STD_LOGIC;
  SIGNAL and_528_nl : STD_LOGIC;
  SIGNAL mux_2958_nl : STD_LOGIC;
  SIGNAL mux_2957_nl : STD_LOGIC;
  SIGNAL nor_452_nl : STD_LOGIC;
  SIGNAL mux_2956_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL mux_2965_nl : STD_LOGIC;
  SIGNAL mux_2964_nl : STD_LOGIC;
  SIGNAL nor_445_nl : STD_LOGIC;
  SIGNAL mux_2963_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL mux_2970_nl : STD_LOGIC;
  SIGNAL mux_2969_nl : STD_LOGIC;
  SIGNAL nor_439_nl : STD_LOGIC;
  SIGNAL mux_2968_nl : STD_LOGIC;
  SIGNAL mux_2967_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL mux_2966_nl : STD_LOGIC;
  SIGNAL mux_2973_nl : STD_LOGIC;
  SIGNAL mux_2972_nl : STD_LOGIC;
  SIGNAL nor_437_nl : STD_LOGIC;
  SIGNAL mux_2971_nl : STD_LOGIC;
  SIGNAL nor_438_nl : STD_LOGIC;
  SIGNAL mux_2979_nl : STD_LOGIC;
  SIGNAL mux_2978_nl : STD_LOGIC;
  SIGNAL mux_2977_nl : STD_LOGIC;
  SIGNAL and_789_nl : STD_LOGIC;
  SIGNAL and_810_nl : STD_LOGIC;
  SIGNAL mux_2976_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL nor_434_nl : STD_LOGIC;
  SIGNAL mux_2975_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL mux_2974_nl : STD_LOGIC;
  SIGNAL and_525_nl : STD_LOGIC;
  SIGNAL nor_436_nl : STD_LOGIC;
  SIGNAL mux_2982_nl : STD_LOGIC;
  SIGNAL mux_2981_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL mux_2980_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL mux_2987_nl : STD_LOGIC;
  SIGNAL mux_2986_nl : STD_LOGIC;
  SIGNAL and_790_nl : STD_LOGIC;
  SIGNAL mux_2985_nl : STD_LOGIC;
  SIGNAL mux_2984_nl : STD_LOGIC;
  SIGNAL and_520_nl : STD_LOGIC;
  SIGNAL mux_2983_nl : STD_LOGIC;
  SIGNAL mux_2990_nl : STD_LOGIC;
  SIGNAL mux_2989_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL mux_2988_nl : STD_LOGIC;
  SIGNAL and_517_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_721_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL and_1047_nl : STD_LOGIC;
  SIGNAL acc_1_nl : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_722_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nand_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux_723_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL STAGE_LOOP_mux_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_and_337_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux_64_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_146_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_or_88_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_and_312_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_147_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_or_89_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_or_90_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_mux_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux1h_148_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_1048_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_tmp_mux_65_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_tmp_or_91_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1267_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1268_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1890_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1891_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1892_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1893_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1894_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1895_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1896_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1269_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1897_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1898_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1899_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1900_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1901_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1902_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1903_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1270_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1271_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1904_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1905_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1906_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1907_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1908_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1909_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1910_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1272_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1273_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1274_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1275_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1911_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1912_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1913_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1914_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1915_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1916_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1917_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1276_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1277_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1278_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1279_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1280_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1281_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1282_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1283_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1918_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1919_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1920_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1921_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1922_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1923_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1924_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1284_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1285_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1286_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1287_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1288_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1289_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1290_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1291_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1292_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1293_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1294_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1295_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1296_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1297_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1298_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1299_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1925_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1926_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1927_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1928_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1929_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1930_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_1931_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1300_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1301_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1302_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1303_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1304_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1305_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1306_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1307_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1308_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1309_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1310_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1311_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1312_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1313_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1314_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1315_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1316_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1317_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1318_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1319_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1320_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1321_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1322_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1323_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1324_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1325_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1326_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1327_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1328_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1329_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_1330_nl : STD_LOGIC;
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT modulo_dev
    PORT (
      base_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1 : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat : STD_LOGIC;

  SIGNAL COMP_LOOP_5_tmp_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL COMP_LOOP_5_tmp_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_5_tmp_lshift_rg_z : STD_LOGIC_VECTOR (10 DOWNTO 0);

  SIGNAL COMP_LOOP_1_tmp_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_1_tmp_lshift_rg_z : STD_LOGIC_VECTOR (9 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_core_wait_dp
    PORT(
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT inPlaceNTT_DIF_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      COMP_LOOP_C_28_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_56_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_84_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_112_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_140_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_168_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_196_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_224_tr0 : IN STD_LOGIC;
      VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_1_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_5_2(input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_8_2(input_7 : STD_LOGIC;
  input_6 : STD_LOGIC;
  input_5 : STD_LOGIC;
  input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
      tmp := sel(5);
      result := result or ( input_5 and tmp);
      tmp := sel(6);
      result := result or ( input_6 and tmp);
      tmp := sel(7);
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_16_2(input_15 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_6_2(input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_7_2(input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_16_2(input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_32_2(input_31 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(31 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_3_2(input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_64_2(input_63 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_62 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_61 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_60 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_59 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_58 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_57 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_56 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_55 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_54 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_53 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_52 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_51 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_50 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_49 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_48 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_47 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_46 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_45 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_44 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_43 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_42 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_41 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_40 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_39 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_38 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_37 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_36 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_35 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_34 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_33 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_32 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(63 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
      tmp := (OTHERS=>sel( 32));
      result := result or ( input_32 and tmp);
      tmp := (OTHERS=>sel( 33));
      result := result or ( input_33 and tmp);
      tmp := (OTHERS=>sel( 34));
      result := result or ( input_34 and tmp);
      tmp := (OTHERS=>sel( 35));
      result := result or ( input_35 and tmp);
      tmp := (OTHERS=>sel( 36));
      result := result or ( input_36 and tmp);
      tmp := (OTHERS=>sel( 37));
      result := result or ( input_37 and tmp);
      tmp := (OTHERS=>sel( 38));
      result := result or ( input_38 and tmp);
      tmp := (OTHERS=>sel( 39));
      result := result or ( input_39 and tmp);
      tmp := (OTHERS=>sel( 40));
      result := result or ( input_40 and tmp);
      tmp := (OTHERS=>sel( 41));
      result := result or ( input_41 and tmp);
      tmp := (OTHERS=>sel( 42));
      result := result or ( input_42 and tmp);
      tmp := (OTHERS=>sel( 43));
      result := result or ( input_43 and tmp);
      tmp := (OTHERS=>sel( 44));
      result := result or ( input_44 and tmp);
      tmp := (OTHERS=>sel( 45));
      result := result or ( input_45 and tmp);
      tmp := (OTHERS=>sel( 46));
      result := result or ( input_46 and tmp);
      tmp := (OTHERS=>sel( 47));
      result := result or ( input_47 and tmp);
      tmp := (OTHERS=>sel( 48));
      result := result or ( input_48 and tmp);
      tmp := (OTHERS=>sel( 49));
      result := result or ( input_49 and tmp);
      tmp := (OTHERS=>sel( 50));
      result := result or ( input_50 and tmp);
      tmp := (OTHERS=>sel( 51));
      result := result or ( input_51 and tmp);
      tmp := (OTHERS=>sel( 52));
      result := result or ( input_52 and tmp);
      tmp := (OTHERS=>sel( 53));
      result := result or ( input_53 and tmp);
      tmp := (OTHERS=>sel( 54));
      result := result or ( input_54 and tmp);
      tmp := (OTHERS=>sel( 55));
      result := result or ( input_55 and tmp);
      tmp := (OTHERS=>sel( 56));
      result := result or ( input_56 and tmp);
      tmp := (OTHERS=>sel( 57));
      result := result or ( input_57 and tmp);
      tmp := (OTHERS=>sel( 58));
      result := result or ( input_58 and tmp);
      tmp := (OTHERS=>sel( 59));
      result := result or ( input_59 and tmp);
      tmp := (OTHERS=>sel( 60));
      result := result or ( input_60 and tmp);
      tmp := (OTHERS=>sel( 61));
      result := result or ( input_61 and tmp);
      tmp := (OTHERS=>sel( 62));
      result := result or ( input_62 and tmp);
      tmp := (OTHERS=>sel( 63));
      result := result or ( input_63 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_65_2(input_64 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_63 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_62 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_61 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_60 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_59 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_58 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_57 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_56 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_55 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_54 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_53 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_52 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_51 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_50 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_49 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_48 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_47 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_46 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_45 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_44 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_43 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_42 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_41 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_40 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_39 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_38 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_37 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_36 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_35 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_34 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_33 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_32 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(64 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
      tmp := (OTHERS=>sel( 32));
      result := result or ( input_32 and tmp);
      tmp := (OTHERS=>sel( 33));
      result := result or ( input_33 and tmp);
      tmp := (OTHERS=>sel( 34));
      result := result or ( input_34 and tmp);
      tmp := (OTHERS=>sel( 35));
      result := result or ( input_35 and tmp);
      tmp := (OTHERS=>sel( 36));
      result := result or ( input_36 and tmp);
      tmp := (OTHERS=>sel( 37));
      result := result or ( input_37 and tmp);
      tmp := (OTHERS=>sel( 38));
      result := result or ( input_38 and tmp);
      tmp := (OTHERS=>sel( 39));
      result := result or ( input_39 and tmp);
      tmp := (OTHERS=>sel( 40));
      result := result or ( input_40 and tmp);
      tmp := (OTHERS=>sel( 41));
      result := result or ( input_41 and tmp);
      tmp := (OTHERS=>sel( 42));
      result := result or ( input_42 and tmp);
      tmp := (OTHERS=>sel( 43));
      result := result or ( input_43 and tmp);
      tmp := (OTHERS=>sel( 44));
      result := result or ( input_44 and tmp);
      tmp := (OTHERS=>sel( 45));
      result := result or ( input_45 and tmp);
      tmp := (OTHERS=>sel( 46));
      result := result or ( input_46 and tmp);
      tmp := (OTHERS=>sel( 47));
      result := result or ( input_47 and tmp);
      tmp := (OTHERS=>sel( 48));
      result := result or ( input_48 and tmp);
      tmp := (OTHERS=>sel( 49));
      result := result or ( input_49 and tmp);
      tmp := (OTHERS=>sel( 50));
      result := result or ( input_50 and tmp);
      tmp := (OTHERS=>sel( 51));
      result := result or ( input_51 and tmp);
      tmp := (OTHERS=>sel( 52));
      result := result or ( input_52 and tmp);
      tmp := (OTHERS=>sel( 53));
      result := result or ( input_53 and tmp);
      tmp := (OTHERS=>sel( 54));
      result := result or ( input_54 and tmp);
      tmp := (OTHERS=>sel( 55));
      result := result or ( input_55 and tmp);
      tmp := (OTHERS=>sel( 56));
      result := result or ( input_56 and tmp);
      tmp := (OTHERS=>sel( 57));
      result := result or ( input_57 and tmp);
      tmp := (OTHERS=>sel( 58));
      result := result or ( input_58 and tmp);
      tmp := (OTHERS=>sel( 59));
      result := result or ( input_59 and tmp);
      tmp := (OTHERS=>sel( 60));
      result := result or ( input_60 and tmp);
      tmp := (OTHERS=>sel( 61));
      result := result or ( input_61 and tmp);
      tmp := (OTHERS=>sel( 62));
      result := result or ( input_62 and tmp);
      tmp := (OTHERS=>sel( 63));
      result := result or ( input_63 and tmp);
      tmp := (OTHERS=>sel( 64));
      result := result or ( input_64 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_68_2(input_67 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_66 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_65 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_64 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_63 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_62 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_61 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_60 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_59 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_58 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_57 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_56 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_55 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_54 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_53 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_52 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_51 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_50 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_49 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_48 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_47 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_46 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_45 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_44 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_43 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_42 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_41 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_40 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_39 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_38 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_37 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_36 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_35 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_34 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_33 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_32 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(67 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
      tmp := (OTHERS=>sel( 32));
      result := result or ( input_32 and tmp);
      tmp := (OTHERS=>sel( 33));
      result := result or ( input_33 and tmp);
      tmp := (OTHERS=>sel( 34));
      result := result or ( input_34 and tmp);
      tmp := (OTHERS=>sel( 35));
      result := result or ( input_35 and tmp);
      tmp := (OTHERS=>sel( 36));
      result := result or ( input_36 and tmp);
      tmp := (OTHERS=>sel( 37));
      result := result or ( input_37 and tmp);
      tmp := (OTHERS=>sel( 38));
      result := result or ( input_38 and tmp);
      tmp := (OTHERS=>sel( 39));
      result := result or ( input_39 and tmp);
      tmp := (OTHERS=>sel( 40));
      result := result or ( input_40 and tmp);
      tmp := (OTHERS=>sel( 41));
      result := result or ( input_41 and tmp);
      tmp := (OTHERS=>sel( 42));
      result := result or ( input_42 and tmp);
      tmp := (OTHERS=>sel( 43));
      result := result or ( input_43 and tmp);
      tmp := (OTHERS=>sel( 44));
      result := result or ( input_44 and tmp);
      tmp := (OTHERS=>sel( 45));
      result := result or ( input_45 and tmp);
      tmp := (OTHERS=>sel( 46));
      result := result or ( input_46 and tmp);
      tmp := (OTHERS=>sel( 47));
      result := result or ( input_47 and tmp);
      tmp := (OTHERS=>sel( 48));
      result := result or ( input_48 and tmp);
      tmp := (OTHERS=>sel( 49));
      result := result or ( input_49 and tmp);
      tmp := (OTHERS=>sel( 50));
      result := result or ( input_50 and tmp);
      tmp := (OTHERS=>sel( 51));
      result := result or ( input_51 and tmp);
      tmp := (OTHERS=>sel( 52));
      result := result or ( input_52 and tmp);
      tmp := (OTHERS=>sel( 53));
      result := result or ( input_53 and tmp);
      tmp := (OTHERS=>sel( 54));
      result := result or ( input_54 and tmp);
      tmp := (OTHERS=>sel( 55));
      result := result or ( input_55 and tmp);
      tmp := (OTHERS=>sel( 56));
      result := result or ( input_56 and tmp);
      tmp := (OTHERS=>sel( 57));
      result := result or ( input_57 and tmp);
      tmp := (OTHERS=>sel( 58));
      result := result or ( input_58 and tmp);
      tmp := (OTHERS=>sel( 59));
      result := result or ( input_59 and tmp);
      tmp := (OTHERS=>sel( 60));
      result := result or ( input_60 and tmp);
      tmp := (OTHERS=>sel( 61));
      result := result or ( input_61 and tmp);
      tmp := (OTHERS=>sel( 62));
      result := result or ( input_62 and tmp);
      tmp := (OTHERS=>sel( 63));
      result := result or ( input_63 and tmp);
      tmp := (OTHERS=>sel( 64));
      result := result or ( input_64 and tmp);
      tmp := (OTHERS=>sel( 65));
      result := result or ( input_65 and tmp);
      tmp := (OTHERS=>sel( 66));
      result := result or ( input_66 and tmp);
      tmp := (OTHERS=>sel( 67));
      result := result or ( input_67 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_8_2(input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_9_2(input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_3_2(input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_9_4_2(input_3 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_11_2_2(input_0 : STD_LOGIC_VECTOR(10 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(10 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(10 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_9_2_2(input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION minimum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1<arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION maximum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1>arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION READSLICE_64_65(input_val:STD_LOGIC_VECTOR(64 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC_VECTOR IS
    CONSTANT min_sat_index:INTEGER:= maximum( index, 0 );
    CONSTANT sat_index:INTEGER:= minimum( min_sat_index, 1);
  BEGIN
    RETURN input_val(sat_index+63 DOWNTO sat_index);
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 5,
      width => 64
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  vec_rsc_triosy_0_63_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_63_lz
    );
  vec_rsc_triosy_0_62_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_62_lz
    );
  vec_rsc_triosy_0_61_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_61_lz
    );
  vec_rsc_triosy_0_60_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_60_lz
    );
  vec_rsc_triosy_0_59_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_59_lz
    );
  vec_rsc_triosy_0_58_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_58_lz
    );
  vec_rsc_triosy_0_57_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_57_lz
    );
  vec_rsc_triosy_0_56_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_56_lz
    );
  vec_rsc_triosy_0_55_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_55_lz
    );
  vec_rsc_triosy_0_54_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_54_lz
    );
  vec_rsc_triosy_0_53_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_53_lz
    );
  vec_rsc_triosy_0_52_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_52_lz
    );
  vec_rsc_triosy_0_51_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_51_lz
    );
  vec_rsc_triosy_0_50_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_50_lz
    );
  vec_rsc_triosy_0_49_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_49_lz
    );
  vec_rsc_triosy_0_48_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_48_lz
    );
  vec_rsc_triosy_0_47_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_47_lz
    );
  vec_rsc_triosy_0_46_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_46_lz
    );
  vec_rsc_triosy_0_45_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_45_lz
    );
  vec_rsc_triosy_0_44_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_44_lz
    );
  vec_rsc_triosy_0_43_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_43_lz
    );
  vec_rsc_triosy_0_42_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_42_lz
    );
  vec_rsc_triosy_0_41_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_41_lz
    );
  vec_rsc_triosy_0_40_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_40_lz
    );
  vec_rsc_triosy_0_39_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_39_lz
    );
  vec_rsc_triosy_0_38_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_38_lz
    );
  vec_rsc_triosy_0_37_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_37_lz
    );
  vec_rsc_triosy_0_36_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_36_lz
    );
  vec_rsc_triosy_0_35_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_35_lz
    );
  vec_rsc_triosy_0_34_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_34_lz
    );
  vec_rsc_triosy_0_33_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_33_lz
    );
  vec_rsc_triosy_0_32_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_32_lz
    );
  vec_rsc_triosy_0_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_31_lz
    );
  vec_rsc_triosy_0_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_30_lz
    );
  vec_rsc_triosy_0_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_29_lz
    );
  vec_rsc_triosy_0_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_28_lz
    );
  vec_rsc_triosy_0_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_27_lz
    );
  vec_rsc_triosy_0_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_26_lz
    );
  vec_rsc_triosy_0_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_25_lz
    );
  vec_rsc_triosy_0_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_24_lz
    );
  vec_rsc_triosy_0_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_23_lz
    );
  vec_rsc_triosy_0_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_22_lz
    );
  vec_rsc_triosy_0_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_21_lz
    );
  vec_rsc_triosy_0_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_20_lz
    );
  vec_rsc_triosy_0_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_19_lz
    );
  vec_rsc_triosy_0_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_18_lz
    );
  vec_rsc_triosy_0_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_17_lz
    );
  vec_rsc_triosy_0_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_16_lz
    );
  vec_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_15_lz
    );
  vec_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_14_lz
    );
  vec_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_13_lz
    );
  vec_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_12_lz
    );
  vec_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_11_lz
    );
  vec_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_10_lz
    );
  vec_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_9_lz
    );
  vec_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_8_lz
    );
  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_7_lz
    );
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_6_lz
    );
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_5_lz
    );
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_4_lz
    );
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_3_lz
    );
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_2_lz
    );
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_1_lz
    );
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => vec_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  twiddle_rsc_triosy_0_63_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_63_lz
    );
  twiddle_rsc_triosy_0_62_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_62_lz
    );
  twiddle_rsc_triosy_0_61_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_61_lz
    );
  twiddle_rsc_triosy_0_60_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_60_lz
    );
  twiddle_rsc_triosy_0_59_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_59_lz
    );
  twiddle_rsc_triosy_0_58_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_58_lz
    );
  twiddle_rsc_triosy_0_57_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_57_lz
    );
  twiddle_rsc_triosy_0_56_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_56_lz
    );
  twiddle_rsc_triosy_0_55_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_55_lz
    );
  twiddle_rsc_triosy_0_54_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_54_lz
    );
  twiddle_rsc_triosy_0_53_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_53_lz
    );
  twiddle_rsc_triosy_0_52_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_52_lz
    );
  twiddle_rsc_triosy_0_51_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_51_lz
    );
  twiddle_rsc_triosy_0_50_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_50_lz
    );
  twiddle_rsc_triosy_0_49_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_49_lz
    );
  twiddle_rsc_triosy_0_48_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_48_lz
    );
  twiddle_rsc_triosy_0_47_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_47_lz
    );
  twiddle_rsc_triosy_0_46_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_46_lz
    );
  twiddle_rsc_triosy_0_45_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_45_lz
    );
  twiddle_rsc_triosy_0_44_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_44_lz
    );
  twiddle_rsc_triosy_0_43_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_43_lz
    );
  twiddle_rsc_triosy_0_42_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_42_lz
    );
  twiddle_rsc_triosy_0_41_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_41_lz
    );
  twiddle_rsc_triosy_0_40_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_40_lz
    );
  twiddle_rsc_triosy_0_39_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_39_lz
    );
  twiddle_rsc_triosy_0_38_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_38_lz
    );
  twiddle_rsc_triosy_0_37_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_37_lz
    );
  twiddle_rsc_triosy_0_36_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_36_lz
    );
  twiddle_rsc_triosy_0_35_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_35_lz
    );
  twiddle_rsc_triosy_0_34_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_34_lz
    );
  twiddle_rsc_triosy_0_33_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_33_lz
    );
  twiddle_rsc_triosy_0_32_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_32_lz
    );
  twiddle_rsc_triosy_0_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_31_lz
    );
  twiddle_rsc_triosy_0_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_30_lz
    );
  twiddle_rsc_triosy_0_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_29_lz
    );
  twiddle_rsc_triosy_0_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_28_lz
    );
  twiddle_rsc_triosy_0_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_27_lz
    );
  twiddle_rsc_triosy_0_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_26_lz
    );
  twiddle_rsc_triosy_0_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_25_lz
    );
  twiddle_rsc_triosy_0_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_24_lz
    );
  twiddle_rsc_triosy_0_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_23_lz
    );
  twiddle_rsc_triosy_0_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_22_lz
    );
  twiddle_rsc_triosy_0_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_21_lz
    );
  twiddle_rsc_triosy_0_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_20_lz
    );
  twiddle_rsc_triosy_0_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_19_lz
    );
  twiddle_rsc_triosy_0_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_18_lz
    );
  twiddle_rsc_triosy_0_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_17_lz
    );
  twiddle_rsc_triosy_0_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_16_lz
    );
  twiddle_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_15_lz
    );
  twiddle_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_14_lz
    );
  twiddle_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_13_lz
    );
  twiddle_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_12_lz
    );
  twiddle_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_11_lz
    );
  twiddle_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_10_lz
    );
  twiddle_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_9_lz
    );
  twiddle_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_8_lz
    );
  twiddle_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_7_lz
    );
  twiddle_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_6_lz
    );
  twiddle_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_5_lz
    );
  twiddle_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_4_lz
    );
  twiddle_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_3_lz
    );
  twiddle_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_2_lz
    );
  twiddle_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_1_lz
    );
  twiddle_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_63_obj_ld_cse,
      lz => twiddle_rsc_triosy_0_0_lz
    );
  COMP_LOOP_1_modulo_dev_cmp : modulo_dev
    PORT MAP(
      base_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat,
      m_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat,
      return_rsc_z => COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1,
      ccs_ccore_start_rsc_dat => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => clk,
      ccs_ccore_srst => rst,
      ccs_ccore_en => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
    );
  COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat <= MUX1HOT_v_64_3_2((READSLICE_64_65(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_724_cse
      & '1') + UNSIGNED((MUX_v_64_2_2((NOT COMP_LOOP_1_acc_8_itm), (NOT z_out_9),
      COMP_LOOP_or_65_itm)) & '1'), 65)), 1)), COMP_LOOP_1_acc_8_itm, z_out_8, STD_LOGIC_VECTOR'(
      COMP_LOOP_or_68_itm & ((NOT (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_3721,
      mux_tmp_2924, fsm_output(6))), or_tmp_3718, fsm_output(2))), (MUX_s_1_2_2(or_tmp_3718,
      (MUX_s_1_2_2(mux_tmp_2924, ((NOT (fsm_output(4))) OR (fsm_output(3)) OR (fsm_output(7))),
      fsm_output(6))), fsm_output(2))), fsm_output(5)))) AND and_dcpl_340) & ((and_dcpl_92
      AND and_dcpl_57) OR (and_dcpl_262 AND and_dcpl_344) OR (and_dcpl_262 AND and_dcpl_347)
      OR (and_dcpl_60 AND and_dcpl_64) OR (and_dcpl_66 AND and_dcpl_57) OR (and_dcpl_355
      AND and_dcpl_110) OR (and_dcpl_355 AND and_dcpl_113) OR (and_dcpl_353 AND and_dcpl_116))));
  COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat <= p_sva;
  COMP_LOOP_1_modulo_dev_cmp_return_rsc_z <= COMP_LOOP_1_modulo_dev_cmp_return_rsc_z_1;
  COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat <= NOT((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(((fsm_output(3))
      OR (NOT (MUX_s_1_2_2(or_364_cse, and_735_cse, fsm_output(0))))), nand_tmp_142,
      fsm_output(6))), ((fsm_output(6)) OR mux_tmp_2939), fsm_output(5))), (MUX_s_1_2_2((MUX_s_1_2_2(mux_tmp_2939,
      ((fsm_output(3)) OR (fsm_output(0)) OR (NOT and_735_cse)), fsm_output(6))),
      (MUX_s_1_2_2(nand_tmp_142, ((fsm_output(3)) OR (NOT((NOT (fsm_output(0))) OR
      (fsm_output(4)))) OR (fsm_output(7))), fsm_output(6))), fsm_output(5))), fsm_output(2)))
      OR (fsm_output(1)));

  COMP_LOOP_5_tmp_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 11
      )
    PORT MAP(
      a => COMP_LOOP_5_tmp_lshift_rg_a,
      s => COMP_LOOP_5_tmp_lshift_rg_s,
      z => COMP_LOOP_5_tmp_lshift_rg_z
    );
  COMP_LOOP_5_tmp_lshift_rg_a(0) <= '1';
  COMP_LOOP_5_tmp_lshift_rg_s <= MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, z_out_4, CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("00000010")));
  z_out <= COMP_LOOP_5_tmp_lshift_rg_z;

  COMP_LOOP_1_tmp_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 10
      )
    PORT MAP(
      a => COMP_LOOP_1_tmp_lshift_rg_a,
      s => COMP_LOOP_1_tmp_lshift_rg_s,
      z => COMP_LOOP_1_tmp_lshift_rg_z
    );
  COMP_LOOP_1_tmp_lshift_rg_a(0) <= '1';
  COMP_LOOP_1_tmp_lshift_rg_s <= MUX_v_4_2_2(z_out_4, COMP_LOOP_1_tmp_acc_cse_sva,
      ((NOT (fsm_output(4))) AND (fsm_output(0)) AND nor_1715_cse AND CONV_SL_1_1(fsm_output(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("01")) AND nor_1716_cse) OR ((NOT (fsm_output(4)))
      AND (NOT (fsm_output(0))) AND nor_1715_cse AND CONV_SL_1_1(fsm_output(2 DOWNTO
      1)=STD_LOGIC_VECTOR'("10")) AND nor_1716_cse));
  z_out_1 <= COMP_LOOP_1_tmp_lshift_rg_z;

  inPlaceNTT_DIF_core_wait_dp_inst : inPlaceNTT_DIF_core_wait_dp
    PORT MAP(
      ensig_cgo_iro => mux_2997_rmff,
      ensig_cgo => reg_ensig_cgo_cse,
      COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en => COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
    );
  inPlaceNTT_DIF_core_core_fsm_inst : inPlaceNTT_DIF_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => inPlaceNTT_DIF_core_core_fsm_inst_fsm_output,
      COMP_LOOP_C_28_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0,
      COMP_LOOP_C_56_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0,
      COMP_LOOP_C_84_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0,
      COMP_LOOP_C_112_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0,
      COMP_LOOP_C_140_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0,
      COMP_LOOP_C_168_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0,
      COMP_LOOP_C_196_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0,
      COMP_LOOP_C_224_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0,
      VEC_LOOP_C_0_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_1_tr0 => inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0
    );
  fsm_output <= inPlaceNTT_DIF_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0 <= NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0 <= NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0 <= NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0 <= NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0 <= NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0 <= NOT COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 <= z_out_3(10);
  inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 <= NOT (z_out_2(4));

  or_595_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  nand_191_cse <= NOT((z_out_7(0)) AND (fsm_output(3)));
  nand_190_cse <= NOT(CONV_SL_1_1(z_out_7(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      (fsm_output(3)));
  nand_188_cse <= NOT(CONV_SL_1_1(z_out_7(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND
      (fsm_output(3)));
  nand_184_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(3)));
  nand_174_cse <= NOT((COMP_LOOP_3_tmp_lshift_ncse_sva(4)) AND (fsm_output(3)));
  nand_175_cse <= NOT((COMP_LOOP_2_tmp_lshift_ncse_sva(5)) AND (fsm_output(3)));
  mux_2995_nl <= MUX_s_1_2_2(mux_tmp_2924, mux_tmp_2927, fsm_output(6));
  mux_2996_nl <= MUX_s_1_2_2(or_tmp_3718, mux_2995_nl, fsm_output(2));
  nor_425_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10"))))
      OR (fsm_output(7)));
  mux_2992_nl <= MUX_s_1_2_2(mux_tmp_2924, nor_425_nl, fsm_output(6));
  mux_2993_nl <= MUX_s_1_2_2(mux_2992_nl, (NOT and_705_cse), fsm_output(2));
  mux_2997_rmff <= MUX_s_1_2_2(mux_2996_nl, mux_2993_nl, fsm_output(5));
  or_4007_cse <= (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(3));
  and_78_cse <= (fsm_output(6)) AND or_4007_cse AND (fsm_output(7));
  nor_1744_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_1046_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  mux_3029_nl <= MUX_s_1_2_2(mux_tmp_2959, mux_tmp_2961, fsm_output(2));
  mux_3030_nl <= MUX_s_1_2_2(mux_3029_nl, mux_tmp_2960, fsm_output(1));
  mux_3031_nl <= MUX_s_1_2_2(mux_3030_nl, (fsm_output(6)), fsm_output(5));
  COMP_LOOP_or_121_cse <= mux_3031_nl OR (fsm_output(7));
  and_507_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  nor_1674_cse <= NOT((fsm_output(2)) OR (fsm_output(6)));
  COMP_LOOP_or_120_rgt <= and_dcpl_259 OR and_dcpl_260 OR and_dcpl_263;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001010"));
  COMP_LOOP_tmp_nor_67_cse <= NOT((z_out_7(4)) OR (z_out_7(2)) OR (z_out_7(1)));
  mux_3044_nl <= MUX_s_1_2_2(mux_tmp_2976, mux_tmp_2975, fsm_output(1));
  mux_3045_nl <= MUX_s_1_2_2(mux_3044_nl, (NOT mux_180_cse), fsm_output(5));
  COMP_LOOP_or_126_cse <= NOT(mux_3045_nl AND (NOT (fsm_output(7))));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_78_cse <= (z_out_7(3)) AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_67_cse;
  nor_358_cse <= NOT((fsm_output(5)) OR (NOT (fsm_output(0))));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001100"));
  COMP_LOOP_tmp_nor_68_cse <= NOT((z_out_7(4)) OR (z_out_7(2)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_79_cse <= (z_out_7(3)) AND (z_out_7(1)) AND COMP_LOOP_tmp_nor_68_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001101"));
  COMP_LOOP_tmp_nor_69_cse <= NOT((z_out_7(4)) OR (z_out_7(2)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_cse <= (z_out_7(3)) AND (z_out_7(1)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_69_cse;
  or_341_cse <= (fsm_output(4)) OR (fsm_output(6));
  and_677_cse <= (fsm_output(3)) AND (fsm_output(4)) AND (fsm_output(6));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001110"));
  COMP_LOOP_tmp_nor_70_cse <= NOT((z_out_7(4)) OR (z_out_7(1)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_nor_70_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001111"));
  COMP_LOOP_tmp_nor_71_cse <= NOT((z_out_7(4)) OR (z_out_7(1)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_cse <= (z_out_7(3)) AND (z_out_7(2)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_71_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_23_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010001"));
  COMP_LOOP_tmp_nor_72_cse <= NOT((z_out_7(4)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_cse <= CONV_SL_1_1(z_out_7(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_tmp_nor_72_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_27_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
  COMP_LOOP_tmp_nor_76_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010100"));
  COMP_LOOP_or_135_cse <= MUX_s_1_2_2(mux_tmp_3003, (fsm_output(7)), fsm_output(5));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_88_cse <= (z_out_7(4)) AND (z_out_7(1)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_76_cse;
  and_640_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"));
  and_639_cse <= (fsm_output(3)) AND (fsm_output(0));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_28_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010110"));
  COMP_LOOP_tmp_nor_77_cse <= NOT((z_out_7(3)) OR (z_out_7(1)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_89_cse <= (z_out_7(4)) AND (z_out_7(2)) AND COMP_LOOP_tmp_nor_77_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_29_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010111"));
  COMP_LOOP_tmp_nor_78_cse <= NOT((z_out_7(3)) OR (z_out_7(1)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_90_cse <= (z_out_7(4)) AND (z_out_7(2)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_78_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_30_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011000"));
  COMP_LOOP_tmp_nor_79_cse <= NOT((z_out_7(3)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_91_cse <= (z_out_7(4)) AND (z_out_7(2)) AND (z_out_7(1))
      AND COMP_LOOP_tmp_nor_79_cse;
  or_359_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  and_673_cse <= (fsm_output(6)) AND (fsm_output(4));
  or_364_cse <= (fsm_output(4)) OR (fsm_output(7));
  COMP_LOOP_or_110_rgt <= and_dcpl_77 OR and_dcpl_259;
  COMP_LOOP_tmp_nor_208_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_244_cse <= CONV_SL_1_1(z_out_7(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_nor_208_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_31_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011001"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_92_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"));
  nor_412_cse <= NOT((NOT (fsm_output(5))) OR (fsm_output(7)));
  or_3900_nl <= and_507_cse OR (fsm_output(7));
  mux_3094_nl <= MUX_s_1_2_2(or_3900_nl, or_tmp_3773, fsm_output(3));
  mux_3095_cse <= MUX_s_1_2_2((fsm_output(7)), mux_3094_nl, fsm_output(0));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_32_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011010"));
  COMP_LOOP_tmp_nor_80_cse <= NOT(CONV_SL_1_1(z_out_7(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_93_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_nor_80_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_33_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011011"));
  COMP_LOOP_tmp_nor_81_cse <= NOT(CONV_SL_1_1(z_out_7(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_94_cse <= (z_out_7(4)) AND (z_out_7(3)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_81_cse;
  or_560_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_742_cse <= MUX_s_1_2_2(or_560_nl, (fsm_output(7)), fsm_output(6));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011100"));
  COMP_LOOP_tmp_nor_82_cse <= NOT((z_out_7(2)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_95_cse <= (z_out_7(4)) AND (z_out_7(3)) AND (z_out_7(1))
      AND COMP_LOOP_tmp_nor_82_cse;
  or_564_cse <= (NOT (fsm_output(5))) OR (fsm_output(7));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_96_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"));
  COMP_LOOP_tmp_nor_83_cse <= NOT(CONV_SL_1_1(z_out_7(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_97_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_tmp_nor_83_cse;
  mux_297_cse <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(6));
  and_808_cse <= (fsm_output(2)) AND (fsm_output(6));
  and_763_cse <= (fsm_output(3)) AND (fsm_output(7));
  or_154_nl <= (fsm_output(2)) OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(3));
  mux_221_cse <= MUX_s_1_2_2(or_80_cse, or_154_nl, fsm_output(1));
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
  COMP_LOOP_tmp_nor_140_cse <= NOT(CONV_SL_1_1(z_out_7(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_tmp_nor_141_cse <= NOT((z_out_7(3)) OR (z_out_7(2)) OR (z_out_7(0)));
  and_493_cse <= (fsm_output(5)) AND (fsm_output(7));
  or_4057_cse <= (fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(3));
  and_736_cse <= or_4057_cse AND (fsm_output(7));
  and_705_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  mux_180_cse <= MUX_s_1_2_2(and_677_cse, and_673_cse, fsm_output(2));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_24_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010010"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_25_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_cse <= (z_out_7(4)) AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_140_cse;
  nor_1683_cse <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_87_cse <= (z_out_7(4)) AND (z_out_7(1)) AND COMP_LOOP_tmp_nor_141_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_98_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"));
  mux_3233_nl <= MUX_s_1_2_2(mux_tmp_3100, mux_tmp_3098, fsm_output(2));
  mux_3234_nl <= MUX_s_1_2_2(mux_3233_nl, mux_tmp_3101, fsm_output(1));
  COMP_LOOP_or_151_cse <= MUX_s_1_2_2(mux_3234_nl, mux_tmp_3119, fsm_output(5));
  mux_3237_nl <= MUX_s_1_2_2(mux_tmp_3169, (fsm_output(7)), fsm_output(6));
  mux_3238_nl <= MUX_s_1_2_2(mux_tmp_656, mux_3237_nl, fsm_output(2));
  COMP_LOOP_or_153_cse <= MUX_s_1_2_2(mux_tmp_3102, mux_3238_nl, fsm_output(5));
  COMP_LOOP_tmp_nor_34_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse <= (z_out_7(5)) AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_34_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_99_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"));
  nor_399_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  or_477_cse <= (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(7));
  and_655_cse <= or_595_cse AND (fsm_output(7));
  nor_398_cse <= NOT((fsm_output(4)) OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  COMP_LOOP_tmp_nor_35_cse <= NOT((z_out_7(4)) OR (z_out_7(3)) OR (z_out_7(2)) OR
      (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse <= (z_out_7(5)) AND (z_out_7(1)) AND COMP_LOOP_tmp_nor_35_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
  COMP_LOOP_tmp_or_cse <= and_dcpl_74 OR and_dcpl_77 OR and_dcpl_258 OR and_dcpl_259
      OR and_dcpl_260 OR and_dcpl_263;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("000101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("000011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("000110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("000111"));
  COMP_LOOP_tmp_nor_63_cse <= NOT((z_out_7(4)) OR (z_out_7(3)) OR (z_out_7(1)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_74_cse <= (z_out_7(2)) AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_63_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001001"));
  COMP_LOOP_tmp_nor_64_cse <= NOT((z_out_7(4)) OR (z_out_7(3)) OR (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_75_cse <= CONV_SL_1_1(z_out_7(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_nor_64_cse;
  COMP_LOOP_tmp_nor_65_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_76_cse <= CONV_SL_1_1(z_out_7(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_tmp_nor_65_cse;
  COMP_LOOP_tmp_or_5_cse <= and_dcpl_74 OR and_dcpl_77 OR and_dcpl_259 OR and_dcpl_260
      OR and_dcpl_263;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_cse <= (z_out_7(5)) AND (z_out_7(1)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_208_cse;
  COMP_LOOP_tmp_nor_37_cse <= NOT((z_out_7(4)) OR (z_out_7(3)) OR (z_out_7(1)) OR
      (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse <= (z_out_7(5)) AND (z_out_7(2)) AND COMP_LOOP_tmp_nor_37_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse <= (z_out_7(5)) AND (z_out_7(2)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_63_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse <= (z_out_7(5)) AND (z_out_7(2)) AND (z_out_7(1))
      AND COMP_LOOP_tmp_nor_64_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse <= (z_out_7(5)) AND (z_out_7(2)) AND (z_out_7(1))
      AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_65_cse;
  COMP_LOOP_tmp_nor_41_cse <= NOT((z_out_7(4)) OR (z_out_7(2)) OR (z_out_7(1)) OR
      (z_out_7(0)));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse <= (z_out_7(5)) AND (z_out_7(3)) AND COMP_LOOP_tmp_nor_41_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse <= (z_out_7(5)) AND (z_out_7(3)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_67_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse <= (z_out_7(5)) AND (z_out_7(3)) AND (z_out_7(1))
      AND COMP_LOOP_tmp_nor_68_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_49_cse <= (z_out_7(5)) AND (z_out_7(3)) AND (z_out_7(1))
      AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_69_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_50_cse <= (z_out_7(5)) AND (z_out_7(3)) AND (z_out_7(2))
      AND COMP_LOOP_tmp_nor_70_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse <= (z_out_7(5)) AND (z_out_7(3)) AND (z_out_7(2))
      AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_71_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_52_cse <= (z_out_7(5)) AND (z_out_7(3)) AND (z_out_7(2))
      AND (z_out_7(1)) AND COMP_LOOP_tmp_nor_72_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse <= (z_out_7(5)) AND (z_out_7(4)) AND (z_out_7(0))
      AND COMP_LOOP_tmp_nor_140_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_56_cse <= (z_out_7(5)) AND (z_out_7(4)) AND (z_out_7(1))
      AND COMP_LOOP_tmp_nor_141_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_57_cse <= (z_out_7(5)) AND (z_out_7(4)) AND (z_out_7(1))
      AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_76_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_58_cse <= (z_out_7(5)) AND (z_out_7(4)) AND (z_out_7(2))
      AND COMP_LOOP_tmp_nor_77_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_59_cse <= (z_out_7(5)) AND (z_out_7(4)) AND (z_out_7(2))
      AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_78_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_60_cse <= (z_out_7(5)) AND (z_out_7(4)) AND (z_out_7(2))
      AND (z_out_7(1)) AND COMP_LOOP_tmp_nor_79_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_61_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_62_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 3)=STD_LOGIC_VECTOR'("111"))
      AND COMP_LOOP_tmp_nor_80_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_63_cse <= (z_out_7(5)) AND (z_out_7(4)) AND (z_out_7(3))
      AND (z_out_7(0)) AND COMP_LOOP_tmp_nor_81_cse;
  COMP_LOOP_tmp_nor_150_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
  COMP_LOOP_or_74_cse <= and_dcpl_260 OR and_dcpl_263;
  COMP_LOOP_tmp_nor_10_cse <= NOT((z_out_7(5)) OR (z_out_7(4)) OR (z_out_7(2)) OR
      (z_out_7(1)) OR (z_out_7(0)));
  COMP_LOOP_tmp_nor_151_cse <= NOT((z_out_7(5)) OR (z_out_7(4)) OR (z_out_7(3)) OR
      (z_out_7(2)) OR (z_out_7(0)));
  COMP_LOOP_tmp_nor_18_cse <= NOT((z_out_7(5)) OR (z_out_7(3)) OR (z_out_7(2)) OR
      (z_out_7(1)) OR (z_out_7(0)));
  COMP_LOOP_tmp_nor_153_cse <= NOT((z_out_7(5)) OR (z_out_7(4)) OR (z_out_7(3)) OR
      (z_out_7(1)) OR (z_out_7(0)));
  COMP_LOOP_or_68_itm <= and_dcpl_258 OR and_dcpl_343 OR and_dcpl_346 OR and_dcpl_349
      OR and_dcpl_351 OR and_dcpl_354 OR and_dcpl_357 OR and_dcpl_359;
  COMP_LOOP_tmp_or_36_cse <= and_dcpl_77 OR and_dcpl_259 OR and_dcpl_260 OR and_dcpl_263;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_64_cse <= (z_out_7(5)) AND (z_out_7(4)) AND (z_out_7(3))
      AND (z_out_7(1)) AND COMP_LOOP_tmp_nor_82_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_65_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_66_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 2)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_tmp_nor_83_cse;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_67_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_68_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_69_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
  COMP_LOOP_tmp_or_43_cse <= and_dcpl_258 OR and_dcpl_261;
  or_80_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"));
  and_478_m1c <= and_dcpl_262 AND and_dcpl_73;
  mux_3357_nl <= MUX_s_1_2_2(not_tmp_868, (fsm_output(7)), fsm_output(6));
  mux_3358_nl <= MUX_s_1_2_2(mux_3357_nl, mux_tmp_3288, fsm_output(2));
  mux_3356_nl <= MUX_s_1_2_2(mux_tmp_3100, mux_tmp_3288, fsm_output(2));
  mux_3359_nl <= MUX_s_1_2_2(mux_3358_nl, mux_3356_nl, fsm_output(1));
  mux_3360_tmp <= MUX_s_1_2_2(mux_3359_nl, (fsm_output(7)), fsm_output(5));
  and_735_cse <= (fsm_output(4)) AND (fsm_output(7));
  COMP_LOOP_1_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "000")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_1_acc_10_itm_10_1_1 <= COMP_LOOP_1_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_acc_psp_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
      DOWNTO 3)) + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0), 7));
  COMP_LOOP_acc_14_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
      DOWNTO 1)) + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "11")),
      9));
  COMP_LOOP_acc_1_cse_4_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
      + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "011")), 10));
  COMP_LOOP_acc_11_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
      DOWNTO 1)) + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "01")),
      9));
  COMP_LOOP_acc_1_cse_2_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
      + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "001")), 10));
  COMP_LOOP_2_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "001")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_2_acc_10_itm_10_1_1 <= COMP_LOOP_2_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_3_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "010")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_3_acc_10_itm_10_1_1 <= COMP_LOOP_3_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_4_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "011")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_4_acc_10_itm_10_1_1 <= COMP_LOOP_4_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_5_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "100")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_5_acc_10_itm_10_1_1 <= COMP_LOOP_5_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_6_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "101")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_6_acc_10_itm_10_1_1 <= COMP_LOOP_6_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_7_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "110")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_7_acc_10_itm_10_1_1 <= COMP_LOOP_7_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_8_acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 &
      STD_LOGIC_VECTOR'( "111")), 10), 11) + UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      11));
  COMP_LOOP_8_acc_10_itm_10_1_1 <= COMP_LOOP_8_acc_10_nl(10 DOWNTO 1);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_274_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(1))
      AND COMP_LOOP_tmp_nor_151_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_276_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(2))
      AND COMP_LOOP_tmp_nor_153_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_280_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(3))
      AND COMP_LOOP_tmp_nor_157_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_288_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(4))
      AND COMP_LOOP_tmp_nor_165_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_304_rgt <= (COMP_LOOP_2_tmp_lshift_ncse_sva(5))
      AND COMP_LOOP_tmp_nor_180_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_243_rgt <= (COMP_LOOP_3_tmp_lshift_ncse_sva(1))
      AND COMP_LOOP_tmp_nor_207_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_245_rgt <= (COMP_LOOP_3_tmp_lshift_ncse_sva(2))
      AND COMP_LOOP_tmp_nor_209_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_249_rgt <= (COMP_LOOP_3_tmp_lshift_ncse_sva(3))
      AND COMP_LOOP_tmp_nor_213_itm;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_257_rgt <= (COMP_LOOP_3_tmp_lshift_ncse_sva(4))
      AND COMP_LOOP_tmp_nor_220_itm;
  nor_tmp_1 <= (fsm_output(4)) AND (fsm_output(0)) AND (fsm_output(3));
  mux_tmp_6 <= MUX_s_1_2_2((fsm_output(4)), or_595_cse, fsm_output(2));
  and_dcpl_8 <= nor_399_cse AND (NOT (fsm_output(5)));
  and_779_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111"));
  or_150_cse <= (fsm_output(0)) OR (fsm_output(3));
  and_tmp_10 <= (fsm_output(4)) AND or_150_cse;
  or_tmp_105 <= (fsm_output(4)) OR and_639_cse;
  or_tmp_118 <= (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_119 <= (fsm_output(3)) OR (fsm_output(7));
  not_tmp_88 <= NOT((fsm_output(4)) OR (fsm_output(7)));
  nor_tmp_99 <= or_341_cse AND (fsm_output(7));
  mux_tmp_206 <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), or_341_cse);
  or_4050_cse <= and_640_cse OR (fsm_output(6));
  mux_tmp_293 <= MUX_s_1_2_2(and_640_cse, (fsm_output(4)), fsm_output(2));
  mux_510_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_118, fsm_output(4));
  mux_tmp_444 <= MUX_s_1_2_2(mux_510_nl, (fsm_output(7)), fsm_output(6));
  or_tmp_404 <= (fsm_output(4)) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_201_nl <= (fsm_output(4)) OR (NOT (fsm_output(7)));
  mux_tmp_656 <= MUX_s_1_2_2(or_201_nl, (fsm_output(7)), fsm_output(6));
  and_dcpl_55 <= NOT((fsm_output(1)) OR (fsm_output(5)));
  and_dcpl_57 <= nor_1674_cse AND and_dcpl_55;
  and_dcpl_58 <= NOT((fsm_output(0)) OR (fsm_output(4)));
  and_dcpl_59 <= NOT((fsm_output(7)) OR (fsm_output(3)));
  and_dcpl_60 <= and_dcpl_59 AND and_dcpl_58;
  and_dcpl_62 <= (NOT (fsm_output(1))) AND (fsm_output(5));
  and_dcpl_64 <= and_808_cse AND and_dcpl_62;
  and_dcpl_65 <= (fsm_output(7)) AND (NOT (fsm_output(3)));
  and_dcpl_66 <= and_dcpl_65 AND and_dcpl_58;
  and_tmp_29 <= (fsm_output(6)) AND and_655_cse;
  mux_tmp_720 <= MUX_s_1_2_2(and_tmp_29, and_705_cse, fsm_output(2));
  and_dcpl_72 <= (fsm_output(1)) AND (NOT (fsm_output(5)));
  and_dcpl_73 <= nor_1674_cse AND and_dcpl_72;
  and_dcpl_74 <= and_dcpl_60 AND and_dcpl_73;
  and_dcpl_75 <= (fsm_output(0)) AND (NOT (fsm_output(4)));
  and_dcpl_76 <= and_dcpl_59 AND and_dcpl_75;
  and_dcpl_77 <= and_dcpl_76 AND and_dcpl_73;
  and_dcpl_78 <= (NOT (fsm_output(6))) AND (fsm_output(2));
  and_dcpl_79 <= and_dcpl_78 AND and_dcpl_72;
  and_dcpl_80 <= (NOT (fsm_output(0))) AND (fsm_output(4));
  and_dcpl_81 <= (NOT (fsm_output(7))) AND (fsm_output(3));
  and_dcpl_82 <= and_dcpl_81 AND and_dcpl_80;
  and_dcpl_84 <= (fsm_output(0)) AND (fsm_output(4));
  and_dcpl_85 <= and_dcpl_81 AND and_dcpl_84;
  and_dcpl_86 <= and_dcpl_85 AND and_dcpl_79;
  and_dcpl_87 <= (fsm_output(1)) AND (fsm_output(5));
  and_dcpl_88 <= nor_1674_cse AND and_dcpl_87;
  and_dcpl_90 <= and_dcpl_85 AND and_dcpl_88;
  and_dcpl_91 <= and_808_cse AND and_dcpl_72;
  and_dcpl_92 <= and_dcpl_59 AND and_dcpl_80;
  and_dcpl_94 <= and_dcpl_59 AND and_dcpl_84;
  and_dcpl_95 <= and_dcpl_94 AND and_dcpl_91;
  and_dcpl_96 <= (fsm_output(6)) AND (NOT (fsm_output(2)));
  and_dcpl_97 <= and_dcpl_96 AND and_dcpl_87;
  and_dcpl_99 <= and_dcpl_94 AND and_dcpl_97;
  and_dcpl_101 <= and_763_cse AND and_dcpl_58;
  and_dcpl_103 <= and_763_cse AND and_dcpl_75;
  and_dcpl_104 <= and_dcpl_103 AND and_dcpl_79;
  and_dcpl_106 <= and_dcpl_103 AND and_dcpl_88;
  and_dcpl_108 <= and_dcpl_65 AND and_dcpl_75;
  and_dcpl_109 <= and_dcpl_108 AND and_dcpl_91;
  and_dcpl_110 <= and_dcpl_78 AND and_dcpl_55;
  and_dcpl_112 <= and_dcpl_85 AND and_dcpl_110;
  and_dcpl_113 <= nor_1674_cse AND and_dcpl_62;
  and_dcpl_115 <= and_dcpl_85 AND and_dcpl_113;
  and_dcpl_116 <= and_808_cse AND and_dcpl_55;
  and_dcpl_118 <= and_dcpl_94 AND and_dcpl_116;
  and_dcpl_119 <= and_dcpl_96 AND and_dcpl_62;
  or_tmp_491 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_495 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_497 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_501 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT and_763_cse);
  or_tmp_535 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_539 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_541 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_545 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (NOT and_763_cse);
  not_tmp_321 <= NOT((VEC_LOOP_j_10_0_sva_9_0(0)) AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_579 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_583 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_585 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_589 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT and_763_cse);
  or_tmp_623 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_627 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_629 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_633 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (NOT and_763_cse);
  not_tmp_330 <= NOT(CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_667 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_671 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_673 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_677 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT and_763_cse);
  or_tmp_711 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_715 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_717 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_721 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (NOT and_763_cse);
  or_tmp_755 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_759 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_761 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_765 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT and_763_cse);
  or_tmp_799 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_803 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_805 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_809 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (NOT and_763_cse);
  not_tmp_347 <= NOT((COMP_LOOP_acc_13_psp_sva(0)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_843 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_847 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_849 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_853 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT and_763_cse);
  or_tmp_887 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_891 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_893 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_897 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (NOT and_763_cse);
  or_tmp_931 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_935 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_937 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_941 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT and_763_cse);
  or_tmp_975 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_979 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_981 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_985 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (NOT and_763_cse);
  or_tmp_1019 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1023 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1025 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1029 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT and_763_cse);
  or_tmp_1063 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1067 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1069 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1073 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (NOT and_763_cse);
  or_tmp_1107 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1111 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1113 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1117 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT and_763_cse);
  or_tmp_1151 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1155 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1157 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1161 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001111"))
      AND and_763_cse);
  or_tmp_1195 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1199 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1201 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1205 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (NOT and_763_cse);
  not_tmp_384 <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(4)) AND (fsm_output(3)) AND
      (fsm_output(7)));
  not_tmp_388 <= NOT((COMP_LOOP_acc_10_cse_10_1_7_sva(4)) AND (fsm_output(3)) AND
      (fsm_output(7)));
  or_tmp_1239 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1243 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1245 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1249 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (NOT and_763_cse);
  or_tmp_1283 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1287 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1289 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1293 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (NOT and_763_cse);
  or_tmp_1327 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1331 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1333 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1337 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (NOT and_763_cse);
  or_tmp_1371 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1375 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1377 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1381 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (NOT and_763_cse);
  or_tmp_1415 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1419 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1421 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1425 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (NOT and_763_cse);
  or_tmp_1459 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1463 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1465 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1469 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (NOT and_763_cse);
  or_tmp_1503 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1507 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1509 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1513 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010111"))
      AND and_763_cse);
  not_tmp_414 <= NOT((COMP_LOOP_acc_13_psp_sva(2)) AND (COMP_LOOP_acc_13_psp_sva(0))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_1547 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1551 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1553 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1557 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (NOT and_763_cse);
  or_tmp_1591 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1595 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1597 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1601 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (NOT and_763_cse);
  or_tmp_1635 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1639 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1641 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1645 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (NOT and_763_cse);
  or_tmp_1679 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1683 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1685 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1689 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011011"))
      AND and_763_cse);
  or_tmp_1723 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1727 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1729 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1733 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (NOT and_763_cse);
  or_tmp_1767 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1771 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1773 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1777 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011101"))
      AND and_763_cse);
  or_tmp_1811 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1815 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1817 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1821 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011110"))
      AND and_763_cse);
  or_tmp_1855 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1859 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  or_tmp_1861 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  or_tmp_1865 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND and_763_cse);
  or_tmp_1898 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1902 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1904 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  not_tmp_452 <= NOT((COMP_LOOP_acc_1_cse_6_sva(5)) AND (fsm_output(3)) AND (fsm_output(7)));
  not_tmp_453 <= NOT((COMP_LOOP_acc_10_cse_10_1_6_sva(5)) AND (fsm_output(3)) AND
      (fsm_output(7)));
  or_tmp_1908 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR not_tmp_453;
  or_tmp_1942 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1946 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1948 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  not_tmp_458 <= NOT((COMP_LOOP_acc_10_cse_10_1_6_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(5))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_1952 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"))
      OR not_tmp_458;
  or_tmp_1986 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_1990 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_1992 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_1996 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR not_tmp_453;
  or_tmp_2030 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2034 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2036 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  not_tmp_467 <= NOT((COMP_LOOP_acc_10_cse_10_1_6_sva(1)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(0))
      AND (COMP_LOOP_acc_10_cse_10_1_6_sva(5)) AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_2040 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"))
      OR not_tmp_467;
  or_tmp_2074 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2078 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2080 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2084 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR not_tmp_453;
  or_tmp_2118 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2122 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2124 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2128 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"))
      OR not_tmp_458;
  or_tmp_2162 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2166 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2168 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2172 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR not_tmp_453;
  or_tmp_2206 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2210 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2212 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  not_tmp_484 <= NOT((COMP_LOOP_acc_10_cse_10_1_6_sva(2)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(1))
      AND (COMP_LOOP_acc_10_cse_10_1_6_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(5))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_2216 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_484;
  or_tmp_2250 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2254 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2256 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2260 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR not_tmp_453;
  or_tmp_2294 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2298 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2300 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2304 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"))
      OR not_tmp_458;
  or_tmp_2338 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2342 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2344 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2348 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR not_tmp_453;
  or_tmp_2382 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2386 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2388 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2392 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("010"))
      OR not_tmp_467;
  or_tmp_2426 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2430 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2432 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2436 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR not_tmp_453;
  or_tmp_2470 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2474 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2476 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2480 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"))
      OR not_tmp_458;
  or_tmp_2514 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2518 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2520 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2524 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR not_tmp_453;
  or_tmp_2558 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2562 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  or_tmp_2564 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  or_tmp_2567 <= (COMP_LOOP_acc_10_cse_10_1_6_sva(4)) OR (NOT((COMP_LOOP_acc_10_cse_10_1_6_sva(3))
      AND (COMP_LOOP_acc_10_cse_10_1_6_sva(2)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(1))
      AND (COMP_LOOP_acc_10_cse_10_1_6_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(5))
      AND (fsm_output(3)) AND (fsm_output(7))));
  or_tmp_2601 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2605 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2607 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  not_tmp_522 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_2611 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR not_tmp_453;
  not_tmp_523 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)) AND (fsm_output(7)));
  not_tmp_527 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_2645 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2649 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2651 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2655 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"))
      OR not_tmp_458;
  or_tmp_2689 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2693 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2695 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2699 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR not_tmp_453;
  or_tmp_2733 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2737 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2739 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2743 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("100"))
      OR not_tmp_467;
  or_tmp_2777 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2781 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2783 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2787 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR not_tmp_453;
  not_tmp_544 <= NOT((COMP_LOOP_acc_10_cse_10_1_7_sva(2)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(5))
      AND (COMP_LOOP_acc_10_cse_10_1_7_sva(4)) AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_2821 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2825 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2827 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2831 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"))
      OR not_tmp_458;
  not_tmp_549 <= NOT((COMP_LOOP_acc_10_cse_10_1_7_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      AND (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(4))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_2865 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2869 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2871 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_2875 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR not_tmp_453;
  or_tmp_2909 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2913 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  or_tmp_2915 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  or_tmp_2919 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_484;
  or_tmp_2953 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_2957 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_2959 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  not_tmp_559 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 3)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_2963 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR not_tmp_453;
  not_tmp_560 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 3)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_2997 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_3001 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_3003 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  not_tmp_565 <= NOT((COMP_LOOP_acc_1_cse_6_sva(0)) AND (COMP_LOOP_acc_1_cse_6_sva(3))
      AND (COMP_LOOP_acc_1_cse_6_sva(4)) AND (COMP_LOOP_acc_1_cse_6_sva(5)) AND (fsm_output(3))
      AND (fsm_output(7)));
  or_tmp_3007 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100"))
      OR not_tmp_458;
  or_tmp_3041 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_3045 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_3047 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_3051 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR not_tmp_453;
  not_tmp_570 <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(1)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      AND (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(4))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_3085 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_3089 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  or_tmp_3091 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  not_tmp_575 <= NOT((COMP_LOOP_acc_1_cse_6_sva(1)) AND (COMP_LOOP_acc_1_cse_6_sva(0))
      AND (COMP_LOOP_acc_1_cse_6_sva(3)) AND (COMP_LOOP_acc_1_cse_6_sva(4)) AND (COMP_LOOP_acc_1_cse_6_sva(5))
      AND (fsm_output(3)) AND (fsm_output(7)));
  or_tmp_3094 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("110"))
      OR not_tmp_467;
  or_tmp_3128 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_3132 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  or_tmp_3134 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_tmp_3138 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR not_tmp_453;
  or_tmp_3172 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_3176 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  or_tmp_3178 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  or_tmp_3182 <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1110"))))
      OR not_tmp_458;
  or_tmp_3215 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_tmp_3219 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  or_tmp_3221 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  or_tmp_3225 <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))))
      OR not_tmp_453;
  or_tmp_3258 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7))));
  or_tmp_3262 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  or_tmp_3264 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  nor_tmp_306 <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)) AND (fsm_output(7));
  nor_tmp_307 <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)) AND (fsm_output(7));
  and_dcpl_258 <= and_dcpl_60 AND and_dcpl_110;
  and_dcpl_259 <= and_dcpl_76 AND and_dcpl_110;
  and_dcpl_260 <= and_dcpl_60 AND and_dcpl_79;
  and_dcpl_261 <= and_dcpl_76 AND and_dcpl_79;
  and_dcpl_262 <= and_dcpl_81 AND and_dcpl_58;
  and_dcpl_263 <= and_dcpl_262 AND and_dcpl_57;
  and_dcpl_264 <= and_dcpl_81 AND and_dcpl_75;
  and_dcpl_265 <= and_dcpl_264 AND and_dcpl_57;
  and_dcpl_268 <= not_tmp_88 AND nor_1683_cse;
  mux_tmp_2924 <= MUX_s_1_2_2((NOT and_763_cse), or_tmp_118, fsm_output(4));
  or_tmp_3717 <= (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_tmp_2927 <= MUX_s_1_2_2(or_tmp_3717, or_tmp_119, fsm_output(4));
  or_tmp_3718 <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(7));
  and_dcpl_340 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  or_tmp_3721 <= (NOT (fsm_output(4))) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  and_dcpl_343 <= and_dcpl_60 AND and_dcpl_113;
  and_dcpl_344 <= and_dcpl_78 AND and_dcpl_62;
  and_dcpl_346 <= and_dcpl_82 AND and_dcpl_344;
  and_dcpl_347 <= and_dcpl_96 AND and_dcpl_55;
  and_dcpl_349 <= and_dcpl_82 AND and_dcpl_347;
  and_dcpl_351 <= and_dcpl_92 AND and_dcpl_64;
  and_dcpl_353 <= and_dcpl_65 AND and_dcpl_80;
  and_dcpl_354 <= and_dcpl_353 AND and_dcpl_57;
  and_dcpl_355 <= and_763_cse AND and_dcpl_80;
  and_dcpl_357 <= and_dcpl_101 AND and_dcpl_344;
  and_dcpl_359 <= and_dcpl_101 AND and_dcpl_347;
  mux_522_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(4));
  mux_3004_nl <= MUX_s_1_2_2(and_735_cse, mux_522_nl, fsm_output(0));
  nand_tmp_142 <= NOT((fsm_output(3)) AND (NOT mux_3004_nl));
  or_3843_nl <= (fsm_output(0)) OR (NOT and_735_cse);
  mux_tmp_2939 <= MUX_s_1_2_2(or_364_cse, or_3843_nl, fsm_output(3));
  or_tmp_3734 <= (fsm_output(5)) OR (NOT (fsm_output(1)));
  and_dcpl_365 <= (NOT (fsm_output(3))) AND (fsm_output(0));
  or_dcpl_122 <= (fsm_output(6)) OR (fsm_output(2)) OR or_tmp_3734;
  or_dcpl_125 <= or_tmp_119 OR (fsm_output(0)) OR (fsm_output(4)) OR or_dcpl_122;
  mux_tmp_2953 <= MUX_s_1_2_2(and_dcpl_60, and_655_cse, fsm_output(6));
  mux_tmp_2955 <= MUX_s_1_2_2((NOT or_477_cse), and_655_cse, fsm_output(6));
  mux_tmp_2956 <= MUX_s_1_2_2(mux_tmp_2955, and_tmp_29, fsm_output(2));
  mux_3021_nl <= MUX_s_1_2_2(mux_tmp_2953, and_78_cse, fsm_output(2));
  mux_3024_nl <= MUX_s_1_2_2(mux_tmp_2956, mux_3021_nl, fsm_output(1));
  mux_3025_itm <= MUX_s_1_2_2(mux_3024_nl, and_705_cse, fsm_output(5));
  mux_tmp_2959 <= MUX_s_1_2_2((NOT or_595_cse), and_640_cse, fsm_output(6));
  mux_tmp_2960 <= MUX_s_1_2_2(mux_tmp_2959, and_677_cse, fsm_output(2));
  mux_tmp_2961 <= MUX_s_1_2_2((NOT or_4007_cse), and_640_cse, fsm_output(6));
  mux_tmp_2965 <= MUX_s_1_2_2((NOT or_595_cse), (fsm_output(4)), fsm_output(6));
  mux_tmp_2966 <= MUX_s_1_2_2(mux_tmp_2959, mux_tmp_2965, fsm_output(2));
  mux_3034_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), and_640_cse, fsm_output(6));
  mux_tmp_2968 <= MUX_s_1_2_2(mux_3034_nl, mux_tmp_2965, fsm_output(2));
  and_dcpl_370 <= and_dcpl_264 AND and_dcpl_113;
  mux_tmp_2971 <= MUX_s_1_2_2(mux_tmp_2959, and_673_cse, fsm_output(2));
  mux_3041_nl <= MUX_s_1_2_2(and_dcpl_365, (fsm_output(3)), fsm_output(4));
  or_tmp_3744 <= (fsm_output(6)) OR mux_3041_nl;
  mux_tmp_2975 <= MUX_s_1_2_2((fsm_output(6)), or_tmp_3744, fsm_output(2));
  or_tmp_3746 <= (fsm_output(6)) OR (NOT((fsm_output(4)) OR (NOT and_639_cse)));
  mux_tmp_2976 <= MUX_s_1_2_2(or_tmp_3746, (fsm_output(6)), fsm_output(2));
  and_dcpl_375 <= and_dcpl_264 AND and_dcpl_88;
  or_tmp_3747 <= (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(3));
  and_dcpl_377 <= and_dcpl_78 AND and_dcpl_87;
  and_dcpl_382 <= and_dcpl_94 AND and_dcpl_377;
  or_3880_nl <= (fsm_output(6)) OR nor_398_cse;
  mux_3057_nl <= MUX_s_1_2_2((fsm_output(6)), or_3880_nl, fsm_output(2));
  mux_3058_itm <= MUX_s_1_2_2(mux_tmp_2976, mux_3057_nl, fsm_output(1));
  and_dcpl_384 <= and_dcpl_85 AND and_dcpl_57;
  mux_tmp_2993 <= MUX_s_1_2_2(or_4050_cse, or_tmp_3744, fsm_output(2));
  mux_tmp_2994 <= MUX_s_1_2_2(or_tmp_3746, or_4050_cse, fsm_output(2));
  or_tmp_3757 <= (NOT((NOT (fsm_output(0))) OR (fsm_output(3)))) OR (fsm_output(7));
  or_tmp_3760 <= and_639_cse OR (fsm_output(7));
  or_3887_nl <= (fsm_output(4)) OR (NOT or_tmp_3760);
  mux_tmp_3001 <= MUX_s_1_2_2(or_3887_nl, (fsm_output(7)), fsm_output(6));
  mux_3069_nl <= MUX_s_1_2_2(mux_tmp_3001, mux_tmp_656, fsm_output(2));
  or_3884_nl <= (fsm_output(4)) OR (NOT or_tmp_3757);
  mux_3065_nl <= MUX_s_1_2_2(or_3884_nl, (fsm_output(7)), fsm_output(6));
  mux_3067_nl <= MUX_s_1_2_2(mux_tmp_656, mux_3065_nl, fsm_output(2));
  mux_tmp_3003 <= MUX_s_1_2_2(mux_3069_nl, mux_3067_nl, fsm_output(1));
  mux_3075_nl <= MUX_s_1_2_2((NOT or_tmp_3757), or_tmp_118, fsm_output(4));
  mux_tmp_3009 <= MUX_s_1_2_2(mux_3075_nl, (fsm_output(7)), fsm_output(6));
  mux_tmp_3012 <= MUX_s_1_2_2(mux_tmp_444, mux_tmp_3009, fsm_output(2));
  mux_tmp_3013 <= MUX_s_1_2_2(mux_tmp_3001, mux_tmp_444, fsm_output(2));
  mux_tmp_3016 <= MUX_s_1_2_2(and_dcpl_59, (fsm_output(7)), or_341_cse);
  and_dcpl_387 <= and_dcpl_264 AND and_dcpl_79;
  or_tmp_3773 <= nor_1744_cse OR (fsm_output(7));
  and_dcpl_388 <= and_dcpl_94 AND and_dcpl_79;
  mux_tmp_3042 <= MUX_s_1_2_2(mux_tmp_2953, and_705_cse, fsm_output(2));
  and_tmp_31 <= (fsm_output(6)) AND (fsm_output(4)) AND or_150_cse;
  or_3906_nl <= (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0))
      OR (fsm_output(3));
  mux_3114_itm <= MUX_s_1_2_2(or_tmp_3747, or_3906_nl, fsm_output(1));
  mux_tmp_3049 <= MUX_s_1_2_2(mux_tmp_2961, and_673_cse, fsm_output(2));
  mux_3117_nl <= MUX_s_1_2_2(mux_tmp_2959, and_tmp_31, fsm_output(2));
  mux_3118_nl <= MUX_s_1_2_2(mux_3117_nl, mux_tmp_3049, fsm_output(1));
  mux_3119_nl <= MUX_s_1_2_2(mux_3118_nl, (fsm_output(6)), fsm_output(5));
  and_dcpl_390 <= NOT(mux_3119_nl OR (fsm_output(7)));
  mux_67_nl <= MUX_s_1_2_2(nor_tmp_1, and_640_cse, or_359_cse);
  mux_3122_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_67_nl), fsm_output(5));
  and_dcpl_392 <= mux_3122_nl AND nor_399_cse;
  and_dcpl_396 <= mux_221_cse AND and_dcpl_8;
  mux_3129_nl <= MUX_s_1_2_2(mux_221_cse, (NOT and_779_cse), fsm_output(5));
  and_dcpl_399 <= mux_3129_nl AND nor_399_cse;
  mux_3133_nl <= MUX_s_1_2_2(mux_tmp_2961, and_677_cse, fsm_output(2));
  mux_3134_nl <= MUX_s_1_2_2(mux_tmp_2960, mux_3133_nl, fsm_output(1));
  mux_3135_nl <= MUX_s_1_2_2(mux_3134_nl, (fsm_output(6)), fsm_output(5));
  and_dcpl_402 <= NOT(mux_3135_nl OR (fsm_output(7)));
  nor_1425_nl <= NOT((fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_tmp_3069 <= MUX_s_1_2_2(nor_1425_nl, (fsm_output(7)), or_341_cse);
  mux_tmp_3070 <= MUX_s_1_2_2(mux_tmp_3069, and_736_cse, fsm_output(2));
  mux_tmp_3078 <= MUX_s_1_2_2(mux_tmp_3016, nor_tmp_99, fsm_output(2));
  mux_3148_nl <= MUX_s_1_2_2((NOT mux_3114_itm), mux_180_cse, fsm_output(5));
  and_dcpl_403 <= NOT(mux_3148_nl OR (fsm_output(7)));
  mux_210_nl <= MUX_s_1_2_2(and_640_cse, and_tmp_10, and_507_cse);
  mux_3150_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_210_nl), fsm_output(5));
  and_dcpl_404 <= mux_3150_nl AND nor_399_cse;
  mux_214_nl <= MUX_s_1_2_2(or_tmp_105, or_595_cse, fsm_output(2));
  mux_215_nl <= MUX_s_1_2_2(mux_tmp_6, mux_214_nl, fsm_output(1));
  mux_3156_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_215_nl), fsm_output(5));
  and_dcpl_406 <= mux_3156_nl AND nor_399_cse;
  mux_217_nl <= MUX_s_1_2_2(or_tmp_105, or_595_cse, or_359_cse);
  mux_3158_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_217_nl), fsm_output(5));
  and_dcpl_407 <= mux_3158_nl AND nor_399_cse;
  mux_tmp_3098 <= MUX_s_1_2_2(and_dcpl_60, (fsm_output(7)), fsm_output(6));
  mux_tmp_3100 <= MUX_s_1_2_2((NOT or_477_cse), (fsm_output(7)), fsm_output(6));
  mux_tmp_3101 <= MUX_s_1_2_2(mux_tmp_3100, and_705_cse, fsm_output(2));
  mux_3166_nl <= MUX_s_1_2_2(mux_tmp_3098, and_705_cse, fsm_output(2));
  mux_tmp_3102 <= MUX_s_1_2_2(mux_tmp_3101, mux_3166_nl, fsm_output(1));
  mux_3173_nl <= MUX_s_1_2_2(mux_tmp_3069, nor_tmp_99, fsm_output(2));
  mux_3174_nl <= MUX_s_1_2_2(mux_tmp_3078, mux_3173_nl, fsm_output(1));
  mux_3175_itm <= MUX_s_1_2_2(mux_3174_nl, (fsm_output(7)), fsm_output(5));
  mux_3176_nl <= MUX_s_1_2_2(nor_tmp_1, and_640_cse, fsm_output(2));
  mux_3177_nl <= MUX_s_1_2_2(and_779_cse, mux_3176_nl, fsm_output(1));
  mux_3178_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_3177_nl), fsm_output(5));
  and_dcpl_410 <= mux_3178_nl AND nor_399_cse;
  mux_3179_nl <= MUX_s_1_2_2(or_4007_cse, (NOT nor_tmp_1), fsm_output(2));
  mux_3180_nl <= MUX_s_1_2_2(or_80_cse, mux_3179_nl, fsm_output(1));
  and_dcpl_411 <= mux_3180_nl AND and_dcpl_8;
  mux_3184_nl <= MUX_s_1_2_2(mux_tmp_2956, mux_tmp_3042, fsm_output(1));
  mux_3185_itm <= MUX_s_1_2_2(mux_3184_nl, and_705_cse, fsm_output(5));
  mux_tmp_3119 <= MUX_s_1_2_2(nor_tmp_99, and_736_cse, fsm_output(2));
  mux_3187_itm <= MUX_s_1_2_2(mux_tmp_3102, mux_tmp_3119, fsm_output(5));
  nor_1524_nl <= NOT((fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(4))
      OR (fsm_output(7)));
  nor_409_nl <= NOT((fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0))
      OR (fsm_output(3)) OR (fsm_output(7)));
  not_tmp_811 <= MUX_s_1_2_2(nor_1524_nl, nor_409_nl, fsm_output(1));
  mux_3199_nl <= MUX_s_1_2_2(mux_tmp_2953, and_tmp_29, fsm_output(2));
  mux_tmp_3133 <= MUX_s_1_2_2(mux_tmp_2956, mux_3199_nl, fsm_output(1));
  mux_3201_itm <= MUX_s_1_2_2(mux_tmp_3133, and_705_cse, fsm_output(5));
  or_tmp_3801 <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(3));
  and_tmp_33 <= (fsm_output(6)) AND or_595_cse;
  and_dcpl_421 <= and_dcpl_85 AND and_dcpl_73;
  mux_tmp_3169 <= MUX_s_1_2_2(or_tmp_3717, or_tmp_118, fsm_output(4));
  mux_tmp_3193 <= MUX_s_1_2_2((NOT (fsm_output(7))), and_655_cse, fsm_output(6));
  nor_400_nl <= NOT((NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(3))) OR (fsm_output(4))))
      OR (fsm_output(7)));
  mux_3262_nl <= MUX_s_1_2_2(nor_400_nl, and_655_cse, fsm_output(6));
  mux_tmp_3196 <= MUX_s_1_2_2(mux_3262_nl, mux_tmp_3193, fsm_output(2));
  and_tmp_35 <= (fsm_output(5)) AND mux_297_cse;
  mux_tmp_3210 <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), or_595_cse);
  and_tmp_36 <= (fsm_output(6)) AND mux_tmp_3210;
  mux_tmp_3213 <= MUX_s_1_2_2(or_tmp_3717, (fsm_output(7)), fsm_output(4));
  mux_tmp_3214 <= MUX_s_1_2_2((NOT or_477_cse), mux_tmp_3213, fsm_output(6));
  nor_1474_nl <= NOT(and_640_cse OR (fsm_output(7)));
  mux_tmp_3218 <= MUX_s_1_2_2(nor_1474_nl, (fsm_output(7)), fsm_output(6));
  mux_75_nl <= MUX_s_1_2_2(or_595_cse, or_4007_cse, fsm_output(2));
  mux_3305_itm <= MUX_s_1_2_2(mux_75_nl, or_80_cse, fsm_output(1));
  or_dcpl_134 <= or_tmp_119 OR (NOT (fsm_output(0))) OR (fsm_output(4));
  nor_1709_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")));
  nor_1710_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  mux_3314_nl <= MUX_s_1_2_2(nor_1709_nl, nor_1710_nl, fsm_output(1));
  and_dcpl_432 <= mux_3314_nl AND (NOT (fsm_output(7))) AND and_dcpl_75 AND nor_1683_cse;
  or_tmp_3833 <= (fsm_output(4)) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  nor_tmp_391 <= (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(7));
  mux_tmp_3280 <= MUX_s_1_2_2((NOT or_477_cse), and_735_cse, fsm_output(6));
  not_tmp_868 <= NOT((fsm_output(4)) OR or_tmp_3760);
  or_dcpl_150 <= or_dcpl_134 OR (fsm_output(6)) OR (NOT (fsm_output(2))) OR or_tmp_3734;
  mux_3354_nl <= MUX_s_1_2_2(and_dcpl_59, and_763_cse, fsm_output(4));
  mux_tmp_3288 <= MUX_s_1_2_2(mux_3354_nl, (fsm_output(7)), fsm_output(6));
  STAGE_LOOP_i_3_0_sva_mx0c1 <= and_dcpl_66 AND and_dcpl_64;
  VEC_LOOP_j_10_0_sva_9_0_mx0c0 <= and_dcpl_76 AND and_dcpl_57;
  mux_3318_nl <= MUX_s_1_2_2(mux_tmp_2927, or_tmp_3833, fsm_output(6));
  mux_3317_nl <= MUX_s_1_2_2((NOT nor_tmp_391), or_tmp_3721, fsm_output(6));
  mux_3319_nl <= MUX_s_1_2_2(mux_3318_nl, mux_3317_nl, fsm_output(2));
  or_3973_nl <= (fsm_output(6)) OR (NOT nor_tmp_391);
  mux_3315_nl <= MUX_s_1_2_2(or_tmp_3833, or_477_cse, fsm_output(6));
  mux_3316_nl <= MUX_s_1_2_2(or_3973_nl, mux_3315_nl, fsm_output(2));
  mux_3320_nl <= MUX_s_1_2_2(mux_3319_nl, mux_3316_nl, fsm_output(5));
  COMP_LOOP_1_acc_8_itm_mx0c4 <= (NOT mux_3320_nl) AND and_dcpl_340;
  mux_3340_nl <= MUX_s_1_2_2(mux_3305_itm, (NOT mux_tmp_6), fsm_output(5));
  and_474_tmp <= mux_3340_nl AND nor_399_cse;
  mux_104_nl <= MUX_s_1_2_2((NOT or_595_cse), or_595_cse, fsm_output(6));
  mux_3342_nl <= MUX_s_1_2_2(mux_104_nl, and_tmp_33, and_507_cse);
  mux_3343_nl <= MUX_s_1_2_2(mux_3342_nl, (fsm_output(6)), fsm_output(5));
  nor_1579_tmp <= NOT(mux_3343_nl OR (fsm_output(7)));
  mux_3345_nl <= MUX_s_1_2_2(or_4057_cse, or_tmp_3801, and_507_cse);
  mux_3344_nl <= MUX_s_1_2_2(and_tmp_33, (fsm_output(6)), fsm_output(2));
  mux_3346_nl <= MUX_s_1_2_2(mux_3345_nl, (NOT mux_3344_nl), fsm_output(5));
  and_476_tmp <= mux_3346_nl AND (NOT (fsm_output(7)));
  nor_tmp_396 <= NOT((NOT(or_595_cse OR CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"))))
      OR (fsm_output(7)));
  and_102_nl <= ((fsm_output(7)) XOR (fsm_output(4))) AND ((fsm_output(3)) XOR (fsm_output(6)))
      AND (NOT (fsm_output(1))) AND ((fsm_output(2)) XOR (fsm_output(5))) AND (fsm_output(0));
  vec_rsc_0_0_i_d_d_pff <= MUX_v_64_2_2(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z,
      COMP_LOOP_1_acc_8_itm, and_102_nl);
  and_114_nl <= and_dcpl_82 AND and_dcpl_79;
  and_120_nl <= and_dcpl_82 AND and_dcpl_88;
  and_124_nl <= and_dcpl_92 AND and_dcpl_91;
  and_129_nl <= and_dcpl_92 AND and_dcpl_97;
  and_133_nl <= and_dcpl_101 AND and_dcpl_79;
  and_136_nl <= and_dcpl_101 AND and_dcpl_88;
  and_138_nl <= and_dcpl_66 AND and_dcpl_91;
  vec_rsc_0_0_i_radr_d_pff <= MUX1HOT_v_4_16_2((COMP_LOOP_1_acc_10_itm_10_1_1(9 DOWNTO
      6)), (COMP_LOOP_acc_psp_sva(6 DOWNTO 3)), (COMP_LOOP_acc_1_cse_2_sva(9 DOWNTO
      6)), (COMP_LOOP_acc_10_cse_10_1_2_sva(9 DOWNTO 6)), (COMP_LOOP_acc_11_psp_sva(8
      DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_3_sva(9 DOWNTO 6)), (COMP_LOOP_acc_1_cse_4_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_10_cse_10_1_4_sva(9 DOWNTO 6)), (COMP_LOOP_acc_13_psp_sva(7
      DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_5_sva(9 DOWNTO 6)), (COMP_LOOP_acc_1_cse_6_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_10_cse_10_1_6_sva(9 DOWNTO 6)), (COMP_LOOP_acc_14_psp_sva(8
      DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_7_sva(9 DOWNTO 6)), (COMP_LOOP_acc_1_cse_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_10_cse_10_1_sva(9 DOWNTO 6)), STD_LOGIC_VECTOR'(
      and_dcpl_74 & and_dcpl_77 & and_114_nl & and_dcpl_86 & and_120_nl & and_dcpl_90
      & and_124_nl & and_dcpl_95 & and_129_nl & and_dcpl_99 & and_133_nl & and_dcpl_104
      & and_136_nl & and_dcpl_106 & and_138_nl & and_dcpl_109));
  and_142_nl <= and_dcpl_82 AND and_dcpl_110;
  and_145_nl <= and_dcpl_82 AND and_dcpl_113;
  and_148_nl <= and_dcpl_92 AND and_dcpl_116;
  and_151_nl <= and_dcpl_92 AND and_dcpl_119;
  and_152_nl <= and_dcpl_94 AND and_dcpl_119;
  and_153_nl <= and_dcpl_101 AND and_dcpl_110;
  and_154_nl <= and_dcpl_103 AND and_dcpl_110;
  and_155_nl <= and_dcpl_101 AND and_dcpl_113;
  and_156_nl <= and_dcpl_103 AND and_dcpl_113;
  and_157_nl <= and_dcpl_66 AND and_dcpl_116;
  and_158_nl <= and_dcpl_108 AND and_dcpl_116;
  and_159_nl <= and_dcpl_66 AND and_dcpl_119;
  and_160_nl <= and_dcpl_108 AND and_dcpl_119;
  vec_rsc_0_0_i_wadr_d_pff <= MUX1HOT_v_4_16_2((COMP_LOOP_acc_10_cse_10_1_1_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_psp_sva(6 DOWNTO 3)), (COMP_LOOP_acc_10_cse_10_1_2_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_1_cse_2_sva(9 DOWNTO 6)), (COMP_LOOP_acc_10_cse_10_1_3_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_11_psp_sva(8 DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_4_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_1_cse_4_sva(9 DOWNTO 6)), (COMP_LOOP_acc_10_cse_10_1_5_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_13_psp_sva(7 DOWNTO 4)), (COMP_LOOP_acc_10_cse_10_1_6_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_1_cse_6_sva(9 DOWNTO 6)), (COMP_LOOP_acc_10_cse_10_1_7_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_14_psp_sva(8 DOWNTO 5)), (COMP_LOOP_acc_10_cse_10_1_sva(9
      DOWNTO 6)), (COMP_LOOP_acc_1_cse_sva(9 DOWNTO 6)), STD_LOGIC_VECTOR'( and_142_nl
      & and_dcpl_112 & and_145_nl & and_dcpl_115 & and_148_nl & and_dcpl_118 & and_151_nl
      & and_152_nl & and_153_nl & and_154_nl & and_155_nl & and_156_nl & and_157_nl
      & and_158_nl & and_159_nl & and_160_nl));
  nor_1414_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT and_763_cse));
  nor_1415_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_802_nl <= MUX_s_1_2_2(nor_1414_nl, nor_1415_nl, fsm_output(0));
  nor_1416_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1417_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_801_nl <= MUX_s_1_2_2(nor_1416_nl, nor_1417_nl, fsm_output(0));
  mux_803_nl <= MUX_s_1_2_2(mux_802_nl, mux_801_nl, fsm_output(4));
  nor_1418_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1419_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_799_nl <= MUX_s_1_2_2(nor_1418_nl, nor_1419_nl, fsm_output(0));
  nor_1420_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1421_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_798_nl <= MUX_s_1_2_2(nor_1420_nl, nor_1421_nl, fsm_output(0));
  mux_800_nl <= MUX_s_1_2_2(mux_799_nl, mux_798_nl, fsm_output(4));
  mux_804_nl <= MUX_s_1_2_2(mux_803_nl, mux_800_nl, fsm_output(6));
  nand_469_nl <= NOT((fsm_output(2)) AND mux_804_nl);
  or_615_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT and_763_cse);
  mux_795_nl <= MUX_s_1_2_2(or_tmp_501, or_615_nl, fsm_output(0));
  or_612_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_794_nl <= MUX_s_1_2_2(or_tmp_497, or_612_nl, fsm_output(0));
  mux_796_nl <= MUX_s_1_2_2(mux_795_nl, mux_794_nl, fsm_output(4));
  or_609_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_792_nl <= MUX_s_1_2_2(or_tmp_495, or_609_nl, fsm_output(0));
  or_606_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_791_nl <= MUX_s_1_2_2(or_tmp_491, or_606_nl, fsm_output(0));
  mux_793_nl <= MUX_s_1_2_2(mux_792_nl, mux_791_nl, fsm_output(4));
  mux_797_nl <= MUX_s_1_2_2(mux_796_nl, mux_793_nl, fsm_output(6));
  or_4142_nl <= (fsm_output(2)) OR mux_797_nl;
  mux_805_nl <= MUX_s_1_2_2(nand_469_nl, or_4142_nl, fsm_output(5));
  vec_rsc_0_0_i_we_d_pff <= NOT(mux_805_nl OR (fsm_output(1)));
  or_648_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_647_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_818_nl <= MUX_s_1_2_2(or_648_nl, or_647_nl, fsm_output(0));
  or_649_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_818_nl;
  or_645_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")) OR (NOT and_763_cse);
  mux_815_nl <= MUX_s_1_2_2(or_645_nl, or_tmp_501, fsm_output(0));
  or_643_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_814_nl <= MUX_s_1_2_2(or_643_nl, or_tmp_497, fsm_output(0));
  mux_816_nl <= MUX_s_1_2_2(mux_815_nl, mux_814_nl, fsm_output(4));
  or_642_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_812_nl <= MUX_s_1_2_2(or_642_nl, or_tmp_495, fsm_output(0));
  or_640_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_811_nl <= MUX_s_1_2_2(or_640_nl, or_tmp_491, fsm_output(0));
  mux_813_nl <= MUX_s_1_2_2(mux_812_nl, mux_811_nl, fsm_output(4));
  mux_817_nl <= MUX_s_1_2_2(mux_816_nl, mux_813_nl, fsm_output(6));
  mux_819_nl <= MUX_s_1_2_2(or_649_nl, mux_817_nl, fsm_output(2));
  or_638_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_636_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT and_763_cse);
  mux_808_nl <= MUX_s_1_2_2(or_638_nl, or_636_nl, fsm_output(0));
  or_634_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_633_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_807_nl <= MUX_s_1_2_2(or_634_nl, or_633_nl, fsm_output(0));
  mux_809_nl <= MUX_s_1_2_2(mux_808_nl, mux_807_nl, fsm_output(4));
  nor_1412_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1413_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_806_nl <= MUX_s_1_2_2(nor_1412_nl, nor_1413_nl, fsm_output(0));
  nand_15_nl <= NOT((fsm_output(4)) AND mux_806_nl);
  mux_810_nl <= MUX_s_1_2_2(mux_809_nl, nand_15_nl, fsm_output(6));
  or_639_nl <= (fsm_output(2)) OR mux_810_nl;
  mux_820_nl <= MUX_s_1_2_2(mux_819_nl, or_639_nl, fsm_output(5));
  vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_820_nl) AND (fsm_output(1));
  nor_1403_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (NOT and_763_cse));
  nor_1404_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_832_nl <= MUX_s_1_2_2(nor_1403_nl, nor_1404_nl, fsm_output(0));
  nor_1405_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1406_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_831_nl <= MUX_s_1_2_2(nor_1405_nl, nor_1406_nl, fsm_output(0));
  mux_833_nl <= MUX_s_1_2_2(mux_832_nl, mux_831_nl, fsm_output(4));
  nor_1407_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1408_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_829_nl <= MUX_s_1_2_2(nor_1407_nl, nor_1408_nl, fsm_output(0));
  nor_1409_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1410_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_828_nl <= MUX_s_1_2_2(nor_1409_nl, nor_1410_nl, fsm_output(0));
  mux_830_nl <= MUX_s_1_2_2(mux_829_nl, mux_828_nl, fsm_output(4));
  mux_834_nl <= MUX_s_1_2_2(mux_833_nl, mux_830_nl, fsm_output(6));
  nand_468_nl <= NOT((fsm_output(2)) AND mux_834_nl);
  or_659_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (NOT and_763_cse);
  mux_825_nl <= MUX_s_1_2_2(or_tmp_545, or_659_nl, fsm_output(0));
  or_656_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_824_nl <= MUX_s_1_2_2(or_tmp_541, or_656_nl, fsm_output(0));
  mux_826_nl <= MUX_s_1_2_2(mux_825_nl, mux_824_nl, fsm_output(4));
  or_653_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_822_nl <= MUX_s_1_2_2(or_tmp_539, or_653_nl, fsm_output(0));
  or_650_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_821_nl <= MUX_s_1_2_2(or_tmp_535, or_650_nl, fsm_output(0));
  mux_823_nl <= MUX_s_1_2_2(mux_822_nl, mux_821_nl, fsm_output(4));
  mux_827_nl <= MUX_s_1_2_2(mux_826_nl, mux_823_nl, fsm_output(6));
  or_4141_nl <= (fsm_output(2)) OR mux_827_nl;
  mux_835_nl <= MUX_s_1_2_2(nand_468_nl, or_4141_nl, fsm_output(5));
  vec_rsc_0_1_i_we_d_pff <= NOT(mux_835_nl OR (fsm_output(1)));
  or_692_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_691_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_848_nl <= MUX_s_1_2_2(or_692_nl, or_691_nl, fsm_output(0));
  or_693_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_848_nl;
  or_689_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000001")) OR (NOT and_763_cse);
  mux_845_nl <= MUX_s_1_2_2(or_689_nl, or_tmp_545, fsm_output(0));
  or_687_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000001")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_844_nl <= MUX_s_1_2_2(or_687_nl, or_tmp_541, fsm_output(0));
  mux_846_nl <= MUX_s_1_2_2(mux_845_nl, mux_844_nl, fsm_output(4));
  or_686_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000001")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_842_nl <= MUX_s_1_2_2(or_686_nl, or_tmp_539, fsm_output(0));
  or_684_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000001")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_841_nl <= MUX_s_1_2_2(or_684_nl, or_tmp_535, fsm_output(0));
  mux_843_nl <= MUX_s_1_2_2(mux_842_nl, mux_841_nl, fsm_output(4));
  mux_847_nl <= MUX_s_1_2_2(mux_846_nl, mux_843_nl, fsm_output(6));
  mux_849_nl <= MUX_s_1_2_2(or_693_nl, mux_847_nl, fsm_output(2));
  or_682_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_680_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (NOT and_763_cse);
  mux_838_nl <= MUX_s_1_2_2(or_682_nl, or_680_nl, fsm_output(0));
  or_678_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_677_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_837_nl <= MUX_s_1_2_2(or_678_nl, or_677_nl, fsm_output(0));
  mux_839_nl <= MUX_s_1_2_2(mux_838_nl, mux_837_nl, fsm_output(4));
  nor_1401_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1402_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_836_nl <= MUX_s_1_2_2(nor_1401_nl, nor_1402_nl, fsm_output(0));
  nand_17_nl <= NOT((fsm_output(4)) AND mux_836_nl);
  mux_840_nl <= MUX_s_1_2_2(mux_839_nl, nand_17_nl, fsm_output(6));
  or_683_nl <= (fsm_output(2)) OR mux_840_nl;
  mux_850_nl <= MUX_s_1_2_2(mux_849_nl, or_683_nl, fsm_output(5));
  vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_850_nl) AND (fsm_output(1));
  nor_1392_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT and_763_cse));
  nor_1393_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_862_nl <= MUX_s_1_2_2(nor_1392_nl, nor_1393_nl, fsm_output(0));
  nor_1394_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1395_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_861_nl <= MUX_s_1_2_2(nor_1394_nl, nor_1395_nl, fsm_output(0));
  mux_863_nl <= MUX_s_1_2_2(mux_862_nl, mux_861_nl, fsm_output(4));
  nor_1396_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1397_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_859_nl <= MUX_s_1_2_2(nor_1396_nl, nor_1397_nl, fsm_output(0));
  nor_1398_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1399_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_858_nl <= MUX_s_1_2_2(nor_1398_nl, nor_1399_nl, fsm_output(0));
  mux_860_nl <= MUX_s_1_2_2(mux_859_nl, mux_858_nl, fsm_output(4));
  mux_864_nl <= MUX_s_1_2_2(mux_863_nl, mux_860_nl, fsm_output(6));
  nand_467_nl <= NOT((fsm_output(2)) AND mux_864_nl);
  or_703_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT and_763_cse);
  mux_855_nl <= MUX_s_1_2_2(or_tmp_589, or_703_nl, fsm_output(0));
  or_700_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_854_nl <= MUX_s_1_2_2(or_tmp_585, or_700_nl, fsm_output(0));
  mux_856_nl <= MUX_s_1_2_2(mux_855_nl, mux_854_nl, fsm_output(4));
  or_697_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_852_nl <= MUX_s_1_2_2(or_tmp_583, or_697_nl, fsm_output(0));
  or_694_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_851_nl <= MUX_s_1_2_2(or_tmp_579, or_694_nl, fsm_output(0));
  mux_853_nl <= MUX_s_1_2_2(mux_852_nl, mux_851_nl, fsm_output(4));
  mux_857_nl <= MUX_s_1_2_2(mux_856_nl, mux_853_nl, fsm_output(6));
  or_4140_nl <= (fsm_output(2)) OR mux_857_nl;
  mux_865_nl <= MUX_s_1_2_2(nand_467_nl, or_4140_nl, fsm_output(5));
  vec_rsc_0_2_i_we_d_pff <= NOT(mux_865_nl OR (fsm_output(1)));
  or_736_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_735_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_878_nl <= MUX_s_1_2_2(or_736_nl, or_735_nl, fsm_output(0));
  or_737_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_878_nl;
  or_733_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000010")) OR (NOT and_763_cse);
  mux_875_nl <= MUX_s_1_2_2(or_733_nl, or_tmp_589, fsm_output(0));
  or_731_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000010")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_874_nl <= MUX_s_1_2_2(or_731_nl, or_tmp_585, fsm_output(0));
  mux_876_nl <= MUX_s_1_2_2(mux_875_nl, mux_874_nl, fsm_output(4));
  or_730_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000010")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_872_nl <= MUX_s_1_2_2(or_730_nl, or_tmp_583, fsm_output(0));
  or_728_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000010")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_871_nl <= MUX_s_1_2_2(or_728_nl, or_tmp_579, fsm_output(0));
  mux_873_nl <= MUX_s_1_2_2(mux_872_nl, mux_871_nl, fsm_output(4));
  mux_877_nl <= MUX_s_1_2_2(mux_876_nl, mux_873_nl, fsm_output(6));
  mux_879_nl <= MUX_s_1_2_2(or_737_nl, mux_877_nl, fsm_output(2));
  or_726_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_724_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT and_763_cse);
  mux_868_nl <= MUX_s_1_2_2(or_726_nl, or_724_nl, fsm_output(0));
  or_722_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_721_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_867_nl <= MUX_s_1_2_2(or_722_nl, or_721_nl, fsm_output(0));
  mux_869_nl <= MUX_s_1_2_2(mux_868_nl, mux_867_nl, fsm_output(4));
  nor_1390_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1391_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_866_nl <= MUX_s_1_2_2(nor_1390_nl, nor_1391_nl, fsm_output(0));
  nand_19_nl <= NOT((fsm_output(4)) AND mux_866_nl);
  mux_870_nl <= MUX_s_1_2_2(mux_869_nl, nand_19_nl, fsm_output(6));
  or_727_nl <= (fsm_output(2)) OR mux_870_nl;
  mux_880_nl <= MUX_s_1_2_2(mux_879_nl, or_727_nl, fsm_output(5));
  vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_880_nl) AND (fsm_output(1));
  nor_1381_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (NOT and_763_cse));
  nor_1382_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR not_tmp_330);
  mux_892_nl <= MUX_s_1_2_2(nor_1381_nl, nor_1382_nl, fsm_output(0));
  nor_1383_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1384_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_891_nl <= MUX_s_1_2_2(nor_1383_nl, nor_1384_nl, fsm_output(0));
  mux_893_nl <= MUX_s_1_2_2(mux_892_nl, mux_891_nl, fsm_output(4));
  nor_1385_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1386_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_889_nl <= MUX_s_1_2_2(nor_1385_nl, nor_1386_nl, fsm_output(0));
  nor_1387_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1388_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_888_nl <= MUX_s_1_2_2(nor_1387_nl, nor_1388_nl, fsm_output(0));
  mux_890_nl <= MUX_s_1_2_2(mux_889_nl, mux_888_nl, fsm_output(4));
  mux_894_nl <= MUX_s_1_2_2(mux_893_nl, mux_890_nl, fsm_output(6));
  nand_466_nl <= NOT((fsm_output(2)) AND mux_894_nl);
  or_747_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (NOT and_763_cse);
  mux_885_nl <= MUX_s_1_2_2(or_tmp_633, or_747_nl, fsm_output(0));
  or_744_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_884_nl <= MUX_s_1_2_2(or_tmp_629, or_744_nl, fsm_output(0));
  mux_886_nl <= MUX_s_1_2_2(mux_885_nl, mux_884_nl, fsm_output(4));
  or_741_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_882_nl <= MUX_s_1_2_2(or_tmp_627, or_741_nl, fsm_output(0));
  or_738_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_881_nl <= MUX_s_1_2_2(or_tmp_623, or_738_nl, fsm_output(0));
  mux_883_nl <= MUX_s_1_2_2(mux_882_nl, mux_881_nl, fsm_output(4));
  mux_887_nl <= MUX_s_1_2_2(mux_886_nl, mux_883_nl, fsm_output(6));
  or_4139_nl <= (fsm_output(2)) OR mux_887_nl;
  mux_895_nl <= MUX_s_1_2_2(nand_466_nl, or_4139_nl, fsm_output(5));
  vec_rsc_0_3_i_we_d_pff <= NOT(mux_895_nl OR (fsm_output(1)));
  or_780_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_779_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_908_nl <= MUX_s_1_2_2(or_780_nl, or_779_nl, fsm_output(0));
  or_781_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_908_nl;
  or_777_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000011")) OR (NOT and_763_cse);
  mux_905_nl <= MUX_s_1_2_2(or_777_nl, or_tmp_633, fsm_output(0));
  or_775_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000011")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_904_nl <= MUX_s_1_2_2(or_775_nl, or_tmp_629, fsm_output(0));
  mux_906_nl <= MUX_s_1_2_2(mux_905_nl, mux_904_nl, fsm_output(4));
  or_774_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000011")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_902_nl <= MUX_s_1_2_2(or_774_nl, or_tmp_627, fsm_output(0));
  or_772_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000011")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_901_nl <= MUX_s_1_2_2(or_772_nl, or_tmp_623, fsm_output(0));
  mux_903_nl <= MUX_s_1_2_2(mux_902_nl, mux_901_nl, fsm_output(4));
  mux_907_nl <= MUX_s_1_2_2(mux_906_nl, mux_903_nl, fsm_output(6));
  mux_909_nl <= MUX_s_1_2_2(or_781_nl, mux_907_nl, fsm_output(2));
  or_770_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_768_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (NOT and_763_cse);
  mux_898_nl <= MUX_s_1_2_2(or_770_nl, or_768_nl, fsm_output(0));
  or_766_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_765_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_897_nl <= MUX_s_1_2_2(or_766_nl, or_765_nl, fsm_output(0));
  mux_899_nl <= MUX_s_1_2_2(mux_898_nl, mux_897_nl, fsm_output(4));
  nor_1379_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1380_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_896_nl <= MUX_s_1_2_2(nor_1379_nl, nor_1380_nl, fsm_output(0));
  nand_21_nl <= NOT((fsm_output(4)) AND mux_896_nl);
  mux_900_nl <= MUX_s_1_2_2(mux_899_nl, nand_21_nl, fsm_output(6));
  or_771_nl <= (fsm_output(2)) OR mux_900_nl;
  mux_910_nl <= MUX_s_1_2_2(mux_909_nl, or_771_nl, fsm_output(5));
  vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_910_nl) AND (fsm_output(1));
  nor_1370_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT and_763_cse));
  nor_1371_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_922_nl <= MUX_s_1_2_2(nor_1370_nl, nor_1371_nl, fsm_output(0));
  nor_1372_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1373_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_921_nl <= MUX_s_1_2_2(nor_1372_nl, nor_1373_nl, fsm_output(0));
  mux_923_nl <= MUX_s_1_2_2(mux_922_nl, mux_921_nl, fsm_output(4));
  nor_1374_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1375_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_919_nl <= MUX_s_1_2_2(nor_1374_nl, nor_1375_nl, fsm_output(0));
  nor_1376_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1377_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_918_nl <= MUX_s_1_2_2(nor_1376_nl, nor_1377_nl, fsm_output(0));
  mux_920_nl <= MUX_s_1_2_2(mux_919_nl, mux_918_nl, fsm_output(4));
  mux_924_nl <= MUX_s_1_2_2(mux_923_nl, mux_920_nl, fsm_output(6));
  nand_465_nl <= NOT((fsm_output(2)) AND mux_924_nl);
  or_791_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT and_763_cse);
  mux_915_nl <= MUX_s_1_2_2(or_tmp_677, or_791_nl, fsm_output(0));
  or_788_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_914_nl <= MUX_s_1_2_2(or_tmp_673, or_788_nl, fsm_output(0));
  mux_916_nl <= MUX_s_1_2_2(mux_915_nl, mux_914_nl, fsm_output(4));
  or_785_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_912_nl <= MUX_s_1_2_2(or_tmp_671, or_785_nl, fsm_output(0));
  or_782_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_911_nl <= MUX_s_1_2_2(or_tmp_667, or_782_nl, fsm_output(0));
  mux_913_nl <= MUX_s_1_2_2(mux_912_nl, mux_911_nl, fsm_output(4));
  mux_917_nl <= MUX_s_1_2_2(mux_916_nl, mux_913_nl, fsm_output(6));
  or_4138_nl <= (fsm_output(2)) OR mux_917_nl;
  mux_925_nl <= MUX_s_1_2_2(nand_465_nl, or_4138_nl, fsm_output(5));
  vec_rsc_0_4_i_we_d_pff <= NOT(mux_925_nl OR (fsm_output(1)));
  or_824_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_823_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_938_nl <= MUX_s_1_2_2(or_824_nl, or_823_nl, fsm_output(0));
  or_825_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_938_nl;
  or_821_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000100")) OR (NOT and_763_cse);
  mux_935_nl <= MUX_s_1_2_2(or_821_nl, or_tmp_677, fsm_output(0));
  or_819_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000100")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_934_nl <= MUX_s_1_2_2(or_819_nl, or_tmp_673, fsm_output(0));
  mux_936_nl <= MUX_s_1_2_2(mux_935_nl, mux_934_nl, fsm_output(4));
  or_818_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000100")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_932_nl <= MUX_s_1_2_2(or_818_nl, or_tmp_671, fsm_output(0));
  or_816_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000100")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_931_nl <= MUX_s_1_2_2(or_816_nl, or_tmp_667, fsm_output(0));
  mux_933_nl <= MUX_s_1_2_2(mux_932_nl, mux_931_nl, fsm_output(4));
  mux_937_nl <= MUX_s_1_2_2(mux_936_nl, mux_933_nl, fsm_output(6));
  mux_939_nl <= MUX_s_1_2_2(or_825_nl, mux_937_nl, fsm_output(2));
  or_814_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_812_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT and_763_cse);
  mux_928_nl <= MUX_s_1_2_2(or_814_nl, or_812_nl, fsm_output(0));
  or_810_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_809_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_927_nl <= MUX_s_1_2_2(or_810_nl, or_809_nl, fsm_output(0));
  mux_929_nl <= MUX_s_1_2_2(mux_928_nl, mux_927_nl, fsm_output(4));
  nor_1368_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1369_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_926_nl <= MUX_s_1_2_2(nor_1368_nl, nor_1369_nl, fsm_output(0));
  nand_23_nl <= NOT((fsm_output(4)) AND mux_926_nl);
  mux_930_nl <= MUX_s_1_2_2(mux_929_nl, nand_23_nl, fsm_output(6));
  or_815_nl <= (fsm_output(2)) OR mux_930_nl;
  mux_940_nl <= MUX_s_1_2_2(mux_939_nl, or_815_nl, fsm_output(5));
  vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_940_nl) AND (fsm_output(1));
  nor_1359_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (NOT and_763_cse));
  nor_1360_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_952_nl <= MUX_s_1_2_2(nor_1359_nl, nor_1360_nl, fsm_output(0));
  nor_1361_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1362_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_951_nl <= MUX_s_1_2_2(nor_1361_nl, nor_1362_nl, fsm_output(0));
  mux_953_nl <= MUX_s_1_2_2(mux_952_nl, mux_951_nl, fsm_output(4));
  nor_1363_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1364_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_949_nl <= MUX_s_1_2_2(nor_1363_nl, nor_1364_nl, fsm_output(0));
  nor_1365_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1366_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_948_nl <= MUX_s_1_2_2(nor_1365_nl, nor_1366_nl, fsm_output(0));
  mux_950_nl <= MUX_s_1_2_2(mux_949_nl, mux_948_nl, fsm_output(4));
  mux_954_nl <= MUX_s_1_2_2(mux_953_nl, mux_950_nl, fsm_output(6));
  nand_464_nl <= NOT((fsm_output(2)) AND mux_954_nl);
  or_835_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (NOT and_763_cse);
  mux_945_nl <= MUX_s_1_2_2(or_tmp_721, or_835_nl, fsm_output(0));
  or_832_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_944_nl <= MUX_s_1_2_2(or_tmp_717, or_832_nl, fsm_output(0));
  mux_946_nl <= MUX_s_1_2_2(mux_945_nl, mux_944_nl, fsm_output(4));
  or_829_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_942_nl <= MUX_s_1_2_2(or_tmp_715, or_829_nl, fsm_output(0));
  or_826_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_941_nl <= MUX_s_1_2_2(or_tmp_711, or_826_nl, fsm_output(0));
  mux_943_nl <= MUX_s_1_2_2(mux_942_nl, mux_941_nl, fsm_output(4));
  mux_947_nl <= MUX_s_1_2_2(mux_946_nl, mux_943_nl, fsm_output(6));
  or_4137_nl <= (fsm_output(2)) OR mux_947_nl;
  mux_955_nl <= MUX_s_1_2_2(nand_464_nl, or_4137_nl, fsm_output(5));
  vec_rsc_0_5_i_we_d_pff <= NOT(mux_955_nl OR (fsm_output(1)));
  or_868_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_867_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_968_nl <= MUX_s_1_2_2(or_868_nl, or_867_nl, fsm_output(0));
  or_869_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_968_nl;
  or_865_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000101")) OR (NOT and_763_cse);
  mux_965_nl <= MUX_s_1_2_2(or_865_nl, or_tmp_721, fsm_output(0));
  or_863_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000101")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_964_nl <= MUX_s_1_2_2(or_863_nl, or_tmp_717, fsm_output(0));
  mux_966_nl <= MUX_s_1_2_2(mux_965_nl, mux_964_nl, fsm_output(4));
  or_862_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000101")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_962_nl <= MUX_s_1_2_2(or_862_nl, or_tmp_715, fsm_output(0));
  or_860_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000101")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_961_nl <= MUX_s_1_2_2(or_860_nl, or_tmp_711, fsm_output(0));
  mux_963_nl <= MUX_s_1_2_2(mux_962_nl, mux_961_nl, fsm_output(4));
  mux_967_nl <= MUX_s_1_2_2(mux_966_nl, mux_963_nl, fsm_output(6));
  mux_969_nl <= MUX_s_1_2_2(or_869_nl, mux_967_nl, fsm_output(2));
  or_858_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_856_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (NOT and_763_cse);
  mux_958_nl <= MUX_s_1_2_2(or_858_nl, or_856_nl, fsm_output(0));
  or_854_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_853_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_957_nl <= MUX_s_1_2_2(or_854_nl, or_853_nl, fsm_output(0));
  mux_959_nl <= MUX_s_1_2_2(mux_958_nl, mux_957_nl, fsm_output(4));
  nor_1357_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1358_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_956_nl <= MUX_s_1_2_2(nor_1357_nl, nor_1358_nl, fsm_output(0));
  nand_25_nl <= NOT((fsm_output(4)) AND mux_956_nl);
  mux_960_nl <= MUX_s_1_2_2(mux_959_nl, nand_25_nl, fsm_output(6));
  or_859_nl <= (fsm_output(2)) OR mux_960_nl;
  mux_970_nl <= MUX_s_1_2_2(mux_969_nl, or_859_nl, fsm_output(5));
  vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_970_nl) AND (fsm_output(1));
  nor_1348_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT and_763_cse));
  nor_1349_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_982_nl <= MUX_s_1_2_2(nor_1348_nl, nor_1349_nl, fsm_output(0));
  nor_1350_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1351_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_981_nl <= MUX_s_1_2_2(nor_1350_nl, nor_1351_nl, fsm_output(0));
  mux_983_nl <= MUX_s_1_2_2(mux_982_nl, mux_981_nl, fsm_output(4));
  nor_1352_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1353_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_979_nl <= MUX_s_1_2_2(nor_1352_nl, nor_1353_nl, fsm_output(0));
  nor_1354_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1355_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_978_nl <= MUX_s_1_2_2(nor_1354_nl, nor_1355_nl, fsm_output(0));
  mux_980_nl <= MUX_s_1_2_2(mux_979_nl, mux_978_nl, fsm_output(4));
  mux_984_nl <= MUX_s_1_2_2(mux_983_nl, mux_980_nl, fsm_output(6));
  nand_463_nl <= NOT((fsm_output(2)) AND mux_984_nl);
  or_879_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT and_763_cse);
  mux_975_nl <= MUX_s_1_2_2(or_tmp_765, or_879_nl, fsm_output(0));
  or_876_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_974_nl <= MUX_s_1_2_2(or_tmp_761, or_876_nl, fsm_output(0));
  mux_976_nl <= MUX_s_1_2_2(mux_975_nl, mux_974_nl, fsm_output(4));
  or_873_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_972_nl <= MUX_s_1_2_2(or_tmp_759, or_873_nl, fsm_output(0));
  or_870_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_971_nl <= MUX_s_1_2_2(or_tmp_755, or_870_nl, fsm_output(0));
  mux_973_nl <= MUX_s_1_2_2(mux_972_nl, mux_971_nl, fsm_output(4));
  mux_977_nl <= MUX_s_1_2_2(mux_976_nl, mux_973_nl, fsm_output(6));
  or_4136_nl <= (fsm_output(2)) OR mux_977_nl;
  mux_985_nl <= MUX_s_1_2_2(nand_463_nl, or_4136_nl, fsm_output(5));
  vec_rsc_0_6_i_we_d_pff <= NOT(mux_985_nl OR (fsm_output(1)));
  or_912_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_911_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_998_nl <= MUX_s_1_2_2(or_912_nl, or_911_nl, fsm_output(0));
  or_913_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_998_nl;
  or_909_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000110")) OR (NOT and_763_cse);
  mux_995_nl <= MUX_s_1_2_2(or_909_nl, or_tmp_765, fsm_output(0));
  or_907_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000110")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_994_nl <= MUX_s_1_2_2(or_907_nl, or_tmp_761, fsm_output(0));
  mux_996_nl <= MUX_s_1_2_2(mux_995_nl, mux_994_nl, fsm_output(4));
  or_906_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000110")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_992_nl <= MUX_s_1_2_2(or_906_nl, or_tmp_759, fsm_output(0));
  or_904_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000110")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_991_nl <= MUX_s_1_2_2(or_904_nl, or_tmp_755, fsm_output(0));
  mux_993_nl <= MUX_s_1_2_2(mux_992_nl, mux_991_nl, fsm_output(4));
  mux_997_nl <= MUX_s_1_2_2(mux_996_nl, mux_993_nl, fsm_output(6));
  mux_999_nl <= MUX_s_1_2_2(or_913_nl, mux_997_nl, fsm_output(2));
  or_902_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_900_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT and_763_cse);
  mux_988_nl <= MUX_s_1_2_2(or_902_nl, or_900_nl, fsm_output(0));
  or_898_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_897_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_987_nl <= MUX_s_1_2_2(or_898_nl, or_897_nl, fsm_output(0));
  mux_989_nl <= MUX_s_1_2_2(mux_988_nl, mux_987_nl, fsm_output(4));
  nor_1346_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1347_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_986_nl <= MUX_s_1_2_2(nor_1346_nl, nor_1347_nl, fsm_output(0));
  nand_27_nl <= NOT((fsm_output(4)) AND mux_986_nl);
  mux_990_nl <= MUX_s_1_2_2(mux_989_nl, nand_27_nl, fsm_output(6));
  or_903_nl <= (fsm_output(2)) OR mux_990_nl;
  mux_1000_nl <= MUX_s_1_2_2(mux_999_nl, or_903_nl, fsm_output(5));
  vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1000_nl) AND (fsm_output(1));
  nor_1337_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (NOT and_763_cse));
  nor_1338_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))
      OR not_tmp_347);
  mux_1012_nl <= MUX_s_1_2_2(nor_1337_nl, nor_1338_nl, fsm_output(0));
  nor_1339_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1340_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1011_nl <= MUX_s_1_2_2(nor_1339_nl, nor_1340_nl, fsm_output(0));
  mux_1013_nl <= MUX_s_1_2_2(mux_1012_nl, mux_1011_nl, fsm_output(4));
  nor_1341_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1342_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1009_nl <= MUX_s_1_2_2(nor_1341_nl, nor_1342_nl, fsm_output(0));
  nor_1343_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1344_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1008_nl <= MUX_s_1_2_2(nor_1343_nl, nor_1344_nl, fsm_output(0));
  mux_1010_nl <= MUX_s_1_2_2(mux_1009_nl, mux_1008_nl, fsm_output(4));
  mux_1014_nl <= MUX_s_1_2_2(mux_1013_nl, mux_1010_nl, fsm_output(6));
  nand_462_nl <= NOT((fsm_output(2)) AND mux_1014_nl);
  or_923_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (NOT and_763_cse);
  mux_1005_nl <= MUX_s_1_2_2(or_tmp_809, or_923_nl, fsm_output(0));
  or_920_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1004_nl <= MUX_s_1_2_2(or_tmp_805, or_920_nl, fsm_output(0));
  mux_1006_nl <= MUX_s_1_2_2(mux_1005_nl, mux_1004_nl, fsm_output(4));
  or_917_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1002_nl <= MUX_s_1_2_2(or_tmp_803, or_917_nl, fsm_output(0));
  or_914_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1001_nl <= MUX_s_1_2_2(or_tmp_799, or_914_nl, fsm_output(0));
  mux_1003_nl <= MUX_s_1_2_2(mux_1002_nl, mux_1001_nl, fsm_output(4));
  mux_1007_nl <= MUX_s_1_2_2(mux_1006_nl, mux_1003_nl, fsm_output(6));
  or_4135_nl <= (fsm_output(2)) OR mux_1007_nl;
  mux_1015_nl <= MUX_s_1_2_2(nand_462_nl, or_4135_nl, fsm_output(5));
  vec_rsc_0_7_i_we_d_pff <= NOT(mux_1015_nl OR (fsm_output(1)));
  or_956_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_955_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1028_nl <= MUX_s_1_2_2(or_956_nl, or_955_nl, fsm_output(0));
  or_957_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1028_nl;
  or_953_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000111")) OR (NOT and_763_cse);
  mux_1025_nl <= MUX_s_1_2_2(or_953_nl, or_tmp_809, fsm_output(0));
  or_951_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000111")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1024_nl <= MUX_s_1_2_2(or_951_nl, or_tmp_805, fsm_output(0));
  mux_1026_nl <= MUX_s_1_2_2(mux_1025_nl, mux_1024_nl, fsm_output(4));
  or_950_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000111")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1022_nl <= MUX_s_1_2_2(or_950_nl, or_tmp_803, fsm_output(0));
  or_948_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000111")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1021_nl <= MUX_s_1_2_2(or_948_nl, or_tmp_799, fsm_output(0));
  mux_1023_nl <= MUX_s_1_2_2(mux_1022_nl, mux_1021_nl, fsm_output(4));
  mux_1027_nl <= MUX_s_1_2_2(mux_1026_nl, mux_1023_nl, fsm_output(6));
  mux_1029_nl <= MUX_s_1_2_2(or_957_nl, mux_1027_nl, fsm_output(2));
  or_946_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_944_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (NOT and_763_cse);
  mux_1018_nl <= MUX_s_1_2_2(or_946_nl, or_944_nl, fsm_output(0));
  or_942_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_941_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1017_nl <= MUX_s_1_2_2(or_942_nl, or_941_nl, fsm_output(0));
  mux_1019_nl <= MUX_s_1_2_2(mux_1018_nl, mux_1017_nl, fsm_output(4));
  nor_1335_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1336_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1016_nl <= MUX_s_1_2_2(nor_1335_nl, nor_1336_nl, fsm_output(0));
  nand_29_nl <= NOT((fsm_output(4)) AND mux_1016_nl);
  mux_1020_nl <= MUX_s_1_2_2(mux_1019_nl, nand_29_nl, fsm_output(6));
  or_947_nl <= (fsm_output(2)) OR mux_1020_nl;
  mux_1030_nl <= MUX_s_1_2_2(mux_1029_nl, or_947_nl, fsm_output(5));
  vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1030_nl) AND (fsm_output(1));
  nor_1326_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT and_763_cse));
  nor_1327_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_1042_nl <= MUX_s_1_2_2(nor_1326_nl, nor_1327_nl, fsm_output(0));
  nor_1328_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1329_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1041_nl <= MUX_s_1_2_2(nor_1328_nl, nor_1329_nl, fsm_output(0));
  mux_1043_nl <= MUX_s_1_2_2(mux_1042_nl, mux_1041_nl, fsm_output(4));
  nor_1330_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1331_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1039_nl <= MUX_s_1_2_2(nor_1330_nl, nor_1331_nl, fsm_output(0));
  nor_1332_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1333_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1038_nl <= MUX_s_1_2_2(nor_1332_nl, nor_1333_nl, fsm_output(0));
  mux_1040_nl <= MUX_s_1_2_2(mux_1039_nl, mux_1038_nl, fsm_output(4));
  mux_1044_nl <= MUX_s_1_2_2(mux_1043_nl, mux_1040_nl, fsm_output(6));
  nand_461_nl <= NOT((fsm_output(2)) AND mux_1044_nl);
  or_967_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT and_763_cse);
  mux_1035_nl <= MUX_s_1_2_2(or_tmp_853, or_967_nl, fsm_output(0));
  or_964_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1034_nl <= MUX_s_1_2_2(or_tmp_849, or_964_nl, fsm_output(0));
  mux_1036_nl <= MUX_s_1_2_2(mux_1035_nl, mux_1034_nl, fsm_output(4));
  or_961_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1032_nl <= MUX_s_1_2_2(or_tmp_847, or_961_nl, fsm_output(0));
  or_958_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1031_nl <= MUX_s_1_2_2(or_tmp_843, or_958_nl, fsm_output(0));
  mux_1033_nl <= MUX_s_1_2_2(mux_1032_nl, mux_1031_nl, fsm_output(4));
  mux_1037_nl <= MUX_s_1_2_2(mux_1036_nl, mux_1033_nl, fsm_output(6));
  or_4134_nl <= (fsm_output(2)) OR mux_1037_nl;
  mux_1045_nl <= MUX_s_1_2_2(nand_461_nl, or_4134_nl, fsm_output(5));
  vec_rsc_0_8_i_we_d_pff <= NOT(mux_1045_nl OR (fsm_output(1)));
  or_1000_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_999_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1058_nl <= MUX_s_1_2_2(or_1000_nl, or_999_nl, fsm_output(0));
  or_1001_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1058_nl;
  or_997_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001000")) OR (NOT and_763_cse);
  mux_1055_nl <= MUX_s_1_2_2(or_997_nl, or_tmp_853, fsm_output(0));
  or_995_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001000")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1054_nl <= MUX_s_1_2_2(or_995_nl, or_tmp_849, fsm_output(0));
  mux_1056_nl <= MUX_s_1_2_2(mux_1055_nl, mux_1054_nl, fsm_output(4));
  or_994_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001000")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1052_nl <= MUX_s_1_2_2(or_994_nl, or_tmp_847, fsm_output(0));
  or_992_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001000")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1051_nl <= MUX_s_1_2_2(or_992_nl, or_tmp_843, fsm_output(0));
  mux_1053_nl <= MUX_s_1_2_2(mux_1052_nl, mux_1051_nl, fsm_output(4));
  mux_1057_nl <= MUX_s_1_2_2(mux_1056_nl, mux_1053_nl, fsm_output(6));
  mux_1059_nl <= MUX_s_1_2_2(or_1001_nl, mux_1057_nl, fsm_output(2));
  or_990_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_988_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT and_763_cse);
  mux_1048_nl <= MUX_s_1_2_2(or_990_nl, or_988_nl, fsm_output(0));
  or_986_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_985_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1047_nl <= MUX_s_1_2_2(or_986_nl, or_985_nl, fsm_output(0));
  mux_1049_nl <= MUX_s_1_2_2(mux_1048_nl, mux_1047_nl, fsm_output(4));
  nor_1324_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1325_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1046_nl <= MUX_s_1_2_2(nor_1324_nl, nor_1325_nl, fsm_output(0));
  nand_31_nl <= NOT((fsm_output(4)) AND mux_1046_nl);
  mux_1050_nl <= MUX_s_1_2_2(mux_1049_nl, nand_31_nl, fsm_output(6));
  or_991_nl <= (fsm_output(2)) OR mux_1050_nl;
  mux_1060_nl <= MUX_s_1_2_2(mux_1059_nl, or_991_nl, fsm_output(5));
  vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1060_nl) AND (fsm_output(1));
  nor_1315_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (NOT and_763_cse));
  nor_1316_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_1072_nl <= MUX_s_1_2_2(nor_1315_nl, nor_1316_nl, fsm_output(0));
  nor_1317_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1318_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1071_nl <= MUX_s_1_2_2(nor_1317_nl, nor_1318_nl, fsm_output(0));
  mux_1073_nl <= MUX_s_1_2_2(mux_1072_nl, mux_1071_nl, fsm_output(4));
  nor_1319_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1320_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1069_nl <= MUX_s_1_2_2(nor_1319_nl, nor_1320_nl, fsm_output(0));
  nor_1321_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1322_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1068_nl <= MUX_s_1_2_2(nor_1321_nl, nor_1322_nl, fsm_output(0));
  mux_1070_nl <= MUX_s_1_2_2(mux_1069_nl, mux_1068_nl, fsm_output(4));
  mux_1074_nl <= MUX_s_1_2_2(mux_1073_nl, mux_1070_nl, fsm_output(6));
  nand_460_nl <= NOT((fsm_output(2)) AND mux_1074_nl);
  or_1011_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (NOT and_763_cse);
  mux_1065_nl <= MUX_s_1_2_2(or_tmp_897, or_1011_nl, fsm_output(0));
  or_1008_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1064_nl <= MUX_s_1_2_2(or_tmp_893, or_1008_nl, fsm_output(0));
  mux_1066_nl <= MUX_s_1_2_2(mux_1065_nl, mux_1064_nl, fsm_output(4));
  or_1005_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1062_nl <= MUX_s_1_2_2(or_tmp_891, or_1005_nl, fsm_output(0));
  or_1002_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1061_nl <= MUX_s_1_2_2(or_tmp_887, or_1002_nl, fsm_output(0));
  mux_1063_nl <= MUX_s_1_2_2(mux_1062_nl, mux_1061_nl, fsm_output(4));
  mux_1067_nl <= MUX_s_1_2_2(mux_1066_nl, mux_1063_nl, fsm_output(6));
  or_4133_nl <= (fsm_output(2)) OR mux_1067_nl;
  mux_1075_nl <= MUX_s_1_2_2(nand_460_nl, or_4133_nl, fsm_output(5));
  vec_rsc_0_9_i_we_d_pff <= NOT(mux_1075_nl OR (fsm_output(1)));
  or_1044_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1043_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1088_nl <= MUX_s_1_2_2(or_1044_nl, or_1043_nl, fsm_output(0));
  or_1045_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1088_nl;
  or_1041_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001001")) OR (NOT and_763_cse);
  mux_1085_nl <= MUX_s_1_2_2(or_1041_nl, or_tmp_897, fsm_output(0));
  or_1039_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001001")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1084_nl <= MUX_s_1_2_2(or_1039_nl, or_tmp_893, fsm_output(0));
  mux_1086_nl <= MUX_s_1_2_2(mux_1085_nl, mux_1084_nl, fsm_output(4));
  or_1038_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001001")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1082_nl <= MUX_s_1_2_2(or_1038_nl, or_tmp_891, fsm_output(0));
  or_1036_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001001")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1081_nl <= MUX_s_1_2_2(or_1036_nl, or_tmp_887, fsm_output(0));
  mux_1083_nl <= MUX_s_1_2_2(mux_1082_nl, mux_1081_nl, fsm_output(4));
  mux_1087_nl <= MUX_s_1_2_2(mux_1086_nl, mux_1083_nl, fsm_output(6));
  mux_1089_nl <= MUX_s_1_2_2(or_1045_nl, mux_1087_nl, fsm_output(2));
  or_1034_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1032_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (NOT and_763_cse);
  mux_1078_nl <= MUX_s_1_2_2(or_1034_nl, or_1032_nl, fsm_output(0));
  or_1030_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1029_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1077_nl <= MUX_s_1_2_2(or_1030_nl, or_1029_nl, fsm_output(0));
  mux_1079_nl <= MUX_s_1_2_2(mux_1078_nl, mux_1077_nl, fsm_output(4));
  nor_1313_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1314_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1076_nl <= MUX_s_1_2_2(nor_1313_nl, nor_1314_nl, fsm_output(0));
  nand_33_nl <= NOT((fsm_output(4)) AND mux_1076_nl);
  mux_1080_nl <= MUX_s_1_2_2(mux_1079_nl, nand_33_nl, fsm_output(6));
  or_1035_nl <= (fsm_output(2)) OR mux_1080_nl;
  mux_1090_nl <= MUX_s_1_2_2(mux_1089_nl, or_1035_nl, fsm_output(5));
  vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1090_nl) AND (fsm_output(1));
  nor_1304_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT and_763_cse));
  nor_1305_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_1102_nl <= MUX_s_1_2_2(nor_1304_nl, nor_1305_nl, fsm_output(0));
  nor_1306_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1307_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1101_nl <= MUX_s_1_2_2(nor_1306_nl, nor_1307_nl, fsm_output(0));
  mux_1103_nl <= MUX_s_1_2_2(mux_1102_nl, mux_1101_nl, fsm_output(4));
  nor_1308_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1309_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1099_nl <= MUX_s_1_2_2(nor_1308_nl, nor_1309_nl, fsm_output(0));
  nor_1310_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1311_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1098_nl <= MUX_s_1_2_2(nor_1310_nl, nor_1311_nl, fsm_output(0));
  mux_1100_nl <= MUX_s_1_2_2(mux_1099_nl, mux_1098_nl, fsm_output(4));
  mux_1104_nl <= MUX_s_1_2_2(mux_1103_nl, mux_1100_nl, fsm_output(6));
  nand_459_nl <= NOT((fsm_output(2)) AND mux_1104_nl);
  or_1055_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT and_763_cse);
  mux_1095_nl <= MUX_s_1_2_2(or_tmp_941, or_1055_nl, fsm_output(0));
  or_1052_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1094_nl <= MUX_s_1_2_2(or_tmp_937, or_1052_nl, fsm_output(0));
  mux_1096_nl <= MUX_s_1_2_2(mux_1095_nl, mux_1094_nl, fsm_output(4));
  or_1049_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1092_nl <= MUX_s_1_2_2(or_tmp_935, or_1049_nl, fsm_output(0));
  or_1046_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1091_nl <= MUX_s_1_2_2(or_tmp_931, or_1046_nl, fsm_output(0));
  mux_1093_nl <= MUX_s_1_2_2(mux_1092_nl, mux_1091_nl, fsm_output(4));
  mux_1097_nl <= MUX_s_1_2_2(mux_1096_nl, mux_1093_nl, fsm_output(6));
  or_4132_nl <= (fsm_output(2)) OR mux_1097_nl;
  mux_1105_nl <= MUX_s_1_2_2(nand_459_nl, or_4132_nl, fsm_output(5));
  vec_rsc_0_10_i_we_d_pff <= NOT(mux_1105_nl OR (fsm_output(1)));
  or_1088_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1087_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1118_nl <= MUX_s_1_2_2(or_1088_nl, or_1087_nl, fsm_output(0));
  or_1089_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1118_nl;
  or_1085_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001010")) OR (NOT and_763_cse);
  mux_1115_nl <= MUX_s_1_2_2(or_1085_nl, or_tmp_941, fsm_output(0));
  or_1083_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001010")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1114_nl <= MUX_s_1_2_2(or_1083_nl, or_tmp_937, fsm_output(0));
  mux_1116_nl <= MUX_s_1_2_2(mux_1115_nl, mux_1114_nl, fsm_output(4));
  or_1082_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001010")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1112_nl <= MUX_s_1_2_2(or_1082_nl, or_tmp_935, fsm_output(0));
  or_1080_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001010")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1111_nl <= MUX_s_1_2_2(or_1080_nl, or_tmp_931, fsm_output(0));
  mux_1113_nl <= MUX_s_1_2_2(mux_1112_nl, mux_1111_nl, fsm_output(4));
  mux_1117_nl <= MUX_s_1_2_2(mux_1116_nl, mux_1113_nl, fsm_output(6));
  mux_1119_nl <= MUX_s_1_2_2(or_1089_nl, mux_1117_nl, fsm_output(2));
  or_1078_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1076_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT and_763_cse);
  mux_1108_nl <= MUX_s_1_2_2(or_1078_nl, or_1076_nl, fsm_output(0));
  or_1074_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1073_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1107_nl <= MUX_s_1_2_2(or_1074_nl, or_1073_nl, fsm_output(0));
  mux_1109_nl <= MUX_s_1_2_2(mux_1108_nl, mux_1107_nl, fsm_output(4));
  nor_1302_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1303_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1106_nl <= MUX_s_1_2_2(nor_1302_nl, nor_1303_nl, fsm_output(0));
  nand_35_nl <= NOT((fsm_output(4)) AND mux_1106_nl);
  mux_1110_nl <= MUX_s_1_2_2(mux_1109_nl, nand_35_nl, fsm_output(6));
  or_1079_nl <= (fsm_output(2)) OR mux_1110_nl;
  mux_1120_nl <= MUX_s_1_2_2(mux_1119_nl, or_1079_nl, fsm_output(5));
  vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1120_nl) AND (fsm_output(1));
  nor_1293_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (NOT and_763_cse));
  nor_1294_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR not_tmp_330);
  mux_1132_nl <= MUX_s_1_2_2(nor_1293_nl, nor_1294_nl, fsm_output(0));
  nor_1295_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1296_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1131_nl <= MUX_s_1_2_2(nor_1295_nl, nor_1296_nl, fsm_output(0));
  mux_1133_nl <= MUX_s_1_2_2(mux_1132_nl, mux_1131_nl, fsm_output(4));
  nor_1297_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1298_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1129_nl <= MUX_s_1_2_2(nor_1297_nl, nor_1298_nl, fsm_output(0));
  nor_1299_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1300_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1128_nl <= MUX_s_1_2_2(nor_1299_nl, nor_1300_nl, fsm_output(0));
  mux_1130_nl <= MUX_s_1_2_2(mux_1129_nl, mux_1128_nl, fsm_output(4));
  mux_1134_nl <= MUX_s_1_2_2(mux_1133_nl, mux_1130_nl, fsm_output(6));
  nand_458_nl <= NOT((fsm_output(2)) AND mux_1134_nl);
  or_1099_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (NOT and_763_cse);
  mux_1125_nl <= MUX_s_1_2_2(or_tmp_985, or_1099_nl, fsm_output(0));
  or_1096_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1124_nl <= MUX_s_1_2_2(or_tmp_981, or_1096_nl, fsm_output(0));
  mux_1126_nl <= MUX_s_1_2_2(mux_1125_nl, mux_1124_nl, fsm_output(4));
  or_1093_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1122_nl <= MUX_s_1_2_2(or_tmp_979, or_1093_nl, fsm_output(0));
  or_1090_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1121_nl <= MUX_s_1_2_2(or_tmp_975, or_1090_nl, fsm_output(0));
  mux_1123_nl <= MUX_s_1_2_2(mux_1122_nl, mux_1121_nl, fsm_output(4));
  mux_1127_nl <= MUX_s_1_2_2(mux_1126_nl, mux_1123_nl, fsm_output(6));
  or_4131_nl <= (fsm_output(2)) OR mux_1127_nl;
  mux_1135_nl <= MUX_s_1_2_2(nand_458_nl, or_4131_nl, fsm_output(5));
  vec_rsc_0_11_i_we_d_pff <= NOT(mux_1135_nl OR (fsm_output(1)));
  or_1132_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1131_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1148_nl <= MUX_s_1_2_2(or_1132_nl, or_1131_nl, fsm_output(0));
  or_1133_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1148_nl;
  or_1129_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001011")) OR (NOT and_763_cse);
  mux_1145_nl <= MUX_s_1_2_2(or_1129_nl, or_tmp_985, fsm_output(0));
  or_1127_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001011")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1144_nl <= MUX_s_1_2_2(or_1127_nl, or_tmp_981, fsm_output(0));
  mux_1146_nl <= MUX_s_1_2_2(mux_1145_nl, mux_1144_nl, fsm_output(4));
  or_1126_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001011")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1142_nl <= MUX_s_1_2_2(or_1126_nl, or_tmp_979, fsm_output(0));
  or_1124_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001011")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1141_nl <= MUX_s_1_2_2(or_1124_nl, or_tmp_975, fsm_output(0));
  mux_1143_nl <= MUX_s_1_2_2(mux_1142_nl, mux_1141_nl, fsm_output(4));
  mux_1147_nl <= MUX_s_1_2_2(mux_1146_nl, mux_1143_nl, fsm_output(6));
  mux_1149_nl <= MUX_s_1_2_2(or_1133_nl, mux_1147_nl, fsm_output(2));
  or_1122_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1120_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (NOT and_763_cse);
  mux_1138_nl <= MUX_s_1_2_2(or_1122_nl, or_1120_nl, fsm_output(0));
  or_1118_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1117_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1137_nl <= MUX_s_1_2_2(or_1118_nl, or_1117_nl, fsm_output(0));
  mux_1139_nl <= MUX_s_1_2_2(mux_1138_nl, mux_1137_nl, fsm_output(4));
  nor_1291_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1292_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1136_nl <= MUX_s_1_2_2(nor_1291_nl, nor_1292_nl, fsm_output(0));
  nand_37_nl <= NOT((fsm_output(4)) AND mux_1136_nl);
  mux_1140_nl <= MUX_s_1_2_2(mux_1139_nl, nand_37_nl, fsm_output(6));
  or_1123_nl <= (fsm_output(2)) OR mux_1140_nl;
  mux_1150_nl <= MUX_s_1_2_2(mux_1149_nl, or_1123_nl, fsm_output(5));
  vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1150_nl) AND (fsm_output(1));
  nor_1282_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT and_763_cse));
  nor_1283_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_1162_nl <= MUX_s_1_2_2(nor_1282_nl, nor_1283_nl, fsm_output(0));
  nor_1284_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1285_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1161_nl <= MUX_s_1_2_2(nor_1284_nl, nor_1285_nl, fsm_output(0));
  mux_1163_nl <= MUX_s_1_2_2(mux_1162_nl, mux_1161_nl, fsm_output(4));
  nor_1286_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1287_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1159_nl <= MUX_s_1_2_2(nor_1286_nl, nor_1287_nl, fsm_output(0));
  nor_1288_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1289_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1158_nl <= MUX_s_1_2_2(nor_1288_nl, nor_1289_nl, fsm_output(0));
  mux_1160_nl <= MUX_s_1_2_2(mux_1159_nl, mux_1158_nl, fsm_output(4));
  mux_1164_nl <= MUX_s_1_2_2(mux_1163_nl, mux_1160_nl, fsm_output(6));
  nand_457_nl <= NOT((fsm_output(2)) AND mux_1164_nl);
  or_1143_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT and_763_cse);
  mux_1155_nl <= MUX_s_1_2_2(or_tmp_1029, or_1143_nl, fsm_output(0));
  or_1140_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1154_nl <= MUX_s_1_2_2(or_tmp_1025, or_1140_nl, fsm_output(0));
  mux_1156_nl <= MUX_s_1_2_2(mux_1155_nl, mux_1154_nl, fsm_output(4));
  or_1137_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1152_nl <= MUX_s_1_2_2(or_tmp_1023, or_1137_nl, fsm_output(0));
  or_1134_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1151_nl <= MUX_s_1_2_2(or_tmp_1019, or_1134_nl, fsm_output(0));
  mux_1153_nl <= MUX_s_1_2_2(mux_1152_nl, mux_1151_nl, fsm_output(4));
  mux_1157_nl <= MUX_s_1_2_2(mux_1156_nl, mux_1153_nl, fsm_output(6));
  or_4130_nl <= (fsm_output(2)) OR mux_1157_nl;
  mux_1165_nl <= MUX_s_1_2_2(nand_457_nl, or_4130_nl, fsm_output(5));
  vec_rsc_0_12_i_we_d_pff <= NOT(mux_1165_nl OR (fsm_output(1)));
  or_1176_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1175_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1178_nl <= MUX_s_1_2_2(or_1176_nl, or_1175_nl, fsm_output(0));
  or_1177_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1178_nl;
  or_1173_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001100")) OR (NOT and_763_cse);
  mux_1175_nl <= MUX_s_1_2_2(or_1173_nl, or_tmp_1029, fsm_output(0));
  or_1171_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001100")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1174_nl <= MUX_s_1_2_2(or_1171_nl, or_tmp_1025, fsm_output(0));
  mux_1176_nl <= MUX_s_1_2_2(mux_1175_nl, mux_1174_nl, fsm_output(4));
  or_1170_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001100")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1172_nl <= MUX_s_1_2_2(or_1170_nl, or_tmp_1023, fsm_output(0));
  or_1168_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001100")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1171_nl <= MUX_s_1_2_2(or_1168_nl, or_tmp_1019, fsm_output(0));
  mux_1173_nl <= MUX_s_1_2_2(mux_1172_nl, mux_1171_nl, fsm_output(4));
  mux_1177_nl <= MUX_s_1_2_2(mux_1176_nl, mux_1173_nl, fsm_output(6));
  mux_1179_nl <= MUX_s_1_2_2(or_1177_nl, mux_1177_nl, fsm_output(2));
  or_1166_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1164_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT and_763_cse);
  mux_1168_nl <= MUX_s_1_2_2(or_1166_nl, or_1164_nl, fsm_output(0));
  or_1162_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1161_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1167_nl <= MUX_s_1_2_2(or_1162_nl, or_1161_nl, fsm_output(0));
  mux_1169_nl <= MUX_s_1_2_2(mux_1168_nl, mux_1167_nl, fsm_output(4));
  nor_1280_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1281_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1166_nl <= MUX_s_1_2_2(nor_1280_nl, nor_1281_nl, fsm_output(0));
  nand_39_nl <= NOT((fsm_output(4)) AND mux_1166_nl);
  mux_1170_nl <= MUX_s_1_2_2(mux_1169_nl, nand_39_nl, fsm_output(6));
  or_1167_nl <= (fsm_output(2)) OR mux_1170_nl;
  mux_1180_nl <= MUX_s_1_2_2(mux_1179_nl, or_1167_nl, fsm_output(5));
  vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1180_nl) AND (fsm_output(1));
  nor_1271_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (NOT and_763_cse));
  nor_1272_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_1192_nl <= MUX_s_1_2_2(nor_1271_nl, nor_1272_nl, fsm_output(0));
  nor_1273_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1274_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1191_nl <= MUX_s_1_2_2(nor_1273_nl, nor_1274_nl, fsm_output(0));
  mux_1193_nl <= MUX_s_1_2_2(mux_1192_nl, mux_1191_nl, fsm_output(4));
  nor_1275_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1276_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1189_nl <= MUX_s_1_2_2(nor_1275_nl, nor_1276_nl, fsm_output(0));
  nor_1277_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1278_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1188_nl <= MUX_s_1_2_2(nor_1277_nl, nor_1278_nl, fsm_output(0));
  mux_1190_nl <= MUX_s_1_2_2(mux_1189_nl, mux_1188_nl, fsm_output(4));
  mux_1194_nl <= MUX_s_1_2_2(mux_1193_nl, mux_1190_nl, fsm_output(6));
  nand_456_nl <= NOT((fsm_output(2)) AND mux_1194_nl);
  or_1187_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (NOT and_763_cse);
  mux_1185_nl <= MUX_s_1_2_2(or_tmp_1073, or_1187_nl, fsm_output(0));
  or_1184_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1184_nl <= MUX_s_1_2_2(or_tmp_1069, or_1184_nl, fsm_output(0));
  mux_1186_nl <= MUX_s_1_2_2(mux_1185_nl, mux_1184_nl, fsm_output(4));
  or_1181_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1182_nl <= MUX_s_1_2_2(or_tmp_1067, or_1181_nl, fsm_output(0));
  or_1178_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1181_nl <= MUX_s_1_2_2(or_tmp_1063, or_1178_nl, fsm_output(0));
  mux_1183_nl <= MUX_s_1_2_2(mux_1182_nl, mux_1181_nl, fsm_output(4));
  mux_1187_nl <= MUX_s_1_2_2(mux_1186_nl, mux_1183_nl, fsm_output(6));
  or_4129_nl <= (fsm_output(2)) OR mux_1187_nl;
  mux_1195_nl <= MUX_s_1_2_2(nand_456_nl, or_4129_nl, fsm_output(5));
  vec_rsc_0_13_i_we_d_pff <= NOT(mux_1195_nl OR (fsm_output(1)));
  or_1220_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1219_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1208_nl <= MUX_s_1_2_2(or_1220_nl, or_1219_nl, fsm_output(0));
  or_1221_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1208_nl;
  or_1217_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001101")) OR (NOT and_763_cse);
  mux_1205_nl <= MUX_s_1_2_2(or_1217_nl, or_tmp_1073, fsm_output(0));
  or_1215_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001101")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1204_nl <= MUX_s_1_2_2(or_1215_nl, or_tmp_1069, fsm_output(0));
  mux_1206_nl <= MUX_s_1_2_2(mux_1205_nl, mux_1204_nl, fsm_output(4));
  or_1214_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001101")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1202_nl <= MUX_s_1_2_2(or_1214_nl, or_tmp_1067, fsm_output(0));
  or_1212_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001101")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1201_nl <= MUX_s_1_2_2(or_1212_nl, or_tmp_1063, fsm_output(0));
  mux_1203_nl <= MUX_s_1_2_2(mux_1202_nl, mux_1201_nl, fsm_output(4));
  mux_1207_nl <= MUX_s_1_2_2(mux_1206_nl, mux_1203_nl, fsm_output(6));
  mux_1209_nl <= MUX_s_1_2_2(or_1221_nl, mux_1207_nl, fsm_output(2));
  or_1210_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1208_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (NOT and_763_cse);
  mux_1198_nl <= MUX_s_1_2_2(or_1210_nl, or_1208_nl, fsm_output(0));
  or_1206_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1205_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1197_nl <= MUX_s_1_2_2(or_1206_nl, or_1205_nl, fsm_output(0));
  mux_1199_nl <= MUX_s_1_2_2(mux_1198_nl, mux_1197_nl, fsm_output(4));
  nor_1269_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1270_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1196_nl <= MUX_s_1_2_2(nor_1269_nl, nor_1270_nl, fsm_output(0));
  nand_41_nl <= NOT((fsm_output(4)) AND mux_1196_nl);
  mux_1200_nl <= MUX_s_1_2_2(mux_1199_nl, nand_41_nl, fsm_output(6));
  or_1211_nl <= (fsm_output(2)) OR mux_1200_nl;
  mux_1210_nl <= MUX_s_1_2_2(mux_1209_nl, or_1211_nl, fsm_output(5));
  vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1210_nl) AND (fsm_output(1));
  nor_1260_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT and_763_cse));
  nor_1261_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_1222_nl <= MUX_s_1_2_2(nor_1260_nl, nor_1261_nl, fsm_output(0));
  nor_1262_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1263_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1221_nl <= MUX_s_1_2_2(nor_1262_nl, nor_1263_nl, fsm_output(0));
  mux_1223_nl <= MUX_s_1_2_2(mux_1222_nl, mux_1221_nl, fsm_output(4));
  nor_1264_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1265_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1219_nl <= MUX_s_1_2_2(nor_1264_nl, nor_1265_nl, fsm_output(0));
  nor_1266_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1267_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1218_nl <= MUX_s_1_2_2(nor_1266_nl, nor_1267_nl, fsm_output(0));
  mux_1220_nl <= MUX_s_1_2_2(mux_1219_nl, mux_1218_nl, fsm_output(4));
  mux_1224_nl <= MUX_s_1_2_2(mux_1223_nl, mux_1220_nl, fsm_output(6));
  nand_455_nl <= NOT((fsm_output(2)) AND mux_1224_nl);
  or_1231_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT and_763_cse);
  mux_1215_nl <= MUX_s_1_2_2(or_tmp_1117, or_1231_nl, fsm_output(0));
  or_1228_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1214_nl <= MUX_s_1_2_2(or_tmp_1113, or_1228_nl, fsm_output(0));
  mux_1216_nl <= MUX_s_1_2_2(mux_1215_nl, mux_1214_nl, fsm_output(4));
  or_1225_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1212_nl <= MUX_s_1_2_2(or_tmp_1111, or_1225_nl, fsm_output(0));
  or_1222_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1211_nl <= MUX_s_1_2_2(or_tmp_1107, or_1222_nl, fsm_output(0));
  mux_1213_nl <= MUX_s_1_2_2(mux_1212_nl, mux_1211_nl, fsm_output(4));
  mux_1217_nl <= MUX_s_1_2_2(mux_1216_nl, mux_1213_nl, fsm_output(6));
  or_4128_nl <= (fsm_output(2)) OR mux_1217_nl;
  mux_1225_nl <= MUX_s_1_2_2(nand_455_nl, or_4128_nl, fsm_output(5));
  vec_rsc_0_14_i_we_d_pff <= NOT(mux_1225_nl OR (fsm_output(1)));
  or_1264_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1263_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1238_nl <= MUX_s_1_2_2(or_1264_nl, or_1263_nl, fsm_output(0));
  or_1265_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1238_nl;
  or_1261_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001110")) OR (NOT and_763_cse);
  mux_1235_nl <= MUX_s_1_2_2(or_1261_nl, or_tmp_1117, fsm_output(0));
  or_1259_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001110")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1234_nl <= MUX_s_1_2_2(or_1259_nl, or_tmp_1113, fsm_output(0));
  mux_1236_nl <= MUX_s_1_2_2(mux_1235_nl, mux_1234_nl, fsm_output(4));
  or_1258_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001110")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1232_nl <= MUX_s_1_2_2(or_1258_nl, or_tmp_1111, fsm_output(0));
  or_1256_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001110")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1231_nl <= MUX_s_1_2_2(or_1256_nl, or_tmp_1107, fsm_output(0));
  mux_1233_nl <= MUX_s_1_2_2(mux_1232_nl, mux_1231_nl, fsm_output(4));
  mux_1237_nl <= MUX_s_1_2_2(mux_1236_nl, mux_1233_nl, fsm_output(6));
  mux_1239_nl <= MUX_s_1_2_2(or_1265_nl, mux_1237_nl, fsm_output(2));
  or_1254_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1252_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT and_763_cse);
  mux_1228_nl <= MUX_s_1_2_2(or_1254_nl, or_1252_nl, fsm_output(0));
  or_1250_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1249_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1227_nl <= MUX_s_1_2_2(or_1250_nl, or_1249_nl, fsm_output(0));
  mux_1229_nl <= MUX_s_1_2_2(mux_1228_nl, mux_1227_nl, fsm_output(4));
  nor_1258_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1259_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1226_nl <= MUX_s_1_2_2(nor_1258_nl, nor_1259_nl, fsm_output(0));
  nand_43_nl <= NOT((fsm_output(4)) AND mux_1226_nl);
  mux_1230_nl <= MUX_s_1_2_2(mux_1229_nl, nand_43_nl, fsm_output(6));
  or_1255_nl <= (fsm_output(2)) OR mux_1230_nl;
  mux_1240_nl <= MUX_s_1_2_2(mux_1239_nl, or_1255_nl, fsm_output(5));
  vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1240_nl) AND (fsm_output(1));
  and_618_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001111"))
      AND and_763_cse;
  nor_1250_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001"))
      OR not_tmp_347);
  mux_1252_nl <= MUX_s_1_2_2(and_618_nl, nor_1250_nl, fsm_output(0));
  nor_1251_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1252_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1251_nl <= MUX_s_1_2_2(nor_1251_nl, nor_1252_nl, fsm_output(0));
  mux_1253_nl <= MUX_s_1_2_2(mux_1252_nl, mux_1251_nl, fsm_output(4));
  nor_1253_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1254_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1249_nl <= MUX_s_1_2_2(nor_1253_nl, nor_1254_nl, fsm_output(0));
  nor_1255_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1256_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1248_nl <= MUX_s_1_2_2(nor_1255_nl, nor_1256_nl, fsm_output(0));
  mux_1250_nl <= MUX_s_1_2_2(mux_1249_nl, mux_1248_nl, fsm_output(4));
  mux_1254_nl <= MUX_s_1_2_2(mux_1253_nl, mux_1250_nl, fsm_output(6));
  nand_454_nl <= NOT((fsm_output(2)) AND mux_1254_nl);
  nand_332_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001111"))
      AND and_763_cse);
  mux_1245_nl <= MUX_s_1_2_2(or_tmp_1161, nand_332_nl, fsm_output(0));
  or_1272_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1244_nl <= MUX_s_1_2_2(or_tmp_1157, or_1272_nl, fsm_output(0));
  mux_1246_nl <= MUX_s_1_2_2(mux_1245_nl, mux_1244_nl, fsm_output(4));
  or_1269_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1242_nl <= MUX_s_1_2_2(or_tmp_1155, or_1269_nl, fsm_output(0));
  or_1266_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1241_nl <= MUX_s_1_2_2(or_tmp_1151, or_1266_nl, fsm_output(0));
  mux_1243_nl <= MUX_s_1_2_2(mux_1242_nl, mux_1241_nl, fsm_output(4));
  mux_1247_nl <= MUX_s_1_2_2(mux_1246_nl, mux_1243_nl, fsm_output(6));
  or_4127_nl <= (fsm_output(2)) OR mux_1247_nl;
  mux_1255_nl <= MUX_s_1_2_2(nand_454_nl, or_4127_nl, fsm_output(5));
  vec_rsc_0_15_i_we_d_pff <= NOT(mux_1255_nl OR (fsm_output(1)));
  or_1308_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1307_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1268_nl <= MUX_s_1_2_2(or_1308_nl, or_1307_nl, fsm_output(0));
  or_1309_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1268_nl;
  nand_330_nl <= NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("001111")) AND and_763_cse);
  mux_1265_nl <= MUX_s_1_2_2(nand_330_nl, or_tmp_1161, fsm_output(0));
  or_1303_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001111")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1264_nl <= MUX_s_1_2_2(or_1303_nl, or_tmp_1157, fsm_output(0));
  mux_1266_nl <= MUX_s_1_2_2(mux_1265_nl, mux_1264_nl, fsm_output(4));
  or_1302_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001111")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1262_nl <= MUX_s_1_2_2(or_1302_nl, or_tmp_1155, fsm_output(0));
  or_1300_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001111")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1261_nl <= MUX_s_1_2_2(or_1300_nl, or_tmp_1151, fsm_output(0));
  mux_1263_nl <= MUX_s_1_2_2(mux_1262_nl, mux_1261_nl, fsm_output(4));
  mux_1267_nl <= MUX_s_1_2_2(mux_1266_nl, mux_1263_nl, fsm_output(6));
  mux_1269_nl <= MUX_s_1_2_2(or_1309_nl, mux_1267_nl, fsm_output(2));
  or_1298_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  nand_331_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("001111"))
      AND and_763_cse);
  mux_1258_nl <= MUX_s_1_2_2(or_1298_nl, nand_331_nl, fsm_output(0));
  or_1294_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1293_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1257_nl <= MUX_s_1_2_2(or_1294_nl, or_1293_nl, fsm_output(0));
  mux_1259_nl <= MUX_s_1_2_2(mux_1258_nl, mux_1257_nl, fsm_output(4));
  nor_1248_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1249_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1256_nl <= MUX_s_1_2_2(nor_1248_nl, nor_1249_nl, fsm_output(0));
  nand_45_nl <= NOT((fsm_output(4)) AND mux_1256_nl);
  mux_1260_nl <= MUX_s_1_2_2(mux_1259_nl, nand_45_nl, fsm_output(6));
  or_1299_nl <= (fsm_output(2)) OR mux_1260_nl;
  mux_1270_nl <= MUX_s_1_2_2(mux_1269_nl, or_1299_nl, fsm_output(5));
  vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1270_nl) AND (fsm_output(1));
  nor_1239_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1240_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_1282_nl <= MUX_s_1_2_2(nor_1239_nl, nor_1240_nl, fsm_output(0));
  nor_1241_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1242_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1281_nl <= MUX_s_1_2_2(nor_1241_nl, nor_1242_nl, fsm_output(0));
  mux_1283_nl <= MUX_s_1_2_2(mux_1282_nl, mux_1281_nl, fsm_output(4));
  nor_1243_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1244_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1279_nl <= MUX_s_1_2_2(nor_1243_nl, nor_1244_nl, fsm_output(0));
  nor_1245_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1246_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1278_nl <= MUX_s_1_2_2(nor_1245_nl, nor_1246_nl, fsm_output(0));
  mux_1280_nl <= MUX_s_1_2_2(mux_1279_nl, mux_1278_nl, fsm_output(4));
  mux_1284_nl <= MUX_s_1_2_2(mux_1283_nl, mux_1280_nl, fsm_output(6));
  nand_453_nl <= NOT((fsm_output(2)) AND mux_1284_nl);
  or_1319_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (NOT and_763_cse);
  mux_1275_nl <= MUX_s_1_2_2(or_tmp_1205, or_1319_nl, fsm_output(0));
  or_1316_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1274_nl <= MUX_s_1_2_2(or_tmp_1201, or_1316_nl, fsm_output(0));
  mux_1276_nl <= MUX_s_1_2_2(mux_1275_nl, mux_1274_nl, fsm_output(4));
  or_1313_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1272_nl <= MUX_s_1_2_2(or_tmp_1199, or_1313_nl, fsm_output(0));
  or_1310_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1271_nl <= MUX_s_1_2_2(or_tmp_1195, or_1310_nl, fsm_output(0));
  mux_1273_nl <= MUX_s_1_2_2(mux_1272_nl, mux_1271_nl, fsm_output(4));
  mux_1277_nl <= MUX_s_1_2_2(mux_1276_nl, mux_1273_nl, fsm_output(6));
  or_4126_nl <= (fsm_output(2)) OR mux_1277_nl;
  mux_1285_nl <= MUX_s_1_2_2(nand_453_nl, or_4126_nl, fsm_output(5));
  vec_rsc_0_16_i_we_d_pff <= NOT(mux_1285_nl OR (fsm_output(1)));
  or_1352_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1351_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1298_nl <= MUX_s_1_2_2(or_1352_nl, or_1351_nl, fsm_output(0));
  or_1353_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1298_nl;
  or_1349_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010000")) OR (NOT and_763_cse);
  mux_1295_nl <= MUX_s_1_2_2(or_1349_nl, or_tmp_1205, fsm_output(0));
  or_1347_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010000")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1294_nl <= MUX_s_1_2_2(or_1347_nl, or_tmp_1201, fsm_output(0));
  mux_1296_nl <= MUX_s_1_2_2(mux_1295_nl, mux_1294_nl, fsm_output(4));
  or_1346_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010000")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1292_nl <= MUX_s_1_2_2(or_1346_nl, or_tmp_1199, fsm_output(0));
  or_1344_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010000")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1291_nl <= MUX_s_1_2_2(or_1344_nl, or_tmp_1195, fsm_output(0));
  mux_1293_nl <= MUX_s_1_2_2(mux_1292_nl, mux_1291_nl, fsm_output(4));
  mux_1297_nl <= MUX_s_1_2_2(mux_1296_nl, mux_1293_nl, fsm_output(6));
  mux_1299_nl <= MUX_s_1_2_2(or_1353_nl, mux_1297_nl, fsm_output(2));
  or_1342_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1340_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1288_nl <= MUX_s_1_2_2(or_1342_nl, or_1340_nl, fsm_output(0));
  or_1338_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1337_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1287_nl <= MUX_s_1_2_2(or_1338_nl, or_1337_nl, fsm_output(0));
  mux_1289_nl <= MUX_s_1_2_2(mux_1288_nl, mux_1287_nl, fsm_output(4));
  nor_1237_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1238_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1286_nl <= MUX_s_1_2_2(nor_1237_nl, nor_1238_nl, fsm_output(0));
  nand_47_nl <= NOT((fsm_output(4)) AND mux_1286_nl);
  mux_1290_nl <= MUX_s_1_2_2(mux_1289_nl, nand_47_nl, fsm_output(6));
  or_1343_nl <= (fsm_output(2)) OR mux_1290_nl;
  mux_1300_nl <= MUX_s_1_2_2(mux_1299_nl, or_1343_nl, fsm_output(5));
  vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1300_nl) AND (fsm_output(1));
  nor_1228_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1229_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_1312_nl <= MUX_s_1_2_2(nor_1228_nl, nor_1229_nl, fsm_output(0));
  nor_1230_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1231_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1311_nl <= MUX_s_1_2_2(nor_1230_nl, nor_1231_nl, fsm_output(0));
  mux_1313_nl <= MUX_s_1_2_2(mux_1312_nl, mux_1311_nl, fsm_output(4));
  nor_1232_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1233_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1309_nl <= MUX_s_1_2_2(nor_1232_nl, nor_1233_nl, fsm_output(0));
  nor_1234_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1235_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1308_nl <= MUX_s_1_2_2(nor_1234_nl, nor_1235_nl, fsm_output(0));
  mux_1310_nl <= MUX_s_1_2_2(mux_1309_nl, mux_1308_nl, fsm_output(4));
  mux_1314_nl <= MUX_s_1_2_2(mux_1313_nl, mux_1310_nl, fsm_output(6));
  nand_452_nl <= NOT((fsm_output(2)) AND mux_1314_nl);
  or_1363_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (NOT and_763_cse);
  mux_1305_nl <= MUX_s_1_2_2(or_tmp_1249, or_1363_nl, fsm_output(0));
  or_1360_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1304_nl <= MUX_s_1_2_2(or_tmp_1245, or_1360_nl, fsm_output(0));
  mux_1306_nl <= MUX_s_1_2_2(mux_1305_nl, mux_1304_nl, fsm_output(4));
  or_1357_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1302_nl <= MUX_s_1_2_2(or_tmp_1243, or_1357_nl, fsm_output(0));
  or_1354_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1301_nl <= MUX_s_1_2_2(or_tmp_1239, or_1354_nl, fsm_output(0));
  mux_1303_nl <= MUX_s_1_2_2(mux_1302_nl, mux_1301_nl, fsm_output(4));
  mux_1307_nl <= MUX_s_1_2_2(mux_1306_nl, mux_1303_nl, fsm_output(6));
  or_4125_nl <= (fsm_output(2)) OR mux_1307_nl;
  mux_1315_nl <= MUX_s_1_2_2(nand_452_nl, or_4125_nl, fsm_output(5));
  vec_rsc_0_17_i_we_d_pff <= NOT(mux_1315_nl OR (fsm_output(1)));
  or_1396_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1395_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1328_nl <= MUX_s_1_2_2(or_1396_nl, or_1395_nl, fsm_output(0));
  or_1397_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1328_nl;
  or_1393_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010001")) OR (NOT and_763_cse);
  mux_1325_nl <= MUX_s_1_2_2(or_1393_nl, or_tmp_1249, fsm_output(0));
  or_1391_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010001")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1324_nl <= MUX_s_1_2_2(or_1391_nl, or_tmp_1245, fsm_output(0));
  mux_1326_nl <= MUX_s_1_2_2(mux_1325_nl, mux_1324_nl, fsm_output(4));
  or_1390_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010001")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1322_nl <= MUX_s_1_2_2(or_1390_nl, or_tmp_1243, fsm_output(0));
  or_1388_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010001")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1321_nl <= MUX_s_1_2_2(or_1388_nl, or_tmp_1239, fsm_output(0));
  mux_1323_nl <= MUX_s_1_2_2(mux_1322_nl, mux_1321_nl, fsm_output(4));
  mux_1327_nl <= MUX_s_1_2_2(mux_1326_nl, mux_1323_nl, fsm_output(6));
  mux_1329_nl <= MUX_s_1_2_2(or_1397_nl, mux_1327_nl, fsm_output(2));
  or_1386_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1384_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1318_nl <= MUX_s_1_2_2(or_1386_nl, or_1384_nl, fsm_output(0));
  or_1382_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1381_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1317_nl <= MUX_s_1_2_2(or_1382_nl, or_1381_nl, fsm_output(0));
  mux_1319_nl <= MUX_s_1_2_2(mux_1318_nl, mux_1317_nl, fsm_output(4));
  nor_1226_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1227_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1316_nl <= MUX_s_1_2_2(nor_1226_nl, nor_1227_nl, fsm_output(0));
  nand_49_nl <= NOT((fsm_output(4)) AND mux_1316_nl);
  mux_1320_nl <= MUX_s_1_2_2(mux_1319_nl, nand_49_nl, fsm_output(6));
  or_1387_nl <= (fsm_output(2)) OR mux_1320_nl;
  mux_1330_nl <= MUX_s_1_2_2(mux_1329_nl, or_1387_nl, fsm_output(5));
  vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1330_nl) AND (fsm_output(1));
  nor_1217_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1218_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_1342_nl <= MUX_s_1_2_2(nor_1217_nl, nor_1218_nl, fsm_output(0));
  nor_1219_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1220_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1341_nl <= MUX_s_1_2_2(nor_1219_nl, nor_1220_nl, fsm_output(0));
  mux_1343_nl <= MUX_s_1_2_2(mux_1342_nl, mux_1341_nl, fsm_output(4));
  nor_1221_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1222_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1339_nl <= MUX_s_1_2_2(nor_1221_nl, nor_1222_nl, fsm_output(0));
  nor_1223_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1224_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1338_nl <= MUX_s_1_2_2(nor_1223_nl, nor_1224_nl, fsm_output(0));
  mux_1340_nl <= MUX_s_1_2_2(mux_1339_nl, mux_1338_nl, fsm_output(4));
  mux_1344_nl <= MUX_s_1_2_2(mux_1343_nl, mux_1340_nl, fsm_output(6));
  nand_451_nl <= NOT((fsm_output(2)) AND mux_1344_nl);
  or_1407_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (NOT and_763_cse);
  mux_1335_nl <= MUX_s_1_2_2(or_tmp_1293, or_1407_nl, fsm_output(0));
  or_1404_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1334_nl <= MUX_s_1_2_2(or_tmp_1289, or_1404_nl, fsm_output(0));
  mux_1336_nl <= MUX_s_1_2_2(mux_1335_nl, mux_1334_nl, fsm_output(4));
  or_1401_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1332_nl <= MUX_s_1_2_2(or_tmp_1287, or_1401_nl, fsm_output(0));
  or_1398_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1331_nl <= MUX_s_1_2_2(or_tmp_1283, or_1398_nl, fsm_output(0));
  mux_1333_nl <= MUX_s_1_2_2(mux_1332_nl, mux_1331_nl, fsm_output(4));
  mux_1337_nl <= MUX_s_1_2_2(mux_1336_nl, mux_1333_nl, fsm_output(6));
  or_4124_nl <= (fsm_output(2)) OR mux_1337_nl;
  mux_1345_nl <= MUX_s_1_2_2(nand_451_nl, or_4124_nl, fsm_output(5));
  vec_rsc_0_18_i_we_d_pff <= NOT(mux_1345_nl OR (fsm_output(1)));
  or_1440_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1439_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1358_nl <= MUX_s_1_2_2(or_1440_nl, or_1439_nl, fsm_output(0));
  or_1441_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1358_nl;
  or_1437_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010010")) OR (NOT and_763_cse);
  mux_1355_nl <= MUX_s_1_2_2(or_1437_nl, or_tmp_1293, fsm_output(0));
  or_1435_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010010")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1354_nl <= MUX_s_1_2_2(or_1435_nl, or_tmp_1289, fsm_output(0));
  mux_1356_nl <= MUX_s_1_2_2(mux_1355_nl, mux_1354_nl, fsm_output(4));
  or_1434_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010010")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1352_nl <= MUX_s_1_2_2(or_1434_nl, or_tmp_1287, fsm_output(0));
  or_1432_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010010")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1351_nl <= MUX_s_1_2_2(or_1432_nl, or_tmp_1283, fsm_output(0));
  mux_1353_nl <= MUX_s_1_2_2(mux_1352_nl, mux_1351_nl, fsm_output(4));
  mux_1357_nl <= MUX_s_1_2_2(mux_1356_nl, mux_1353_nl, fsm_output(6));
  mux_1359_nl <= MUX_s_1_2_2(or_1441_nl, mux_1357_nl, fsm_output(2));
  or_1430_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1428_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1348_nl <= MUX_s_1_2_2(or_1430_nl, or_1428_nl, fsm_output(0));
  or_1426_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1425_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1347_nl <= MUX_s_1_2_2(or_1426_nl, or_1425_nl, fsm_output(0));
  mux_1349_nl <= MUX_s_1_2_2(mux_1348_nl, mux_1347_nl, fsm_output(4));
  nor_1215_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1216_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1346_nl <= MUX_s_1_2_2(nor_1215_nl, nor_1216_nl, fsm_output(0));
  nand_51_nl <= NOT((fsm_output(4)) AND mux_1346_nl);
  mux_1350_nl <= MUX_s_1_2_2(mux_1349_nl, nand_51_nl, fsm_output(6));
  or_1431_nl <= (fsm_output(2)) OR mux_1350_nl;
  mux_1360_nl <= MUX_s_1_2_2(mux_1359_nl, or_1431_nl, fsm_output(5));
  vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1360_nl) AND (fsm_output(1));
  nor_1206_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1207_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR not_tmp_330);
  mux_1372_nl <= MUX_s_1_2_2(nor_1206_nl, nor_1207_nl, fsm_output(0));
  nor_1208_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1209_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1371_nl <= MUX_s_1_2_2(nor_1208_nl, nor_1209_nl, fsm_output(0));
  mux_1373_nl <= MUX_s_1_2_2(mux_1372_nl, mux_1371_nl, fsm_output(4));
  nor_1210_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1211_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1369_nl <= MUX_s_1_2_2(nor_1210_nl, nor_1211_nl, fsm_output(0));
  nor_1212_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1213_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1368_nl <= MUX_s_1_2_2(nor_1212_nl, nor_1213_nl, fsm_output(0));
  mux_1370_nl <= MUX_s_1_2_2(mux_1369_nl, mux_1368_nl, fsm_output(4));
  mux_1374_nl <= MUX_s_1_2_2(mux_1373_nl, mux_1370_nl, fsm_output(6));
  nand_450_nl <= NOT((fsm_output(2)) AND mux_1374_nl);
  or_1451_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (NOT and_763_cse);
  mux_1365_nl <= MUX_s_1_2_2(or_tmp_1337, or_1451_nl, fsm_output(0));
  or_1448_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1364_nl <= MUX_s_1_2_2(or_tmp_1333, or_1448_nl, fsm_output(0));
  mux_1366_nl <= MUX_s_1_2_2(mux_1365_nl, mux_1364_nl, fsm_output(4));
  or_1445_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1362_nl <= MUX_s_1_2_2(or_tmp_1331, or_1445_nl, fsm_output(0));
  or_1442_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1361_nl <= MUX_s_1_2_2(or_tmp_1327, or_1442_nl, fsm_output(0));
  mux_1363_nl <= MUX_s_1_2_2(mux_1362_nl, mux_1361_nl, fsm_output(4));
  mux_1367_nl <= MUX_s_1_2_2(mux_1366_nl, mux_1363_nl, fsm_output(6));
  or_4123_nl <= (fsm_output(2)) OR mux_1367_nl;
  mux_1375_nl <= MUX_s_1_2_2(nand_450_nl, or_4123_nl, fsm_output(5));
  vec_rsc_0_19_i_we_d_pff <= NOT(mux_1375_nl OR (fsm_output(1)));
  or_1484_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1483_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1388_nl <= MUX_s_1_2_2(or_1484_nl, or_1483_nl, fsm_output(0));
  or_1485_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1388_nl;
  or_1481_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010011")) OR (NOT and_763_cse);
  mux_1385_nl <= MUX_s_1_2_2(or_1481_nl, or_tmp_1337, fsm_output(0));
  or_1479_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010011")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1384_nl <= MUX_s_1_2_2(or_1479_nl, or_tmp_1333, fsm_output(0));
  mux_1386_nl <= MUX_s_1_2_2(mux_1385_nl, mux_1384_nl, fsm_output(4));
  or_1478_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010011")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1382_nl <= MUX_s_1_2_2(or_1478_nl, or_tmp_1331, fsm_output(0));
  or_1476_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010011")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1381_nl <= MUX_s_1_2_2(or_1476_nl, or_tmp_1327, fsm_output(0));
  mux_1383_nl <= MUX_s_1_2_2(mux_1382_nl, mux_1381_nl, fsm_output(4));
  mux_1387_nl <= MUX_s_1_2_2(mux_1386_nl, mux_1383_nl, fsm_output(6));
  mux_1389_nl <= MUX_s_1_2_2(or_1485_nl, mux_1387_nl, fsm_output(2));
  or_1474_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1472_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1378_nl <= MUX_s_1_2_2(or_1474_nl, or_1472_nl, fsm_output(0));
  or_1470_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1469_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1377_nl <= MUX_s_1_2_2(or_1470_nl, or_1469_nl, fsm_output(0));
  mux_1379_nl <= MUX_s_1_2_2(mux_1378_nl, mux_1377_nl, fsm_output(4));
  nor_1204_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1205_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1376_nl <= MUX_s_1_2_2(nor_1204_nl, nor_1205_nl, fsm_output(0));
  nand_53_nl <= NOT((fsm_output(4)) AND mux_1376_nl);
  mux_1380_nl <= MUX_s_1_2_2(mux_1379_nl, nand_53_nl, fsm_output(6));
  or_1475_nl <= (fsm_output(2)) OR mux_1380_nl;
  mux_1390_nl <= MUX_s_1_2_2(mux_1389_nl, or_1475_nl, fsm_output(5));
  vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1390_nl) AND (fsm_output(1));
  nor_1195_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1196_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_1402_nl <= MUX_s_1_2_2(nor_1195_nl, nor_1196_nl, fsm_output(0));
  nor_1197_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1198_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1401_nl <= MUX_s_1_2_2(nor_1197_nl, nor_1198_nl, fsm_output(0));
  mux_1403_nl <= MUX_s_1_2_2(mux_1402_nl, mux_1401_nl, fsm_output(4));
  nor_1199_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1200_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1399_nl <= MUX_s_1_2_2(nor_1199_nl, nor_1200_nl, fsm_output(0));
  nor_1201_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1202_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1398_nl <= MUX_s_1_2_2(nor_1201_nl, nor_1202_nl, fsm_output(0));
  mux_1400_nl <= MUX_s_1_2_2(mux_1399_nl, mux_1398_nl, fsm_output(4));
  mux_1404_nl <= MUX_s_1_2_2(mux_1403_nl, mux_1400_nl, fsm_output(6));
  nand_449_nl <= NOT((fsm_output(2)) AND mux_1404_nl);
  or_1495_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (NOT and_763_cse);
  mux_1395_nl <= MUX_s_1_2_2(or_tmp_1381, or_1495_nl, fsm_output(0));
  or_1492_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1394_nl <= MUX_s_1_2_2(or_tmp_1377, or_1492_nl, fsm_output(0));
  mux_1396_nl <= MUX_s_1_2_2(mux_1395_nl, mux_1394_nl, fsm_output(4));
  or_1489_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1392_nl <= MUX_s_1_2_2(or_tmp_1375, or_1489_nl, fsm_output(0));
  or_1486_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1391_nl <= MUX_s_1_2_2(or_tmp_1371, or_1486_nl, fsm_output(0));
  mux_1393_nl <= MUX_s_1_2_2(mux_1392_nl, mux_1391_nl, fsm_output(4));
  mux_1397_nl <= MUX_s_1_2_2(mux_1396_nl, mux_1393_nl, fsm_output(6));
  or_4122_nl <= (fsm_output(2)) OR mux_1397_nl;
  mux_1405_nl <= MUX_s_1_2_2(nand_449_nl, or_4122_nl, fsm_output(5));
  vec_rsc_0_20_i_we_d_pff <= NOT(mux_1405_nl OR (fsm_output(1)));
  or_1528_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1527_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1418_nl <= MUX_s_1_2_2(or_1528_nl, or_1527_nl, fsm_output(0));
  or_1529_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1418_nl;
  or_1525_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010100")) OR (NOT and_763_cse);
  mux_1415_nl <= MUX_s_1_2_2(or_1525_nl, or_tmp_1381, fsm_output(0));
  or_1523_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010100")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1414_nl <= MUX_s_1_2_2(or_1523_nl, or_tmp_1377, fsm_output(0));
  mux_1416_nl <= MUX_s_1_2_2(mux_1415_nl, mux_1414_nl, fsm_output(4));
  or_1522_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010100")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1412_nl <= MUX_s_1_2_2(or_1522_nl, or_tmp_1375, fsm_output(0));
  or_1520_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010100")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1411_nl <= MUX_s_1_2_2(or_1520_nl, or_tmp_1371, fsm_output(0));
  mux_1413_nl <= MUX_s_1_2_2(mux_1412_nl, mux_1411_nl, fsm_output(4));
  mux_1417_nl <= MUX_s_1_2_2(mux_1416_nl, mux_1413_nl, fsm_output(6));
  mux_1419_nl <= MUX_s_1_2_2(or_1529_nl, mux_1417_nl, fsm_output(2));
  or_1518_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1516_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1408_nl <= MUX_s_1_2_2(or_1518_nl, or_1516_nl, fsm_output(0));
  or_1514_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1513_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1407_nl <= MUX_s_1_2_2(or_1514_nl, or_1513_nl, fsm_output(0));
  mux_1409_nl <= MUX_s_1_2_2(mux_1408_nl, mux_1407_nl, fsm_output(4));
  nor_1193_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1194_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1406_nl <= MUX_s_1_2_2(nor_1193_nl, nor_1194_nl, fsm_output(0));
  nand_55_nl <= NOT((fsm_output(4)) AND mux_1406_nl);
  mux_1410_nl <= MUX_s_1_2_2(mux_1409_nl, nand_55_nl, fsm_output(6));
  or_1519_nl <= (fsm_output(2)) OR mux_1410_nl;
  mux_1420_nl <= MUX_s_1_2_2(mux_1419_nl, or_1519_nl, fsm_output(5));
  vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1420_nl) AND (fsm_output(1));
  nor_1184_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1185_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_1432_nl <= MUX_s_1_2_2(nor_1184_nl, nor_1185_nl, fsm_output(0));
  nor_1186_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1187_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1431_nl <= MUX_s_1_2_2(nor_1186_nl, nor_1187_nl, fsm_output(0));
  mux_1433_nl <= MUX_s_1_2_2(mux_1432_nl, mux_1431_nl, fsm_output(4));
  nor_1188_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1189_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1429_nl <= MUX_s_1_2_2(nor_1188_nl, nor_1189_nl, fsm_output(0));
  nor_1190_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1191_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1428_nl <= MUX_s_1_2_2(nor_1190_nl, nor_1191_nl, fsm_output(0));
  mux_1430_nl <= MUX_s_1_2_2(mux_1429_nl, mux_1428_nl, fsm_output(4));
  mux_1434_nl <= MUX_s_1_2_2(mux_1433_nl, mux_1430_nl, fsm_output(6));
  nand_448_nl <= NOT((fsm_output(2)) AND mux_1434_nl);
  or_1539_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (NOT and_763_cse);
  mux_1425_nl <= MUX_s_1_2_2(or_tmp_1425, or_1539_nl, fsm_output(0));
  or_1536_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1424_nl <= MUX_s_1_2_2(or_tmp_1421, or_1536_nl, fsm_output(0));
  mux_1426_nl <= MUX_s_1_2_2(mux_1425_nl, mux_1424_nl, fsm_output(4));
  or_1533_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1422_nl <= MUX_s_1_2_2(or_tmp_1419, or_1533_nl, fsm_output(0));
  or_1530_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1421_nl <= MUX_s_1_2_2(or_tmp_1415, or_1530_nl, fsm_output(0));
  mux_1423_nl <= MUX_s_1_2_2(mux_1422_nl, mux_1421_nl, fsm_output(4));
  mux_1427_nl <= MUX_s_1_2_2(mux_1426_nl, mux_1423_nl, fsm_output(6));
  or_4121_nl <= (fsm_output(2)) OR mux_1427_nl;
  mux_1435_nl <= MUX_s_1_2_2(nand_448_nl, or_4121_nl, fsm_output(5));
  vec_rsc_0_21_i_we_d_pff <= NOT(mux_1435_nl OR (fsm_output(1)));
  or_1572_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1571_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1448_nl <= MUX_s_1_2_2(or_1572_nl, or_1571_nl, fsm_output(0));
  or_1573_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1448_nl;
  or_1569_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010101")) OR (NOT and_763_cse);
  mux_1445_nl <= MUX_s_1_2_2(or_1569_nl, or_tmp_1425, fsm_output(0));
  or_1567_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010101")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1444_nl <= MUX_s_1_2_2(or_1567_nl, or_tmp_1421, fsm_output(0));
  mux_1446_nl <= MUX_s_1_2_2(mux_1445_nl, mux_1444_nl, fsm_output(4));
  or_1566_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010101")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1442_nl <= MUX_s_1_2_2(or_1566_nl, or_tmp_1419, fsm_output(0));
  or_1564_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010101")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1441_nl <= MUX_s_1_2_2(or_1564_nl, or_tmp_1415, fsm_output(0));
  mux_1443_nl <= MUX_s_1_2_2(mux_1442_nl, mux_1441_nl, fsm_output(4));
  mux_1447_nl <= MUX_s_1_2_2(mux_1446_nl, mux_1443_nl, fsm_output(6));
  mux_1449_nl <= MUX_s_1_2_2(or_1573_nl, mux_1447_nl, fsm_output(2));
  or_1562_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1560_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(0))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1438_nl <= MUX_s_1_2_2(or_1562_nl, or_1560_nl, fsm_output(0));
  or_1558_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1557_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1437_nl <= MUX_s_1_2_2(or_1558_nl, or_1557_nl, fsm_output(0));
  mux_1439_nl <= MUX_s_1_2_2(mux_1438_nl, mux_1437_nl, fsm_output(4));
  nor_1182_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1183_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1436_nl <= MUX_s_1_2_2(nor_1182_nl, nor_1183_nl, fsm_output(0));
  nand_57_nl <= NOT((fsm_output(4)) AND mux_1436_nl);
  mux_1440_nl <= MUX_s_1_2_2(mux_1439_nl, nand_57_nl, fsm_output(6));
  or_1563_nl <= (fsm_output(2)) OR mux_1440_nl;
  mux_1450_nl <= MUX_s_1_2_2(mux_1449_nl, or_1563_nl, fsm_output(5));
  vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1450_nl) AND (fsm_output(1));
  nor_1173_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1174_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_1462_nl <= MUX_s_1_2_2(nor_1173_nl, nor_1174_nl, fsm_output(0));
  nor_1175_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1176_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1461_nl <= MUX_s_1_2_2(nor_1175_nl, nor_1176_nl, fsm_output(0));
  mux_1463_nl <= MUX_s_1_2_2(mux_1462_nl, mux_1461_nl, fsm_output(4));
  nor_1177_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1178_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1459_nl <= MUX_s_1_2_2(nor_1177_nl, nor_1178_nl, fsm_output(0));
  nor_1179_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1180_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1458_nl <= MUX_s_1_2_2(nor_1179_nl, nor_1180_nl, fsm_output(0));
  mux_1460_nl <= MUX_s_1_2_2(mux_1459_nl, mux_1458_nl, fsm_output(4));
  mux_1464_nl <= MUX_s_1_2_2(mux_1463_nl, mux_1460_nl, fsm_output(6));
  nand_447_nl <= NOT((fsm_output(2)) AND mux_1464_nl);
  or_1583_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (NOT and_763_cse);
  mux_1455_nl <= MUX_s_1_2_2(or_tmp_1469, or_1583_nl, fsm_output(0));
  or_1580_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1454_nl <= MUX_s_1_2_2(or_tmp_1465, or_1580_nl, fsm_output(0));
  mux_1456_nl <= MUX_s_1_2_2(mux_1455_nl, mux_1454_nl, fsm_output(4));
  or_1577_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1452_nl <= MUX_s_1_2_2(or_tmp_1463, or_1577_nl, fsm_output(0));
  or_1574_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1451_nl <= MUX_s_1_2_2(or_tmp_1459, or_1574_nl, fsm_output(0));
  mux_1453_nl <= MUX_s_1_2_2(mux_1452_nl, mux_1451_nl, fsm_output(4));
  mux_1457_nl <= MUX_s_1_2_2(mux_1456_nl, mux_1453_nl, fsm_output(6));
  or_4120_nl <= (fsm_output(2)) OR mux_1457_nl;
  mux_1465_nl <= MUX_s_1_2_2(nand_447_nl, or_4120_nl, fsm_output(5));
  vec_rsc_0_22_i_we_d_pff <= NOT(mux_1465_nl OR (fsm_output(1)));
  or_1616_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1615_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1478_nl <= MUX_s_1_2_2(or_1616_nl, or_1615_nl, fsm_output(0));
  or_1617_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1478_nl;
  or_1613_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010110")) OR (NOT and_763_cse);
  mux_1475_nl <= MUX_s_1_2_2(or_1613_nl, or_tmp_1469, fsm_output(0));
  or_1611_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010110")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1474_nl <= MUX_s_1_2_2(or_1611_nl, or_tmp_1465, fsm_output(0));
  mux_1476_nl <= MUX_s_1_2_2(mux_1475_nl, mux_1474_nl, fsm_output(4));
  or_1610_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010110")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1472_nl <= MUX_s_1_2_2(or_1610_nl, or_tmp_1463, fsm_output(0));
  or_1608_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010110")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1471_nl <= MUX_s_1_2_2(or_1608_nl, or_tmp_1459, fsm_output(0));
  mux_1473_nl <= MUX_s_1_2_2(mux_1472_nl, mux_1471_nl, fsm_output(4));
  mux_1477_nl <= MUX_s_1_2_2(mux_1476_nl, mux_1473_nl, fsm_output(6));
  mux_1479_nl <= MUX_s_1_2_2(or_1617_nl, mux_1477_nl, fsm_output(2));
  or_1606_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1604_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1468_nl <= MUX_s_1_2_2(or_1606_nl, or_1604_nl, fsm_output(0));
  or_1602_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1601_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1467_nl <= MUX_s_1_2_2(or_1602_nl, or_1601_nl, fsm_output(0));
  mux_1469_nl <= MUX_s_1_2_2(mux_1468_nl, mux_1467_nl, fsm_output(4));
  nor_1171_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1172_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1466_nl <= MUX_s_1_2_2(nor_1171_nl, nor_1172_nl, fsm_output(0));
  nand_59_nl <= NOT((fsm_output(4)) AND mux_1466_nl);
  mux_1470_nl <= MUX_s_1_2_2(mux_1469_nl, nand_59_nl, fsm_output(6));
  or_1607_nl <= (fsm_output(2)) OR mux_1470_nl;
  mux_1480_nl <= MUX_s_1_2_2(mux_1479_nl, or_1607_nl, fsm_output(5));
  vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1480_nl) AND (fsm_output(1));
  nor_1162_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1163_nl <= NOT((COMP_LOOP_acc_13_psp_sva(3)) OR (COMP_LOOP_acc_13_psp_sva(1))
      OR not_tmp_414);
  mux_1492_nl <= MUX_s_1_2_2(nor_1162_nl, nor_1163_nl, fsm_output(0));
  nor_1164_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1165_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1491_nl <= MUX_s_1_2_2(nor_1164_nl, nor_1165_nl, fsm_output(0));
  mux_1493_nl <= MUX_s_1_2_2(mux_1492_nl, mux_1491_nl, fsm_output(4));
  nor_1166_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1167_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1489_nl <= MUX_s_1_2_2(nor_1166_nl, nor_1167_nl, fsm_output(0));
  nor_1168_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1169_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1488_nl <= MUX_s_1_2_2(nor_1168_nl, nor_1169_nl, fsm_output(0));
  mux_1490_nl <= MUX_s_1_2_2(mux_1489_nl, mux_1488_nl, fsm_output(4));
  mux_1494_nl <= MUX_s_1_2_2(mux_1493_nl, mux_1490_nl, fsm_output(6));
  nand_446_nl <= NOT((fsm_output(2)) AND mux_1494_nl);
  nand_326_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("010111"))
      AND and_763_cse);
  mux_1485_nl <= MUX_s_1_2_2(or_tmp_1513, nand_326_nl, fsm_output(0));
  or_1624_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1484_nl <= MUX_s_1_2_2(or_tmp_1509, or_1624_nl, fsm_output(0));
  mux_1486_nl <= MUX_s_1_2_2(mux_1485_nl, mux_1484_nl, fsm_output(4));
  or_1621_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1482_nl <= MUX_s_1_2_2(or_tmp_1507, or_1621_nl, fsm_output(0));
  or_1618_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1481_nl <= MUX_s_1_2_2(or_tmp_1503, or_1618_nl, fsm_output(0));
  mux_1483_nl <= MUX_s_1_2_2(mux_1482_nl, mux_1481_nl, fsm_output(4));
  mux_1487_nl <= MUX_s_1_2_2(mux_1486_nl, mux_1483_nl, fsm_output(6));
  or_4119_nl <= (fsm_output(2)) OR mux_1487_nl;
  mux_1495_nl <= MUX_s_1_2_2(nand_446_nl, or_4119_nl, fsm_output(5));
  vec_rsc_0_23_i_we_d_pff <= NOT(mux_1495_nl OR (fsm_output(1)));
  or_1660_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1659_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1508_nl <= MUX_s_1_2_2(or_1660_nl, or_1659_nl, fsm_output(0));
  or_1661_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1508_nl;
  nand_325_nl <= NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("010111")) AND and_763_cse);
  mux_1505_nl <= MUX_s_1_2_2(nand_325_nl, or_tmp_1513, fsm_output(0));
  or_1655_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010111")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1504_nl <= MUX_s_1_2_2(or_1655_nl, or_tmp_1509, fsm_output(0));
  mux_1506_nl <= MUX_s_1_2_2(mux_1505_nl, mux_1504_nl, fsm_output(4));
  or_1654_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010111")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1502_nl <= MUX_s_1_2_2(or_1654_nl, or_tmp_1507, fsm_output(0));
  or_1652_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010111")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1501_nl <= MUX_s_1_2_2(or_1652_nl, or_tmp_1503, fsm_output(0));
  mux_1503_nl <= MUX_s_1_2_2(mux_1502_nl, mux_1501_nl, fsm_output(4));
  mux_1507_nl <= MUX_s_1_2_2(mux_1506_nl, mux_1503_nl, fsm_output(6));
  mux_1509_nl <= MUX_s_1_2_2(or_1661_nl, mux_1507_nl, fsm_output(2));
  or_1650_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1648_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(0))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1498_nl <= MUX_s_1_2_2(or_1650_nl, or_1648_nl, fsm_output(0));
  or_1646_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1645_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1497_nl <= MUX_s_1_2_2(or_1646_nl, or_1645_nl, fsm_output(0));
  mux_1499_nl <= MUX_s_1_2_2(mux_1498_nl, mux_1497_nl, fsm_output(4));
  nor_1160_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1161_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1496_nl <= MUX_s_1_2_2(nor_1160_nl, nor_1161_nl, fsm_output(0));
  nand_61_nl <= NOT((fsm_output(4)) AND mux_1496_nl);
  mux_1500_nl <= MUX_s_1_2_2(mux_1499_nl, nand_61_nl, fsm_output(6));
  or_1651_nl <= (fsm_output(2)) OR mux_1500_nl;
  mux_1510_nl <= MUX_s_1_2_2(mux_1509_nl, or_1651_nl, fsm_output(5));
  vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1510_nl) AND (fsm_output(1));
  nor_1151_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1152_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_1522_nl <= MUX_s_1_2_2(nor_1151_nl, nor_1152_nl, fsm_output(0));
  nor_1153_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1154_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1521_nl <= MUX_s_1_2_2(nor_1153_nl, nor_1154_nl, fsm_output(0));
  mux_1523_nl <= MUX_s_1_2_2(mux_1522_nl, mux_1521_nl, fsm_output(4));
  nor_1155_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1156_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1519_nl <= MUX_s_1_2_2(nor_1155_nl, nor_1156_nl, fsm_output(0));
  nor_1157_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1158_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1518_nl <= MUX_s_1_2_2(nor_1157_nl, nor_1158_nl, fsm_output(0));
  mux_1520_nl <= MUX_s_1_2_2(mux_1519_nl, mux_1518_nl, fsm_output(4));
  mux_1524_nl <= MUX_s_1_2_2(mux_1523_nl, mux_1520_nl, fsm_output(6));
  nand_445_nl <= NOT((fsm_output(2)) AND mux_1524_nl);
  or_1671_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (NOT and_763_cse);
  mux_1515_nl <= MUX_s_1_2_2(or_tmp_1557, or_1671_nl, fsm_output(0));
  or_1668_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1514_nl <= MUX_s_1_2_2(or_tmp_1553, or_1668_nl, fsm_output(0));
  mux_1516_nl <= MUX_s_1_2_2(mux_1515_nl, mux_1514_nl, fsm_output(4));
  or_1665_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1512_nl <= MUX_s_1_2_2(or_tmp_1551, or_1665_nl, fsm_output(0));
  or_1662_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1511_nl <= MUX_s_1_2_2(or_tmp_1547, or_1662_nl, fsm_output(0));
  mux_1513_nl <= MUX_s_1_2_2(mux_1512_nl, mux_1511_nl, fsm_output(4));
  mux_1517_nl <= MUX_s_1_2_2(mux_1516_nl, mux_1513_nl, fsm_output(6));
  or_4118_nl <= (fsm_output(2)) OR mux_1517_nl;
  mux_1525_nl <= MUX_s_1_2_2(nand_445_nl, or_4118_nl, fsm_output(5));
  vec_rsc_0_24_i_we_d_pff <= NOT(mux_1525_nl OR (fsm_output(1)));
  or_1704_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1703_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1538_nl <= MUX_s_1_2_2(or_1704_nl, or_1703_nl, fsm_output(0));
  or_1705_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1538_nl;
  or_1701_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011000")) OR (NOT and_763_cse);
  mux_1535_nl <= MUX_s_1_2_2(or_1701_nl, or_tmp_1557, fsm_output(0));
  or_1699_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011000")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1534_nl <= MUX_s_1_2_2(or_1699_nl, or_tmp_1553, fsm_output(0));
  mux_1536_nl <= MUX_s_1_2_2(mux_1535_nl, mux_1534_nl, fsm_output(4));
  or_1698_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011000")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1532_nl <= MUX_s_1_2_2(or_1698_nl, or_tmp_1551, fsm_output(0));
  or_1696_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011000")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1531_nl <= MUX_s_1_2_2(or_1696_nl, or_tmp_1547, fsm_output(0));
  mux_1533_nl <= MUX_s_1_2_2(mux_1532_nl, mux_1531_nl, fsm_output(4));
  mux_1537_nl <= MUX_s_1_2_2(mux_1536_nl, mux_1533_nl, fsm_output(6));
  mux_1539_nl <= MUX_s_1_2_2(or_1705_nl, mux_1537_nl, fsm_output(2));
  or_1694_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1692_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1528_nl <= MUX_s_1_2_2(or_1694_nl, or_1692_nl, fsm_output(0));
  or_1690_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1689_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1527_nl <= MUX_s_1_2_2(or_1690_nl, or_1689_nl, fsm_output(0));
  mux_1529_nl <= MUX_s_1_2_2(mux_1528_nl, mux_1527_nl, fsm_output(4));
  nor_1149_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1150_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1526_nl <= MUX_s_1_2_2(nor_1149_nl, nor_1150_nl, fsm_output(0));
  nand_63_nl <= NOT((fsm_output(4)) AND mux_1526_nl);
  mux_1530_nl <= MUX_s_1_2_2(mux_1529_nl, nand_63_nl, fsm_output(6));
  or_1695_nl <= (fsm_output(2)) OR mux_1530_nl;
  mux_1540_nl <= MUX_s_1_2_2(mux_1539_nl, or_1695_nl, fsm_output(5));
  vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1540_nl) AND (fsm_output(1));
  nor_1140_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1141_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_1552_nl <= MUX_s_1_2_2(nor_1140_nl, nor_1141_nl, fsm_output(0));
  nor_1142_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1143_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1551_nl <= MUX_s_1_2_2(nor_1142_nl, nor_1143_nl, fsm_output(0));
  mux_1553_nl <= MUX_s_1_2_2(mux_1552_nl, mux_1551_nl, fsm_output(4));
  nor_1144_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1145_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1549_nl <= MUX_s_1_2_2(nor_1144_nl, nor_1145_nl, fsm_output(0));
  nor_1146_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1147_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1548_nl <= MUX_s_1_2_2(nor_1146_nl, nor_1147_nl, fsm_output(0));
  mux_1550_nl <= MUX_s_1_2_2(mux_1549_nl, mux_1548_nl, fsm_output(4));
  mux_1554_nl <= MUX_s_1_2_2(mux_1553_nl, mux_1550_nl, fsm_output(6));
  nand_444_nl <= NOT((fsm_output(2)) AND mux_1554_nl);
  or_1715_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (NOT and_763_cse);
  mux_1545_nl <= MUX_s_1_2_2(or_tmp_1601, or_1715_nl, fsm_output(0));
  or_1712_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1544_nl <= MUX_s_1_2_2(or_tmp_1597, or_1712_nl, fsm_output(0));
  mux_1546_nl <= MUX_s_1_2_2(mux_1545_nl, mux_1544_nl, fsm_output(4));
  or_1709_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1542_nl <= MUX_s_1_2_2(or_tmp_1595, or_1709_nl, fsm_output(0));
  or_1706_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1541_nl <= MUX_s_1_2_2(or_tmp_1591, or_1706_nl, fsm_output(0));
  mux_1543_nl <= MUX_s_1_2_2(mux_1542_nl, mux_1541_nl, fsm_output(4));
  mux_1547_nl <= MUX_s_1_2_2(mux_1546_nl, mux_1543_nl, fsm_output(6));
  or_4117_nl <= (fsm_output(2)) OR mux_1547_nl;
  mux_1555_nl <= MUX_s_1_2_2(nand_444_nl, or_4117_nl, fsm_output(5));
  vec_rsc_0_25_i_we_d_pff <= NOT(mux_1555_nl OR (fsm_output(1)));
  or_1748_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1747_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1568_nl <= MUX_s_1_2_2(or_1748_nl, or_1747_nl, fsm_output(0));
  or_1749_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1568_nl;
  or_1745_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011001")) OR (NOT and_763_cse);
  mux_1565_nl <= MUX_s_1_2_2(or_1745_nl, or_tmp_1601, fsm_output(0));
  or_1743_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011001")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1564_nl <= MUX_s_1_2_2(or_1743_nl, or_tmp_1597, fsm_output(0));
  mux_1566_nl <= MUX_s_1_2_2(mux_1565_nl, mux_1564_nl, fsm_output(4));
  or_1742_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011001")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1562_nl <= MUX_s_1_2_2(or_1742_nl, or_tmp_1595, fsm_output(0));
  or_1740_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011001")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1561_nl <= MUX_s_1_2_2(or_1740_nl, or_tmp_1591, fsm_output(0));
  mux_1563_nl <= MUX_s_1_2_2(mux_1562_nl, mux_1561_nl, fsm_output(4));
  mux_1567_nl <= MUX_s_1_2_2(mux_1566_nl, mux_1563_nl, fsm_output(6));
  mux_1569_nl <= MUX_s_1_2_2(or_1749_nl, mux_1567_nl, fsm_output(2));
  or_1738_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1736_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1558_nl <= MUX_s_1_2_2(or_1738_nl, or_1736_nl, fsm_output(0));
  or_1734_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1733_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1557_nl <= MUX_s_1_2_2(or_1734_nl, or_1733_nl, fsm_output(0));
  mux_1559_nl <= MUX_s_1_2_2(mux_1558_nl, mux_1557_nl, fsm_output(4));
  nor_1138_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1139_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1556_nl <= MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, fsm_output(0));
  nand_65_nl <= NOT((fsm_output(4)) AND mux_1556_nl);
  mux_1560_nl <= MUX_s_1_2_2(mux_1559_nl, nand_65_nl, fsm_output(6));
  or_1739_nl <= (fsm_output(2)) OR mux_1560_nl;
  mux_1570_nl <= MUX_s_1_2_2(mux_1569_nl, or_1739_nl, fsm_output(5));
  vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1570_nl) AND (fsm_output(1));
  nor_1129_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(1))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1130_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_1582_nl <= MUX_s_1_2_2(nor_1129_nl, nor_1130_nl, fsm_output(0));
  nor_1131_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1132_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1581_nl <= MUX_s_1_2_2(nor_1131_nl, nor_1132_nl, fsm_output(0));
  mux_1583_nl <= MUX_s_1_2_2(mux_1582_nl, mux_1581_nl, fsm_output(4));
  nor_1133_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1134_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1579_nl <= MUX_s_1_2_2(nor_1133_nl, nor_1134_nl, fsm_output(0));
  nor_1135_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1136_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1578_nl <= MUX_s_1_2_2(nor_1135_nl, nor_1136_nl, fsm_output(0));
  mux_1580_nl <= MUX_s_1_2_2(mux_1579_nl, mux_1578_nl, fsm_output(4));
  mux_1584_nl <= MUX_s_1_2_2(mux_1583_nl, mux_1580_nl, fsm_output(6));
  nand_443_nl <= NOT((fsm_output(2)) AND mux_1584_nl);
  or_1759_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (NOT and_763_cse);
  mux_1575_nl <= MUX_s_1_2_2(or_tmp_1645, or_1759_nl, fsm_output(0));
  or_1756_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1574_nl <= MUX_s_1_2_2(or_tmp_1641, or_1756_nl, fsm_output(0));
  mux_1576_nl <= MUX_s_1_2_2(mux_1575_nl, mux_1574_nl, fsm_output(4));
  or_1753_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1572_nl <= MUX_s_1_2_2(or_tmp_1639, or_1753_nl, fsm_output(0));
  or_1750_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1571_nl <= MUX_s_1_2_2(or_tmp_1635, or_1750_nl, fsm_output(0));
  mux_1573_nl <= MUX_s_1_2_2(mux_1572_nl, mux_1571_nl, fsm_output(4));
  mux_1577_nl <= MUX_s_1_2_2(mux_1576_nl, mux_1573_nl, fsm_output(6));
  or_4116_nl <= (fsm_output(2)) OR mux_1577_nl;
  mux_1585_nl <= MUX_s_1_2_2(nand_443_nl, or_4116_nl, fsm_output(5));
  vec_rsc_0_26_i_we_d_pff <= NOT(mux_1585_nl OR (fsm_output(1)));
  or_1792_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1791_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1598_nl <= MUX_s_1_2_2(or_1792_nl, or_1791_nl, fsm_output(0));
  or_1793_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1598_nl;
  or_1789_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011010")) OR (NOT and_763_cse);
  mux_1595_nl <= MUX_s_1_2_2(or_1789_nl, or_tmp_1645, fsm_output(0));
  or_1787_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011010")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1594_nl <= MUX_s_1_2_2(or_1787_nl, or_tmp_1641, fsm_output(0));
  mux_1596_nl <= MUX_s_1_2_2(mux_1595_nl, mux_1594_nl, fsm_output(4));
  or_1786_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011010")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1592_nl <= MUX_s_1_2_2(or_1786_nl, or_tmp_1639, fsm_output(0));
  or_1784_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011010")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1591_nl <= MUX_s_1_2_2(or_1784_nl, or_tmp_1635, fsm_output(0));
  mux_1593_nl <= MUX_s_1_2_2(mux_1592_nl, mux_1591_nl, fsm_output(4));
  mux_1597_nl <= MUX_s_1_2_2(mux_1596_nl, mux_1593_nl, fsm_output(6));
  mux_1599_nl <= MUX_s_1_2_2(or_1793_nl, mux_1597_nl, fsm_output(2));
  or_1782_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1780_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1588_nl <= MUX_s_1_2_2(or_1782_nl, or_1780_nl, fsm_output(0));
  or_1778_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1777_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1587_nl <= MUX_s_1_2_2(or_1778_nl, or_1777_nl, fsm_output(0));
  mux_1589_nl <= MUX_s_1_2_2(mux_1588_nl, mux_1587_nl, fsm_output(4));
  nor_1127_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1128_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1586_nl <= MUX_s_1_2_2(nor_1127_nl, nor_1128_nl, fsm_output(0));
  nand_67_nl <= NOT((fsm_output(4)) AND mux_1586_nl);
  mux_1590_nl <= MUX_s_1_2_2(mux_1589_nl, nand_67_nl, fsm_output(6));
  or_1783_nl <= (fsm_output(2)) OR mux_1590_nl;
  mux_1600_nl <= MUX_s_1_2_2(mux_1599_nl, or_1783_nl, fsm_output(5));
  vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1600_nl) AND (fsm_output(1));
  nor_1118_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(1))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1119_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR not_tmp_330);
  mux_1612_nl <= MUX_s_1_2_2(nor_1118_nl, nor_1119_nl, fsm_output(0));
  nor_1120_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1121_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1611_nl <= MUX_s_1_2_2(nor_1120_nl, nor_1121_nl, fsm_output(0));
  mux_1613_nl <= MUX_s_1_2_2(mux_1612_nl, mux_1611_nl, fsm_output(4));
  nor_1122_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1123_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1609_nl <= MUX_s_1_2_2(nor_1122_nl, nor_1123_nl, fsm_output(0));
  nor_1124_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1125_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1608_nl <= MUX_s_1_2_2(nor_1124_nl, nor_1125_nl, fsm_output(0));
  mux_1610_nl <= MUX_s_1_2_2(mux_1609_nl, mux_1608_nl, fsm_output(4));
  mux_1614_nl <= MUX_s_1_2_2(mux_1613_nl, mux_1610_nl, fsm_output(6));
  nand_442_nl <= NOT((fsm_output(2)) AND mux_1614_nl);
  nand_324_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011011"))
      AND and_763_cse);
  mux_1605_nl <= MUX_s_1_2_2(or_tmp_1689, nand_324_nl, fsm_output(0));
  or_1800_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1604_nl <= MUX_s_1_2_2(or_tmp_1685, or_1800_nl, fsm_output(0));
  mux_1606_nl <= MUX_s_1_2_2(mux_1605_nl, mux_1604_nl, fsm_output(4));
  or_1797_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1602_nl <= MUX_s_1_2_2(or_tmp_1683, or_1797_nl, fsm_output(0));
  or_1794_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1601_nl <= MUX_s_1_2_2(or_tmp_1679, or_1794_nl, fsm_output(0));
  mux_1603_nl <= MUX_s_1_2_2(mux_1602_nl, mux_1601_nl, fsm_output(4));
  mux_1607_nl <= MUX_s_1_2_2(mux_1606_nl, mux_1603_nl, fsm_output(6));
  or_4115_nl <= (fsm_output(2)) OR mux_1607_nl;
  mux_1615_nl <= MUX_s_1_2_2(nand_442_nl, or_4115_nl, fsm_output(5));
  vec_rsc_0_27_i_we_d_pff <= NOT(mux_1615_nl OR (fsm_output(1)));
  or_1836_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1835_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1628_nl <= MUX_s_1_2_2(or_1836_nl, or_1835_nl, fsm_output(0));
  or_1837_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1628_nl;
  nand_323_nl <= NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("011011")) AND and_763_cse);
  mux_1625_nl <= MUX_s_1_2_2(nand_323_nl, or_tmp_1689, fsm_output(0));
  or_1831_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011011")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1624_nl <= MUX_s_1_2_2(or_1831_nl, or_tmp_1685, fsm_output(0));
  mux_1626_nl <= MUX_s_1_2_2(mux_1625_nl, mux_1624_nl, fsm_output(4));
  or_1830_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011011")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1622_nl <= MUX_s_1_2_2(or_1830_nl, or_tmp_1683, fsm_output(0));
  or_1828_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011011")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1621_nl <= MUX_s_1_2_2(or_1828_nl, or_tmp_1679, fsm_output(0));
  mux_1623_nl <= MUX_s_1_2_2(mux_1622_nl, mux_1621_nl, fsm_output(4));
  mux_1627_nl <= MUX_s_1_2_2(mux_1626_nl, mux_1623_nl, fsm_output(6));
  mux_1629_nl <= MUX_s_1_2_2(or_1837_nl, mux_1627_nl, fsm_output(2));
  or_1826_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1824_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1618_nl <= MUX_s_1_2_2(or_1826_nl, or_1824_nl, fsm_output(0));
  or_1822_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1821_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1617_nl <= MUX_s_1_2_2(or_1822_nl, or_1821_nl, fsm_output(0));
  mux_1619_nl <= MUX_s_1_2_2(mux_1618_nl, mux_1617_nl, fsm_output(4));
  nor_1116_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1117_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1616_nl <= MUX_s_1_2_2(nor_1116_nl, nor_1117_nl, fsm_output(0));
  nand_69_nl <= NOT((fsm_output(4)) AND mux_1616_nl);
  mux_1620_nl <= MUX_s_1_2_2(mux_1619_nl, nand_69_nl, fsm_output(6));
  or_1827_nl <= (fsm_output(2)) OR mux_1620_nl;
  mux_1630_nl <= MUX_s_1_2_2(mux_1629_nl, or_1827_nl, fsm_output(5));
  vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1630_nl) AND (fsm_output(1));
  nor_1107_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1108_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_1642_nl <= MUX_s_1_2_2(nor_1107_nl, nor_1108_nl, fsm_output(0));
  nor_1109_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1110_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1641_nl <= MUX_s_1_2_2(nor_1109_nl, nor_1110_nl, fsm_output(0));
  mux_1643_nl <= MUX_s_1_2_2(mux_1642_nl, mux_1641_nl, fsm_output(4));
  nor_1111_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1112_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1639_nl <= MUX_s_1_2_2(nor_1111_nl, nor_1112_nl, fsm_output(0));
  nor_1113_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1114_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1638_nl <= MUX_s_1_2_2(nor_1113_nl, nor_1114_nl, fsm_output(0));
  mux_1640_nl <= MUX_s_1_2_2(mux_1639_nl, mux_1638_nl, fsm_output(4));
  mux_1644_nl <= MUX_s_1_2_2(mux_1643_nl, mux_1640_nl, fsm_output(6));
  nand_441_nl <= NOT((fsm_output(2)) AND mux_1644_nl);
  or_1847_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (NOT and_763_cse);
  mux_1635_nl <= MUX_s_1_2_2(or_tmp_1733, or_1847_nl, fsm_output(0));
  or_1844_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1634_nl <= MUX_s_1_2_2(or_tmp_1729, or_1844_nl, fsm_output(0));
  mux_1636_nl <= MUX_s_1_2_2(mux_1635_nl, mux_1634_nl, fsm_output(4));
  or_1841_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1632_nl <= MUX_s_1_2_2(or_tmp_1727, or_1841_nl, fsm_output(0));
  or_1838_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1631_nl <= MUX_s_1_2_2(or_tmp_1723, or_1838_nl, fsm_output(0));
  mux_1633_nl <= MUX_s_1_2_2(mux_1632_nl, mux_1631_nl, fsm_output(4));
  mux_1637_nl <= MUX_s_1_2_2(mux_1636_nl, mux_1633_nl, fsm_output(6));
  or_4114_nl <= (fsm_output(2)) OR mux_1637_nl;
  mux_1645_nl <= MUX_s_1_2_2(nand_441_nl, or_4114_nl, fsm_output(5));
  vec_rsc_0_28_i_we_d_pff <= NOT(mux_1645_nl OR (fsm_output(1)));
  or_1880_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1879_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1658_nl <= MUX_s_1_2_2(or_1880_nl, or_1879_nl, fsm_output(0));
  or_1881_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1658_nl;
  or_1877_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011100")) OR (NOT and_763_cse);
  mux_1655_nl <= MUX_s_1_2_2(or_1877_nl, or_tmp_1733, fsm_output(0));
  or_1875_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011100")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1654_nl <= MUX_s_1_2_2(or_1875_nl, or_tmp_1729, fsm_output(0));
  mux_1656_nl <= MUX_s_1_2_2(mux_1655_nl, mux_1654_nl, fsm_output(4));
  or_1874_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011100")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1652_nl <= MUX_s_1_2_2(or_1874_nl, or_tmp_1727, fsm_output(0));
  or_1872_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011100")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1651_nl <= MUX_s_1_2_2(or_1872_nl, or_tmp_1723, fsm_output(0));
  mux_1653_nl <= MUX_s_1_2_2(mux_1652_nl, mux_1651_nl, fsm_output(4));
  mux_1657_nl <= MUX_s_1_2_2(mux_1656_nl, mux_1653_nl, fsm_output(6));
  mux_1659_nl <= MUX_s_1_2_2(or_1881_nl, mux_1657_nl, fsm_output(2));
  or_1870_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_1868_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1648_nl <= MUX_s_1_2_2(or_1870_nl, or_1868_nl, fsm_output(0));
  or_1866_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1865_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1647_nl <= MUX_s_1_2_2(or_1866_nl, or_1865_nl, fsm_output(0));
  mux_1649_nl <= MUX_s_1_2_2(mux_1648_nl, mux_1647_nl, fsm_output(4));
  nor_1105_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1106_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1646_nl <= MUX_s_1_2_2(nor_1105_nl, nor_1106_nl, fsm_output(0));
  nand_71_nl <= NOT((fsm_output(4)) AND mux_1646_nl);
  mux_1650_nl <= MUX_s_1_2_2(mux_1649_nl, nand_71_nl, fsm_output(6));
  or_1871_nl <= (fsm_output(2)) OR mux_1650_nl;
  mux_1660_nl <= MUX_s_1_2_2(mux_1659_nl, or_1871_nl, fsm_output(5));
  vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1660_nl) AND (fsm_output(1));
  nor_1096_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  nor_1097_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_1672_nl <= MUX_s_1_2_2(nor_1096_nl, nor_1097_nl, fsm_output(0));
  nor_1098_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1099_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1671_nl <= MUX_s_1_2_2(nor_1098_nl, nor_1099_nl, fsm_output(0));
  mux_1673_nl <= MUX_s_1_2_2(mux_1672_nl, mux_1671_nl, fsm_output(4));
  nor_1100_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1101_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1669_nl <= MUX_s_1_2_2(nor_1100_nl, nor_1101_nl, fsm_output(0));
  nor_1102_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1103_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1668_nl <= MUX_s_1_2_2(nor_1102_nl, nor_1103_nl, fsm_output(0));
  mux_1670_nl <= MUX_s_1_2_2(mux_1669_nl, mux_1668_nl, fsm_output(4));
  mux_1674_nl <= MUX_s_1_2_2(mux_1673_nl, mux_1670_nl, fsm_output(6));
  nand_440_nl <= NOT((fsm_output(2)) AND mux_1674_nl);
  nand_322_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011101"))
      AND and_763_cse);
  mux_1665_nl <= MUX_s_1_2_2(or_tmp_1777, nand_322_nl, fsm_output(0));
  or_1888_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1664_nl <= MUX_s_1_2_2(or_tmp_1773, or_1888_nl, fsm_output(0));
  mux_1666_nl <= MUX_s_1_2_2(mux_1665_nl, mux_1664_nl, fsm_output(4));
  or_1885_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1662_nl <= MUX_s_1_2_2(or_tmp_1771, or_1885_nl, fsm_output(0));
  or_1882_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1661_nl <= MUX_s_1_2_2(or_tmp_1767, or_1882_nl, fsm_output(0));
  mux_1663_nl <= MUX_s_1_2_2(mux_1662_nl, mux_1661_nl, fsm_output(4));
  mux_1667_nl <= MUX_s_1_2_2(mux_1666_nl, mux_1663_nl, fsm_output(6));
  or_4113_nl <= (fsm_output(2)) OR mux_1667_nl;
  mux_1675_nl <= MUX_s_1_2_2(nand_440_nl, or_4113_nl, fsm_output(5));
  vec_rsc_0_29_i_we_d_pff <= NOT(mux_1675_nl OR (fsm_output(1)));
  or_1924_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1923_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1688_nl <= MUX_s_1_2_2(or_1924_nl, or_1923_nl, fsm_output(0));
  or_1925_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1688_nl;
  nand_321_nl <= NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("011101")) AND and_763_cse);
  mux_1685_nl <= MUX_s_1_2_2(nand_321_nl, or_tmp_1777, fsm_output(0));
  or_1919_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011101")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1684_nl <= MUX_s_1_2_2(or_1919_nl, or_tmp_1773, fsm_output(0));
  mux_1686_nl <= MUX_s_1_2_2(mux_1685_nl, mux_1684_nl, fsm_output(4));
  or_1918_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011101")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1682_nl <= MUX_s_1_2_2(or_1918_nl, or_tmp_1771, fsm_output(0));
  or_1916_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011101")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1681_nl <= MUX_s_1_2_2(or_1916_nl, or_tmp_1767, fsm_output(0));
  mux_1683_nl <= MUX_s_1_2_2(mux_1682_nl, mux_1681_nl, fsm_output(4));
  mux_1687_nl <= MUX_s_1_2_2(mux_1686_nl, mux_1683_nl, fsm_output(6));
  mux_1689_nl <= MUX_s_1_2_2(or_1925_nl, mux_1687_nl, fsm_output(2));
  or_1914_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_1912_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(0))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1678_nl <= MUX_s_1_2_2(or_1914_nl, or_1912_nl, fsm_output(0));
  or_1910_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1909_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1677_nl <= MUX_s_1_2_2(or_1910_nl, or_1909_nl, fsm_output(0));
  mux_1679_nl <= MUX_s_1_2_2(mux_1678_nl, mux_1677_nl, fsm_output(4));
  nor_1094_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1095_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1676_nl <= MUX_s_1_2_2(nor_1094_nl, nor_1095_nl, fsm_output(0));
  nand_73_nl <= NOT((fsm_output(4)) AND mux_1676_nl);
  mux_1680_nl <= MUX_s_1_2_2(mux_1679_nl, nand_73_nl, fsm_output(6));
  or_1915_nl <= (fsm_output(2)) OR mux_1680_nl;
  mux_1690_nl <= MUX_s_1_2_2(mux_1689_nl, or_1915_nl, fsm_output(5));
  vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1690_nl) AND (fsm_output(1));
  nor_1086_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(2)))
      OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(1))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) OR not_tmp_384);
  and_602_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND and_763_cse;
  mux_1702_nl <= MUX_s_1_2_2(nor_1086_nl, and_602_nl, fsm_output(0));
  nor_1087_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1088_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1701_nl <= MUX_s_1_2_2(nor_1087_nl, nor_1088_nl, fsm_output(0));
  mux_1703_nl <= MUX_s_1_2_2(mux_1702_nl, mux_1701_nl, fsm_output(4));
  nor_1089_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1090_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1699_nl <= MUX_s_1_2_2(nor_1089_nl, nor_1090_nl, fsm_output(0));
  nor_1091_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1092_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1698_nl <= MUX_s_1_2_2(nor_1091_nl, nor_1092_nl, fsm_output(0));
  mux_1700_nl <= MUX_s_1_2_2(mux_1699_nl, mux_1698_nl, fsm_output(4));
  mux_1704_nl <= MUX_s_1_2_2(mux_1703_nl, mux_1700_nl, fsm_output(6));
  nand_439_nl <= NOT((fsm_output(2)) AND mux_1704_nl);
  nand_320_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011110"))
      AND and_763_cse);
  mux_1695_nl <= MUX_s_1_2_2(or_tmp_1821, nand_320_nl, fsm_output(0));
  or_1932_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1694_nl <= MUX_s_1_2_2(or_tmp_1817, or_1932_nl, fsm_output(0));
  mux_1696_nl <= MUX_s_1_2_2(mux_1695_nl, mux_1694_nl, fsm_output(4));
  or_1929_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1692_nl <= MUX_s_1_2_2(or_tmp_1815, or_1929_nl, fsm_output(0));
  or_1926_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1691_nl <= MUX_s_1_2_2(or_tmp_1811, or_1926_nl, fsm_output(0));
  mux_1693_nl <= MUX_s_1_2_2(mux_1692_nl, mux_1691_nl, fsm_output(4));
  mux_1697_nl <= MUX_s_1_2_2(mux_1696_nl, mux_1693_nl, fsm_output(6));
  or_4112_nl <= (fsm_output(2)) OR mux_1697_nl;
  mux_1705_nl <= MUX_s_1_2_2(nand_439_nl, or_4112_nl, fsm_output(5));
  vec_rsc_0_30_i_we_d_pff <= NOT(mux_1705_nl OR (fsm_output(1)));
  or_1968_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_1967_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1718_nl <= MUX_s_1_2_2(or_1968_nl, or_1967_nl, fsm_output(0));
  or_1969_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1718_nl;
  nand_318_nl <= NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("011110")) AND and_763_cse);
  mux_1715_nl <= MUX_s_1_2_2(nand_318_nl, or_tmp_1821, fsm_output(0));
  or_1963_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011110")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1714_nl <= MUX_s_1_2_2(or_1963_nl, or_tmp_1817, fsm_output(0));
  mux_1716_nl <= MUX_s_1_2_2(mux_1715_nl, mux_1714_nl, fsm_output(4));
  or_1962_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011110")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1712_nl <= MUX_s_1_2_2(or_1962_nl, or_tmp_1815, fsm_output(0));
  or_1960_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011110")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1711_nl <= MUX_s_1_2_2(or_1960_nl, or_tmp_1811, fsm_output(0));
  mux_1713_nl <= MUX_s_1_2_2(mux_1712_nl, mux_1711_nl, fsm_output(4));
  mux_1717_nl <= MUX_s_1_2_2(mux_1716_nl, mux_1713_nl, fsm_output(6));
  mux_1719_nl <= MUX_s_1_2_2(or_1969_nl, mux_1717_nl, fsm_output(2));
  nand_319_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND and_763_cse);
  or_1956_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(2)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) OR not_tmp_388;
  mux_1708_nl <= MUX_s_1_2_2(nand_319_nl, or_1956_nl, fsm_output(0));
  or_1954_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_1953_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1707_nl <= MUX_s_1_2_2(or_1954_nl, or_1953_nl, fsm_output(0));
  mux_1709_nl <= MUX_s_1_2_2(mux_1708_nl, mux_1707_nl, fsm_output(4));
  nor_1084_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1085_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1706_nl <= MUX_s_1_2_2(nor_1084_nl, nor_1085_nl, fsm_output(0));
  nand_75_nl <= NOT((fsm_output(4)) AND mux_1706_nl);
  mux_1710_nl <= MUX_s_1_2_2(mux_1709_nl, nand_75_nl, fsm_output(6));
  or_1959_nl <= (fsm_output(2)) OR mux_1710_nl;
  mux_1720_nl <= MUX_s_1_2_2(mux_1719_nl, or_1959_nl, fsm_output(5));
  vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1720_nl) AND (fsm_output(1));
  nor_1077_nl <= NOT((NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      AND (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      AND (NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(5))))) OR not_tmp_384);
  nor_1078_nl <= NOT((COMP_LOOP_acc_13_psp_sva(3)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(3)) AND (fsm_output(7)))));
  mux_1732_nl <= MUX_s_1_2_2(nor_1077_nl, nor_1078_nl, fsm_output(0));
  and_599_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_600_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  mux_1731_nl <= MUX_s_1_2_2(and_599_nl, and_600_nl, fsm_output(0));
  mux_1733_nl <= MUX_s_1_2_2(mux_1732_nl, mux_1731_nl, fsm_output(4));
  and_811_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7));
  and_818_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT (fsm_output(3))) AND (fsm_output(7));
  mux_1729_nl <= MUX_s_1_2_2(and_811_nl, and_818_nl, fsm_output(0));
  nor_1081_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1082_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1728_nl <= MUX_s_1_2_2(nor_1081_nl, nor_1082_nl, fsm_output(0));
  mux_1730_nl <= MUX_s_1_2_2(mux_1729_nl, mux_1728_nl, fsm_output(4));
  mux_1734_nl <= MUX_s_1_2_2(mux_1733_nl, mux_1730_nl, fsm_output(6));
  nand_438_nl <= NOT((fsm_output(2)) AND mux_1734_nl);
  nand_313_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND and_763_cse);
  mux_1725_nl <= MUX_s_1_2_2(or_tmp_1865, nand_313_nl, fsm_output(0));
  nand_314_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_1724_nl <= MUX_s_1_2_2(or_tmp_1861, nand_314_nl, fsm_output(0));
  mux_1726_nl <= MUX_s_1_2_2(mux_1725_nl, mux_1724_nl, fsm_output(4));
  nand_478_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_1722_nl <= MUX_s_1_2_2(or_tmp_1859, nand_478_nl, fsm_output(0));
  or_1970_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1721_nl <= MUX_s_1_2_2(or_tmp_1855, or_1970_nl, fsm_output(0));
  mux_1723_nl <= MUX_s_1_2_2(mux_1722_nl, mux_1721_nl, fsm_output(4));
  mux_1727_nl <= MUX_s_1_2_2(mux_1726_nl, mux_1723_nl, fsm_output(6));
  or_4111_nl <= (fsm_output(2)) OR mux_1727_nl;
  mux_1735_nl <= MUX_s_1_2_2(nand_438_nl, or_4111_nl, fsm_output(5));
  vec_rsc_0_31_i_we_d_pff <= NOT(mux_1735_nl OR (fsm_output(1)));
  or_2011_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2010_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1748_nl <= MUX_s_1_2_2(or_2011_nl, or_2010_nl, fsm_output(0));
  or_2012_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1748_nl;
  nand_302_nl <= NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("011111")) AND and_763_cse);
  mux_1745_nl <= MUX_s_1_2_2(nand_302_nl, or_tmp_1865, fsm_output(0));
  nand_303_nl <= NOT(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("011111")) AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_1744_nl <= MUX_s_1_2_2(nand_303_nl, or_tmp_1861, fsm_output(0));
  mux_1746_nl <= MUX_s_1_2_2(mux_1745_nl, mux_1744_nl, fsm_output(4));
  nand_404_nl <= NOT(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("011111")) AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_1742_nl <= MUX_s_1_2_2(nand_404_nl, or_tmp_1859, fsm_output(0));
  or_2003_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011111")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1741_nl <= MUX_s_1_2_2(or_2003_nl, or_tmp_1855, fsm_output(0));
  mux_1743_nl <= MUX_s_1_2_2(mux_1742_nl, mux_1741_nl, fsm_output(4));
  mux_1747_nl <= MUX_s_1_2_2(mux_1746_nl, mux_1743_nl, fsm_output(6));
  mux_1749_nl <= MUX_s_1_2_2(or_2012_nl, mux_1747_nl, fsm_output(2));
  or_2001_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)) OR not_tmp_321;
  or_1999_nl <= (NOT((COMP_LOOP_acc_10_cse_10_1_7_sva(1)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      AND (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      AND (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(5))))) OR not_tmp_388;
  mux_1738_nl <= MUX_s_1_2_2(or_2001_nl, or_1999_nl, fsm_output(0));
  nand_307_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))
      AND COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
      (fsm_output(3)) AND (NOT (fsm_output(7))));
  nand_308_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_1737_nl <= MUX_s_1_2_2(nand_307_nl, nand_308_nl, fsm_output(0));
  mux_1739_nl <= MUX_s_1_2_2(mux_1738_nl, mux_1737_nl, fsm_output(4));
  nor_1075_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1076_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1736_nl <= MUX_s_1_2_2(nor_1075_nl, nor_1076_nl, fsm_output(0));
  nand_77_nl <= NOT((fsm_output(4)) AND mux_1736_nl);
  mux_1740_nl <= MUX_s_1_2_2(mux_1739_nl, nand_77_nl, fsm_output(6));
  or_2002_nl <= (fsm_output(2)) OR mux_1740_nl;
  mux_1750_nl <= MUX_s_1_2_2(mux_1749_nl, or_2002_nl, fsm_output(5));
  vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1750_nl) AND (fsm_output(1));
  nor_1066_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (NOT and_763_cse));
  nor_1067_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_1762_nl <= MUX_s_1_2_2(nor_1066_nl, nor_1067_nl, fsm_output(0));
  nor_1068_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1069_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1761_nl <= MUX_s_1_2_2(nor_1068_nl, nor_1069_nl, fsm_output(0));
  mux_1763_nl <= MUX_s_1_2_2(mux_1762_nl, mux_1761_nl, fsm_output(4));
  nor_1070_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1071_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1759_nl <= MUX_s_1_2_2(nor_1070_nl, nor_1071_nl, fsm_output(0));
  nor_1072_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1073_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1758_nl <= MUX_s_1_2_2(nor_1072_nl, nor_1073_nl, fsm_output(0));
  mux_1760_nl <= MUX_s_1_2_2(mux_1759_nl, mux_1758_nl, fsm_output(4));
  mux_1764_nl <= MUX_s_1_2_2(mux_1763_nl, mux_1760_nl, fsm_output(6));
  nand_437_nl <= NOT((fsm_output(2)) AND mux_1764_nl);
  or_2022_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR not_tmp_452;
  mux_1755_nl <= MUX_s_1_2_2(or_tmp_1908, or_2022_nl, fsm_output(0));
  or_2019_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1754_nl <= MUX_s_1_2_2(or_tmp_1904, or_2019_nl, fsm_output(0));
  mux_1756_nl <= MUX_s_1_2_2(mux_1755_nl, mux_1754_nl, fsm_output(4));
  or_2016_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1752_nl <= MUX_s_1_2_2(or_tmp_1902, or_2016_nl, fsm_output(0));
  or_2013_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1751_nl <= MUX_s_1_2_2(or_tmp_1898, or_2013_nl, fsm_output(0));
  mux_1753_nl <= MUX_s_1_2_2(mux_1752_nl, mux_1751_nl, fsm_output(4));
  mux_1757_nl <= MUX_s_1_2_2(mux_1756_nl, mux_1753_nl, fsm_output(6));
  or_4110_nl <= (fsm_output(2)) OR mux_1757_nl;
  mux_1765_nl <= MUX_s_1_2_2(nand_437_nl, or_4110_nl, fsm_output(5));
  vec_rsc_0_32_i_we_d_pff <= NOT(mux_1765_nl OR (fsm_output(1)));
  or_2055_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2054_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1778_nl <= MUX_s_1_2_2(or_2055_nl, or_2054_nl, fsm_output(0));
  or_2056_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1778_nl;
  or_2052_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")) OR not_tmp_452;
  mux_1775_nl <= MUX_s_1_2_2(or_2052_nl, or_tmp_1908, fsm_output(0));
  or_2050_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100000")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1774_nl <= MUX_s_1_2_2(or_2050_nl, or_tmp_1904, fsm_output(0));
  mux_1776_nl <= MUX_s_1_2_2(mux_1775_nl, mux_1774_nl, fsm_output(4));
  or_2049_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100000")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1772_nl <= MUX_s_1_2_2(or_2049_nl, or_tmp_1902, fsm_output(0));
  or_2047_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100000")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1771_nl <= MUX_s_1_2_2(or_2047_nl, or_tmp_1898, fsm_output(0));
  mux_1773_nl <= MUX_s_1_2_2(mux_1772_nl, mux_1771_nl, fsm_output(4));
  mux_1777_nl <= MUX_s_1_2_2(mux_1776_nl, mux_1773_nl, fsm_output(6));
  mux_1779_nl <= MUX_s_1_2_2(or_2056_nl, mux_1777_nl, fsm_output(2));
  or_2045_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2043_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (NOT and_763_cse);
  mux_1768_nl <= MUX_s_1_2_2(or_2045_nl, or_2043_nl, fsm_output(0));
  or_2041_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2040_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1767_nl <= MUX_s_1_2_2(or_2041_nl, or_2040_nl, fsm_output(0));
  mux_1769_nl <= MUX_s_1_2_2(mux_1768_nl, mux_1767_nl, fsm_output(4));
  nor_1064_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1065_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1766_nl <= MUX_s_1_2_2(nor_1064_nl, nor_1065_nl, fsm_output(0));
  nand_79_nl <= NOT((fsm_output(4)) AND mux_1766_nl);
  mux_1770_nl <= MUX_s_1_2_2(mux_1769_nl, nand_79_nl, fsm_output(6));
  or_2046_nl <= (fsm_output(2)) OR mux_1770_nl;
  mux_1780_nl <= MUX_s_1_2_2(mux_1779_nl, or_2046_nl, fsm_output(5));
  vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1780_nl) AND (fsm_output(1));
  nor_1055_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (NOT and_763_cse));
  nor_1056_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_1792_nl <= MUX_s_1_2_2(nor_1055_nl, nor_1056_nl, fsm_output(0));
  nor_1057_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1058_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1791_nl <= MUX_s_1_2_2(nor_1057_nl, nor_1058_nl, fsm_output(0));
  mux_1793_nl <= MUX_s_1_2_2(mux_1792_nl, mux_1791_nl, fsm_output(4));
  nor_1059_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1060_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1789_nl <= MUX_s_1_2_2(nor_1059_nl, nor_1060_nl, fsm_output(0));
  nor_1061_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1062_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1788_nl <= MUX_s_1_2_2(nor_1061_nl, nor_1062_nl, fsm_output(0));
  mux_1790_nl <= MUX_s_1_2_2(mux_1789_nl, mux_1788_nl, fsm_output(4));
  mux_1794_nl <= MUX_s_1_2_2(mux_1793_nl, mux_1790_nl, fsm_output(6));
  nand_436_nl <= NOT((fsm_output(2)) AND mux_1794_nl);
  or_2066_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR not_tmp_452;
  mux_1785_nl <= MUX_s_1_2_2(or_tmp_1952, or_2066_nl, fsm_output(0));
  or_2063_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1784_nl <= MUX_s_1_2_2(or_tmp_1948, or_2063_nl, fsm_output(0));
  mux_1786_nl <= MUX_s_1_2_2(mux_1785_nl, mux_1784_nl, fsm_output(4));
  or_2060_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1782_nl <= MUX_s_1_2_2(or_tmp_1946, or_2060_nl, fsm_output(0));
  or_2057_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1781_nl <= MUX_s_1_2_2(or_tmp_1942, or_2057_nl, fsm_output(0));
  mux_1783_nl <= MUX_s_1_2_2(mux_1782_nl, mux_1781_nl, fsm_output(4));
  mux_1787_nl <= MUX_s_1_2_2(mux_1786_nl, mux_1783_nl, fsm_output(6));
  or_4109_nl <= (fsm_output(2)) OR mux_1787_nl;
  mux_1795_nl <= MUX_s_1_2_2(nand_436_nl, or_4109_nl, fsm_output(5));
  vec_rsc_0_33_i_we_d_pff <= NOT(mux_1795_nl OR (fsm_output(1)));
  or_2099_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2098_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1808_nl <= MUX_s_1_2_2(or_2099_nl, or_2098_nl, fsm_output(0));
  or_2100_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1808_nl;
  or_2096_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00001")) OR not_tmp_452;
  mux_1805_nl <= MUX_s_1_2_2(or_2096_nl, or_tmp_1952, fsm_output(0));
  or_2094_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100001")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1804_nl <= MUX_s_1_2_2(or_2094_nl, or_tmp_1948, fsm_output(0));
  mux_1806_nl <= MUX_s_1_2_2(mux_1805_nl, mux_1804_nl, fsm_output(4));
  or_2093_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100001")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1802_nl <= MUX_s_1_2_2(or_2093_nl, or_tmp_1946, fsm_output(0));
  or_2091_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100001")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1801_nl <= MUX_s_1_2_2(or_2091_nl, or_tmp_1942, fsm_output(0));
  mux_1803_nl <= MUX_s_1_2_2(mux_1802_nl, mux_1801_nl, fsm_output(4));
  mux_1807_nl <= MUX_s_1_2_2(mux_1806_nl, mux_1803_nl, fsm_output(6));
  mux_1809_nl <= MUX_s_1_2_2(or_2100_nl, mux_1807_nl, fsm_output(2));
  or_2089_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_2087_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (NOT and_763_cse);
  mux_1798_nl <= MUX_s_1_2_2(or_2089_nl, or_2087_nl, fsm_output(0));
  or_2085_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2084_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1797_nl <= MUX_s_1_2_2(or_2085_nl, or_2084_nl, fsm_output(0));
  mux_1799_nl <= MUX_s_1_2_2(mux_1798_nl, mux_1797_nl, fsm_output(4));
  nor_1053_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1054_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1796_nl <= MUX_s_1_2_2(nor_1053_nl, nor_1054_nl, fsm_output(0));
  nand_81_nl <= NOT((fsm_output(4)) AND mux_1796_nl);
  mux_1800_nl <= MUX_s_1_2_2(mux_1799_nl, nand_81_nl, fsm_output(6));
  or_2090_nl <= (fsm_output(2)) OR mux_1800_nl;
  mux_1810_nl <= MUX_s_1_2_2(mux_1809_nl, or_2090_nl, fsm_output(5));
  vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1810_nl) AND (fsm_output(1));
  nor_1044_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (NOT and_763_cse));
  nor_1045_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_1822_nl <= MUX_s_1_2_2(nor_1044_nl, nor_1045_nl, fsm_output(0));
  nor_1046_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1047_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1821_nl <= MUX_s_1_2_2(nor_1046_nl, nor_1047_nl, fsm_output(0));
  mux_1823_nl <= MUX_s_1_2_2(mux_1822_nl, mux_1821_nl, fsm_output(4));
  nor_1048_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1049_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1819_nl <= MUX_s_1_2_2(nor_1048_nl, nor_1049_nl, fsm_output(0));
  nor_1050_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1051_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1818_nl <= MUX_s_1_2_2(nor_1050_nl, nor_1051_nl, fsm_output(0));
  mux_1820_nl <= MUX_s_1_2_2(mux_1819_nl, mux_1818_nl, fsm_output(4));
  mux_1824_nl <= MUX_s_1_2_2(mux_1823_nl, mux_1820_nl, fsm_output(6));
  nand_435_nl <= NOT((fsm_output(2)) AND mux_1824_nl);
  or_2110_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR not_tmp_452;
  mux_1815_nl <= MUX_s_1_2_2(or_tmp_1996, or_2110_nl, fsm_output(0));
  or_2107_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1814_nl <= MUX_s_1_2_2(or_tmp_1992, or_2107_nl, fsm_output(0));
  mux_1816_nl <= MUX_s_1_2_2(mux_1815_nl, mux_1814_nl, fsm_output(4));
  or_2104_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1812_nl <= MUX_s_1_2_2(or_tmp_1990, or_2104_nl, fsm_output(0));
  or_2101_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1811_nl <= MUX_s_1_2_2(or_tmp_1986, or_2101_nl, fsm_output(0));
  mux_1813_nl <= MUX_s_1_2_2(mux_1812_nl, mux_1811_nl, fsm_output(4));
  mux_1817_nl <= MUX_s_1_2_2(mux_1816_nl, mux_1813_nl, fsm_output(6));
  or_4108_nl <= (fsm_output(2)) OR mux_1817_nl;
  mux_1825_nl <= MUX_s_1_2_2(nand_435_nl, or_4108_nl, fsm_output(5));
  vec_rsc_0_34_i_we_d_pff <= NOT(mux_1825_nl OR (fsm_output(1)));
  or_2143_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2142_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1838_nl <= MUX_s_1_2_2(or_2143_nl, or_2142_nl, fsm_output(0));
  or_2144_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1838_nl;
  or_2140_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00010")) OR not_tmp_452;
  mux_1835_nl <= MUX_s_1_2_2(or_2140_nl, or_tmp_1996, fsm_output(0));
  or_2138_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100010")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1834_nl <= MUX_s_1_2_2(or_2138_nl, or_tmp_1992, fsm_output(0));
  mux_1836_nl <= MUX_s_1_2_2(mux_1835_nl, mux_1834_nl, fsm_output(4));
  or_2137_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100010")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1832_nl <= MUX_s_1_2_2(or_2137_nl, or_tmp_1990, fsm_output(0));
  or_2135_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100010")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1831_nl <= MUX_s_1_2_2(or_2135_nl, or_tmp_1986, fsm_output(0));
  mux_1833_nl <= MUX_s_1_2_2(mux_1832_nl, mux_1831_nl, fsm_output(4));
  mux_1837_nl <= MUX_s_1_2_2(mux_1836_nl, mux_1833_nl, fsm_output(6));
  mux_1839_nl <= MUX_s_1_2_2(or_2144_nl, mux_1837_nl, fsm_output(2));
  or_2133_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2131_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (NOT and_763_cse);
  mux_1828_nl <= MUX_s_1_2_2(or_2133_nl, or_2131_nl, fsm_output(0));
  or_2129_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2128_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1827_nl <= MUX_s_1_2_2(or_2129_nl, or_2128_nl, fsm_output(0));
  mux_1829_nl <= MUX_s_1_2_2(mux_1828_nl, mux_1827_nl, fsm_output(4));
  nor_1042_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1043_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1826_nl <= MUX_s_1_2_2(nor_1042_nl, nor_1043_nl, fsm_output(0));
  nand_83_nl <= NOT((fsm_output(4)) AND mux_1826_nl);
  mux_1830_nl <= MUX_s_1_2_2(mux_1829_nl, nand_83_nl, fsm_output(6));
  or_2134_nl <= (fsm_output(2)) OR mux_1830_nl;
  mux_1840_nl <= MUX_s_1_2_2(mux_1839_nl, or_2134_nl, fsm_output(5));
  vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1840_nl) AND (fsm_output(1));
  nor_1033_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (NOT and_763_cse));
  nor_1034_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR not_tmp_330);
  mux_1852_nl <= MUX_s_1_2_2(nor_1033_nl, nor_1034_nl, fsm_output(0));
  nor_1035_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1036_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1851_nl <= MUX_s_1_2_2(nor_1035_nl, nor_1036_nl, fsm_output(0));
  mux_1853_nl <= MUX_s_1_2_2(mux_1852_nl, mux_1851_nl, fsm_output(4));
  nor_1037_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1038_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1849_nl <= MUX_s_1_2_2(nor_1037_nl, nor_1038_nl, fsm_output(0));
  nor_1039_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1040_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1848_nl <= MUX_s_1_2_2(nor_1039_nl, nor_1040_nl, fsm_output(0));
  mux_1850_nl <= MUX_s_1_2_2(mux_1849_nl, mux_1848_nl, fsm_output(4));
  mux_1854_nl <= MUX_s_1_2_2(mux_1853_nl, mux_1850_nl, fsm_output(6));
  nand_434_nl <= NOT((fsm_output(2)) AND mux_1854_nl);
  or_2154_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR not_tmp_452;
  mux_1845_nl <= MUX_s_1_2_2(or_tmp_2040, or_2154_nl, fsm_output(0));
  or_2151_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1844_nl <= MUX_s_1_2_2(or_tmp_2036, or_2151_nl, fsm_output(0));
  mux_1846_nl <= MUX_s_1_2_2(mux_1845_nl, mux_1844_nl, fsm_output(4));
  or_2148_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1842_nl <= MUX_s_1_2_2(or_tmp_2034, or_2148_nl, fsm_output(0));
  or_2145_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1841_nl <= MUX_s_1_2_2(or_tmp_2030, or_2145_nl, fsm_output(0));
  mux_1843_nl <= MUX_s_1_2_2(mux_1842_nl, mux_1841_nl, fsm_output(4));
  mux_1847_nl <= MUX_s_1_2_2(mux_1846_nl, mux_1843_nl, fsm_output(6));
  or_4107_nl <= (fsm_output(2)) OR mux_1847_nl;
  mux_1855_nl <= MUX_s_1_2_2(nand_434_nl, or_4107_nl, fsm_output(5));
  vec_rsc_0_35_i_we_d_pff <= NOT(mux_1855_nl OR (fsm_output(1)));
  or_2187_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2186_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1868_nl <= MUX_s_1_2_2(or_2187_nl, or_2186_nl, fsm_output(0));
  or_2188_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1868_nl;
  or_2184_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00011")) OR not_tmp_452;
  mux_1865_nl <= MUX_s_1_2_2(or_2184_nl, or_tmp_2040, fsm_output(0));
  or_2182_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100011")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1864_nl <= MUX_s_1_2_2(or_2182_nl, or_tmp_2036, fsm_output(0));
  mux_1866_nl <= MUX_s_1_2_2(mux_1865_nl, mux_1864_nl, fsm_output(4));
  or_2181_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100011")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1862_nl <= MUX_s_1_2_2(or_2181_nl, or_tmp_2034, fsm_output(0));
  or_2179_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100011")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1861_nl <= MUX_s_1_2_2(or_2179_nl, or_tmp_2030, fsm_output(0));
  mux_1863_nl <= MUX_s_1_2_2(mux_1862_nl, mux_1861_nl, fsm_output(4));
  mux_1867_nl <= MUX_s_1_2_2(mux_1866_nl, mux_1863_nl, fsm_output(6));
  mux_1869_nl <= MUX_s_1_2_2(or_2188_nl, mux_1867_nl, fsm_output(2));
  or_2177_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_2175_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (NOT and_763_cse);
  mux_1858_nl <= MUX_s_1_2_2(or_2177_nl, or_2175_nl, fsm_output(0));
  or_2173_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2172_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1857_nl <= MUX_s_1_2_2(or_2173_nl, or_2172_nl, fsm_output(0));
  mux_1859_nl <= MUX_s_1_2_2(mux_1858_nl, mux_1857_nl, fsm_output(4));
  nor_1031_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1032_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1856_nl <= MUX_s_1_2_2(nor_1031_nl, nor_1032_nl, fsm_output(0));
  nand_85_nl <= NOT((fsm_output(4)) AND mux_1856_nl);
  mux_1860_nl <= MUX_s_1_2_2(mux_1859_nl, nand_85_nl, fsm_output(6));
  or_2178_nl <= (fsm_output(2)) OR mux_1860_nl;
  mux_1870_nl <= MUX_s_1_2_2(mux_1869_nl, or_2178_nl, fsm_output(5));
  vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1870_nl) AND (fsm_output(1));
  nor_1022_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (NOT and_763_cse));
  nor_1023_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_1882_nl <= MUX_s_1_2_2(nor_1022_nl, nor_1023_nl, fsm_output(0));
  nor_1024_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1025_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1881_nl <= MUX_s_1_2_2(nor_1024_nl, nor_1025_nl, fsm_output(0));
  mux_1883_nl <= MUX_s_1_2_2(mux_1882_nl, mux_1881_nl, fsm_output(4));
  nor_1026_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1027_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1879_nl <= MUX_s_1_2_2(nor_1026_nl, nor_1027_nl, fsm_output(0));
  nor_1028_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1029_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1878_nl <= MUX_s_1_2_2(nor_1028_nl, nor_1029_nl, fsm_output(0));
  mux_1880_nl <= MUX_s_1_2_2(mux_1879_nl, mux_1878_nl, fsm_output(4));
  mux_1884_nl <= MUX_s_1_2_2(mux_1883_nl, mux_1880_nl, fsm_output(6));
  nand_433_nl <= NOT((fsm_output(2)) AND mux_1884_nl);
  or_2198_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR not_tmp_452;
  mux_1875_nl <= MUX_s_1_2_2(or_tmp_2084, or_2198_nl, fsm_output(0));
  or_2195_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1874_nl <= MUX_s_1_2_2(or_tmp_2080, or_2195_nl, fsm_output(0));
  mux_1876_nl <= MUX_s_1_2_2(mux_1875_nl, mux_1874_nl, fsm_output(4));
  or_2192_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1872_nl <= MUX_s_1_2_2(or_tmp_2078, or_2192_nl, fsm_output(0));
  or_2189_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1871_nl <= MUX_s_1_2_2(or_tmp_2074, or_2189_nl, fsm_output(0));
  mux_1873_nl <= MUX_s_1_2_2(mux_1872_nl, mux_1871_nl, fsm_output(4));
  mux_1877_nl <= MUX_s_1_2_2(mux_1876_nl, mux_1873_nl, fsm_output(6));
  or_4106_nl <= (fsm_output(2)) OR mux_1877_nl;
  mux_1885_nl <= MUX_s_1_2_2(nand_433_nl, or_4106_nl, fsm_output(5));
  vec_rsc_0_36_i_we_d_pff <= NOT(mux_1885_nl OR (fsm_output(1)));
  or_2231_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2230_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1898_nl <= MUX_s_1_2_2(or_2231_nl, or_2230_nl, fsm_output(0));
  or_2232_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1898_nl;
  or_2228_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00100")) OR not_tmp_452;
  mux_1895_nl <= MUX_s_1_2_2(or_2228_nl, or_tmp_2084, fsm_output(0));
  or_2226_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100100")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1894_nl <= MUX_s_1_2_2(or_2226_nl, or_tmp_2080, fsm_output(0));
  mux_1896_nl <= MUX_s_1_2_2(mux_1895_nl, mux_1894_nl, fsm_output(4));
  or_2225_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100100")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1892_nl <= MUX_s_1_2_2(or_2225_nl, or_tmp_2078, fsm_output(0));
  or_2223_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100100")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1891_nl <= MUX_s_1_2_2(or_2223_nl, or_tmp_2074, fsm_output(0));
  mux_1893_nl <= MUX_s_1_2_2(mux_1892_nl, mux_1891_nl, fsm_output(4));
  mux_1897_nl <= MUX_s_1_2_2(mux_1896_nl, mux_1893_nl, fsm_output(6));
  mux_1899_nl <= MUX_s_1_2_2(or_2232_nl, mux_1897_nl, fsm_output(2));
  or_2221_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2219_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (NOT and_763_cse);
  mux_1888_nl <= MUX_s_1_2_2(or_2221_nl, or_2219_nl, fsm_output(0));
  or_2217_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2216_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1887_nl <= MUX_s_1_2_2(or_2217_nl, or_2216_nl, fsm_output(0));
  mux_1889_nl <= MUX_s_1_2_2(mux_1888_nl, mux_1887_nl, fsm_output(4));
  nor_1020_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1021_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1886_nl <= MUX_s_1_2_2(nor_1020_nl, nor_1021_nl, fsm_output(0));
  nand_87_nl <= NOT((fsm_output(4)) AND mux_1886_nl);
  mux_1890_nl <= MUX_s_1_2_2(mux_1889_nl, nand_87_nl, fsm_output(6));
  or_2222_nl <= (fsm_output(2)) OR mux_1890_nl;
  mux_1900_nl <= MUX_s_1_2_2(mux_1899_nl, or_2222_nl, fsm_output(5));
  vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1900_nl) AND (fsm_output(1));
  nor_1011_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (NOT and_763_cse));
  nor_1012_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_1912_nl <= MUX_s_1_2_2(nor_1011_nl, nor_1012_nl, fsm_output(0));
  nor_1013_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1014_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1911_nl <= MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, fsm_output(0));
  mux_1913_nl <= MUX_s_1_2_2(mux_1912_nl, mux_1911_nl, fsm_output(4));
  nor_1015_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1016_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1909_nl <= MUX_s_1_2_2(nor_1015_nl, nor_1016_nl, fsm_output(0));
  nor_1017_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1018_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1908_nl <= MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, fsm_output(0));
  mux_1910_nl <= MUX_s_1_2_2(mux_1909_nl, mux_1908_nl, fsm_output(4));
  mux_1914_nl <= MUX_s_1_2_2(mux_1913_nl, mux_1910_nl, fsm_output(6));
  nand_432_nl <= NOT((fsm_output(2)) AND mux_1914_nl);
  or_2242_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR not_tmp_452;
  mux_1905_nl <= MUX_s_1_2_2(or_tmp_2128, or_2242_nl, fsm_output(0));
  or_2239_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1904_nl <= MUX_s_1_2_2(or_tmp_2124, or_2239_nl, fsm_output(0));
  mux_1906_nl <= MUX_s_1_2_2(mux_1905_nl, mux_1904_nl, fsm_output(4));
  or_2236_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1902_nl <= MUX_s_1_2_2(or_tmp_2122, or_2236_nl, fsm_output(0));
  or_2233_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1901_nl <= MUX_s_1_2_2(or_tmp_2118, or_2233_nl, fsm_output(0));
  mux_1903_nl <= MUX_s_1_2_2(mux_1902_nl, mux_1901_nl, fsm_output(4));
  mux_1907_nl <= MUX_s_1_2_2(mux_1906_nl, mux_1903_nl, fsm_output(6));
  or_4105_nl <= (fsm_output(2)) OR mux_1907_nl;
  mux_1915_nl <= MUX_s_1_2_2(nand_432_nl, or_4105_nl, fsm_output(5));
  vec_rsc_0_37_i_we_d_pff <= NOT(mux_1915_nl OR (fsm_output(1)));
  or_2275_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2274_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1928_nl <= MUX_s_1_2_2(or_2275_nl, or_2274_nl, fsm_output(0));
  or_2276_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1928_nl;
  or_2272_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00101")) OR not_tmp_452;
  mux_1925_nl <= MUX_s_1_2_2(or_2272_nl, or_tmp_2128, fsm_output(0));
  or_2270_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100101")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1924_nl <= MUX_s_1_2_2(or_2270_nl, or_tmp_2124, fsm_output(0));
  mux_1926_nl <= MUX_s_1_2_2(mux_1925_nl, mux_1924_nl, fsm_output(4));
  or_2269_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100101")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1922_nl <= MUX_s_1_2_2(or_2269_nl, or_tmp_2122, fsm_output(0));
  or_2267_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100101")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1921_nl <= MUX_s_1_2_2(or_2267_nl, or_tmp_2118, fsm_output(0));
  mux_1923_nl <= MUX_s_1_2_2(mux_1922_nl, mux_1921_nl, fsm_output(4));
  mux_1927_nl <= MUX_s_1_2_2(mux_1926_nl, mux_1923_nl, fsm_output(6));
  mux_1929_nl <= MUX_s_1_2_2(or_2276_nl, mux_1927_nl, fsm_output(2));
  or_2265_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_2263_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (NOT and_763_cse);
  mux_1918_nl <= MUX_s_1_2_2(or_2265_nl, or_2263_nl, fsm_output(0));
  or_2261_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2260_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1917_nl <= MUX_s_1_2_2(or_2261_nl, or_2260_nl, fsm_output(0));
  mux_1919_nl <= MUX_s_1_2_2(mux_1918_nl, mux_1917_nl, fsm_output(4));
  nor_1009_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1010_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1916_nl <= MUX_s_1_2_2(nor_1009_nl, nor_1010_nl, fsm_output(0));
  nand_89_nl <= NOT((fsm_output(4)) AND mux_1916_nl);
  mux_1920_nl <= MUX_s_1_2_2(mux_1919_nl, nand_89_nl, fsm_output(6));
  or_2266_nl <= (fsm_output(2)) OR mux_1920_nl;
  mux_1930_nl <= MUX_s_1_2_2(mux_1929_nl, or_2266_nl, fsm_output(5));
  vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1930_nl) AND (fsm_output(1));
  nor_1000_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (NOT and_763_cse));
  nor_1001_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_1942_nl <= MUX_s_1_2_2(nor_1000_nl, nor_1001_nl, fsm_output(0));
  nor_1002_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_1003_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1941_nl <= MUX_s_1_2_2(nor_1002_nl, nor_1003_nl, fsm_output(0));
  mux_1943_nl <= MUX_s_1_2_2(mux_1942_nl, mux_1941_nl, fsm_output(4));
  nor_1004_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_1005_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1939_nl <= MUX_s_1_2_2(nor_1004_nl, nor_1005_nl, fsm_output(0));
  nor_1006_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1007_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1938_nl <= MUX_s_1_2_2(nor_1006_nl, nor_1007_nl, fsm_output(0));
  mux_1940_nl <= MUX_s_1_2_2(mux_1939_nl, mux_1938_nl, fsm_output(4));
  mux_1944_nl <= MUX_s_1_2_2(mux_1943_nl, mux_1940_nl, fsm_output(6));
  nand_431_nl <= NOT((fsm_output(2)) AND mux_1944_nl);
  or_2286_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR not_tmp_452;
  mux_1935_nl <= MUX_s_1_2_2(or_tmp_2172, or_2286_nl, fsm_output(0));
  or_2283_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1934_nl <= MUX_s_1_2_2(or_tmp_2168, or_2283_nl, fsm_output(0));
  mux_1936_nl <= MUX_s_1_2_2(mux_1935_nl, mux_1934_nl, fsm_output(4));
  or_2280_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1932_nl <= MUX_s_1_2_2(or_tmp_2166, or_2280_nl, fsm_output(0));
  or_2277_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1931_nl <= MUX_s_1_2_2(or_tmp_2162, or_2277_nl, fsm_output(0));
  mux_1933_nl <= MUX_s_1_2_2(mux_1932_nl, mux_1931_nl, fsm_output(4));
  mux_1937_nl <= MUX_s_1_2_2(mux_1936_nl, mux_1933_nl, fsm_output(6));
  or_4104_nl <= (fsm_output(2)) OR mux_1937_nl;
  mux_1945_nl <= MUX_s_1_2_2(nand_431_nl, or_4104_nl, fsm_output(5));
  vec_rsc_0_38_i_we_d_pff <= NOT(mux_1945_nl OR (fsm_output(1)));
  or_2319_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2318_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1958_nl <= MUX_s_1_2_2(or_2319_nl, or_2318_nl, fsm_output(0));
  or_2320_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1958_nl;
  or_2316_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00110")) OR not_tmp_452;
  mux_1955_nl <= MUX_s_1_2_2(or_2316_nl, or_tmp_2172, fsm_output(0));
  or_2314_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100110")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1954_nl <= MUX_s_1_2_2(or_2314_nl, or_tmp_2168, fsm_output(0));
  mux_1956_nl <= MUX_s_1_2_2(mux_1955_nl, mux_1954_nl, fsm_output(4));
  or_2313_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100110")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1952_nl <= MUX_s_1_2_2(or_2313_nl, or_tmp_2166, fsm_output(0));
  or_2311_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100110")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1951_nl <= MUX_s_1_2_2(or_2311_nl, or_tmp_2162, fsm_output(0));
  mux_1953_nl <= MUX_s_1_2_2(mux_1952_nl, mux_1951_nl, fsm_output(4));
  mux_1957_nl <= MUX_s_1_2_2(mux_1956_nl, mux_1953_nl, fsm_output(6));
  mux_1959_nl <= MUX_s_1_2_2(or_2320_nl, mux_1957_nl, fsm_output(2));
  or_2309_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2307_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (NOT and_763_cse);
  mux_1948_nl <= MUX_s_1_2_2(or_2309_nl, or_2307_nl, fsm_output(0));
  or_2305_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2304_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1947_nl <= MUX_s_1_2_2(or_2305_nl, or_2304_nl, fsm_output(0));
  mux_1949_nl <= MUX_s_1_2_2(mux_1948_nl, mux_1947_nl, fsm_output(4));
  nor_998_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_999_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1946_nl <= MUX_s_1_2_2(nor_998_nl, nor_999_nl, fsm_output(0));
  nand_91_nl <= NOT((fsm_output(4)) AND mux_1946_nl);
  mux_1950_nl <= MUX_s_1_2_2(mux_1949_nl, nand_91_nl, fsm_output(6));
  or_2310_nl <= (fsm_output(2)) OR mux_1950_nl;
  mux_1960_nl <= MUX_s_1_2_2(mux_1959_nl, or_2310_nl, fsm_output(5));
  vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1960_nl) AND (fsm_output(1));
  and_590_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("100111"))
      AND and_763_cse;
  nor_990_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("100"))
      OR not_tmp_347);
  mux_1972_nl <= MUX_s_1_2_2(and_590_nl, nor_990_nl, fsm_output(0));
  nor_991_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_992_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_1971_nl <= MUX_s_1_2_2(nor_991_nl, nor_992_nl, fsm_output(0));
  mux_1973_nl <= MUX_s_1_2_2(mux_1972_nl, mux_1971_nl, fsm_output(4));
  nor_993_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_994_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1969_nl <= MUX_s_1_2_2(nor_993_nl, nor_994_nl, fsm_output(0));
  nor_995_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_996_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1968_nl <= MUX_s_1_2_2(nor_995_nl, nor_996_nl, fsm_output(0));
  mux_1970_nl <= MUX_s_1_2_2(mux_1969_nl, mux_1968_nl, fsm_output(4));
  mux_1974_nl <= MUX_s_1_2_2(mux_1973_nl, mux_1970_nl, fsm_output(6));
  nand_430_nl <= NOT((fsm_output(2)) AND mux_1974_nl);
  or_2330_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR not_tmp_452;
  mux_1965_nl <= MUX_s_1_2_2(or_tmp_2216, or_2330_nl, fsm_output(0));
  or_2327_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1964_nl <= MUX_s_1_2_2(or_tmp_2212, or_2327_nl, fsm_output(0));
  mux_1966_nl <= MUX_s_1_2_2(mux_1965_nl, mux_1964_nl, fsm_output(4));
  or_2324_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1962_nl <= MUX_s_1_2_2(or_tmp_2210, or_2324_nl, fsm_output(0));
  or_2321_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1961_nl <= MUX_s_1_2_2(or_tmp_2206, or_2321_nl, fsm_output(0));
  mux_1963_nl <= MUX_s_1_2_2(mux_1962_nl, mux_1961_nl, fsm_output(4));
  mux_1967_nl <= MUX_s_1_2_2(mux_1966_nl, mux_1963_nl, fsm_output(6));
  or_4103_nl <= (fsm_output(2)) OR mux_1967_nl;
  mux_1975_nl <= MUX_s_1_2_2(nand_430_nl, or_4103_nl, fsm_output(5));
  vec_rsc_0_39_i_we_d_pff <= NOT(mux_1975_nl OR (fsm_output(1)));
  or_2363_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2362_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1988_nl <= MUX_s_1_2_2(or_2363_nl, or_2362_nl, fsm_output(0));
  or_2364_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_1988_nl;
  or_2360_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00111")) OR not_tmp_452;
  mux_1985_nl <= MUX_s_1_2_2(or_2360_nl, or_tmp_2216, fsm_output(0));
  or_2358_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100111")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1984_nl <= MUX_s_1_2_2(or_2358_nl, or_tmp_2212, fsm_output(0));
  mux_1986_nl <= MUX_s_1_2_2(mux_1985_nl, mux_1984_nl, fsm_output(4));
  or_2357_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100111")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1982_nl <= MUX_s_1_2_2(or_2357_nl, or_tmp_2210, fsm_output(0));
  or_2355_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100111")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_1981_nl <= MUX_s_1_2_2(or_2355_nl, or_tmp_2206, fsm_output(0));
  mux_1983_nl <= MUX_s_1_2_2(mux_1982_nl, mux_1981_nl, fsm_output(4));
  mux_1987_nl <= MUX_s_1_2_2(mux_1986_nl, mux_1983_nl, fsm_output(6));
  mux_1989_nl <= MUX_s_1_2_2(or_2364_nl, mux_1987_nl, fsm_output(2));
  or_2353_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  nand_296_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("100111"))
      AND and_763_cse);
  mux_1978_nl <= MUX_s_1_2_2(or_2353_nl, nand_296_nl, fsm_output(0));
  or_2349_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2348_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1977_nl <= MUX_s_1_2_2(or_2349_nl, or_2348_nl, fsm_output(0));
  mux_1979_nl <= MUX_s_1_2_2(mux_1978_nl, mux_1977_nl, fsm_output(4));
  nor_988_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_989_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1976_nl <= MUX_s_1_2_2(nor_988_nl, nor_989_nl, fsm_output(0));
  nand_93_nl <= NOT((fsm_output(4)) AND mux_1976_nl);
  mux_1980_nl <= MUX_s_1_2_2(mux_1979_nl, nand_93_nl, fsm_output(6));
  or_2354_nl <= (fsm_output(2)) OR mux_1980_nl;
  mux_1990_nl <= MUX_s_1_2_2(mux_1989_nl, or_2354_nl, fsm_output(5));
  vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_1990_nl) AND (fsm_output(1));
  nor_979_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (NOT and_763_cse));
  nor_980_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_2002_nl <= MUX_s_1_2_2(nor_979_nl, nor_980_nl, fsm_output(0));
  nor_981_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_982_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2001_nl <= MUX_s_1_2_2(nor_981_nl, nor_982_nl, fsm_output(0));
  mux_2003_nl <= MUX_s_1_2_2(mux_2002_nl, mux_2001_nl, fsm_output(4));
  nor_983_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_984_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_1999_nl <= MUX_s_1_2_2(nor_983_nl, nor_984_nl, fsm_output(0));
  nor_985_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_986_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_1998_nl <= MUX_s_1_2_2(nor_985_nl, nor_986_nl, fsm_output(0));
  mux_2000_nl <= MUX_s_1_2_2(mux_1999_nl, mux_1998_nl, fsm_output(4));
  mux_2004_nl <= MUX_s_1_2_2(mux_2003_nl, mux_2000_nl, fsm_output(6));
  nand_429_nl <= NOT((fsm_output(2)) AND mux_2004_nl);
  or_2374_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR not_tmp_452;
  mux_1995_nl <= MUX_s_1_2_2(or_tmp_2260, or_2374_nl, fsm_output(0));
  or_2371_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_1994_nl <= MUX_s_1_2_2(or_tmp_2256, or_2371_nl, fsm_output(0));
  mux_1996_nl <= MUX_s_1_2_2(mux_1995_nl, mux_1994_nl, fsm_output(4));
  or_2368_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_1992_nl <= MUX_s_1_2_2(or_tmp_2254, or_2368_nl, fsm_output(0));
  or_2365_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_1991_nl <= MUX_s_1_2_2(or_tmp_2250, or_2365_nl, fsm_output(0));
  mux_1993_nl <= MUX_s_1_2_2(mux_1992_nl, mux_1991_nl, fsm_output(4));
  mux_1997_nl <= MUX_s_1_2_2(mux_1996_nl, mux_1993_nl, fsm_output(6));
  or_4102_nl <= (fsm_output(2)) OR mux_1997_nl;
  mux_2005_nl <= MUX_s_1_2_2(nand_429_nl, or_4102_nl, fsm_output(5));
  vec_rsc_0_40_i_we_d_pff <= NOT(mux_2005_nl OR (fsm_output(1)));
  or_2407_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2406_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2018_nl <= MUX_s_1_2_2(or_2407_nl, or_2406_nl, fsm_output(0));
  or_2408_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2018_nl;
  or_2404_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01000")) OR not_tmp_452;
  mux_2015_nl <= MUX_s_1_2_2(or_2404_nl, or_tmp_2260, fsm_output(0));
  or_2402_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101000")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2014_nl <= MUX_s_1_2_2(or_2402_nl, or_tmp_2256, fsm_output(0));
  mux_2016_nl <= MUX_s_1_2_2(mux_2015_nl, mux_2014_nl, fsm_output(4));
  or_2401_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101000")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2012_nl <= MUX_s_1_2_2(or_2401_nl, or_tmp_2254, fsm_output(0));
  or_2399_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101000")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2011_nl <= MUX_s_1_2_2(or_2399_nl, or_tmp_2250, fsm_output(0));
  mux_2013_nl <= MUX_s_1_2_2(mux_2012_nl, mux_2011_nl, fsm_output(4));
  mux_2017_nl <= MUX_s_1_2_2(mux_2016_nl, mux_2013_nl, fsm_output(6));
  mux_2019_nl <= MUX_s_1_2_2(or_2408_nl, mux_2017_nl, fsm_output(2));
  or_2397_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2395_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (NOT and_763_cse);
  mux_2008_nl <= MUX_s_1_2_2(or_2397_nl, or_2395_nl, fsm_output(0));
  or_2393_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2392_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2007_nl <= MUX_s_1_2_2(or_2393_nl, or_2392_nl, fsm_output(0));
  mux_2009_nl <= MUX_s_1_2_2(mux_2008_nl, mux_2007_nl, fsm_output(4));
  nor_977_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_978_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2006_nl <= MUX_s_1_2_2(nor_977_nl, nor_978_nl, fsm_output(0));
  nand_95_nl <= NOT((fsm_output(4)) AND mux_2006_nl);
  mux_2010_nl <= MUX_s_1_2_2(mux_2009_nl, nand_95_nl, fsm_output(6));
  or_2398_nl <= (fsm_output(2)) OR mux_2010_nl;
  mux_2020_nl <= MUX_s_1_2_2(mux_2019_nl, or_2398_nl, fsm_output(5));
  vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2020_nl) AND (fsm_output(1));
  nor_968_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (NOT and_763_cse));
  nor_969_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_2032_nl <= MUX_s_1_2_2(nor_968_nl, nor_969_nl, fsm_output(0));
  nor_970_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_971_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2031_nl <= MUX_s_1_2_2(nor_970_nl, nor_971_nl, fsm_output(0));
  mux_2033_nl <= MUX_s_1_2_2(mux_2032_nl, mux_2031_nl, fsm_output(4));
  nor_972_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_973_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2029_nl <= MUX_s_1_2_2(nor_972_nl, nor_973_nl, fsm_output(0));
  nor_974_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_975_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2028_nl <= MUX_s_1_2_2(nor_974_nl, nor_975_nl, fsm_output(0));
  mux_2030_nl <= MUX_s_1_2_2(mux_2029_nl, mux_2028_nl, fsm_output(4));
  mux_2034_nl <= MUX_s_1_2_2(mux_2033_nl, mux_2030_nl, fsm_output(6));
  nand_428_nl <= NOT((fsm_output(2)) AND mux_2034_nl);
  or_2418_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR not_tmp_452;
  mux_2025_nl <= MUX_s_1_2_2(or_tmp_2304, or_2418_nl, fsm_output(0));
  or_2415_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2024_nl <= MUX_s_1_2_2(or_tmp_2300, or_2415_nl, fsm_output(0));
  mux_2026_nl <= MUX_s_1_2_2(mux_2025_nl, mux_2024_nl, fsm_output(4));
  or_2412_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2022_nl <= MUX_s_1_2_2(or_tmp_2298, or_2412_nl, fsm_output(0));
  or_2409_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2021_nl <= MUX_s_1_2_2(or_tmp_2294, or_2409_nl, fsm_output(0));
  mux_2023_nl <= MUX_s_1_2_2(mux_2022_nl, mux_2021_nl, fsm_output(4));
  mux_2027_nl <= MUX_s_1_2_2(mux_2026_nl, mux_2023_nl, fsm_output(6));
  or_4101_nl <= (fsm_output(2)) OR mux_2027_nl;
  mux_2035_nl <= MUX_s_1_2_2(nand_428_nl, or_4101_nl, fsm_output(5));
  vec_rsc_0_41_i_we_d_pff <= NOT(mux_2035_nl OR (fsm_output(1)));
  or_2451_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2450_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2048_nl <= MUX_s_1_2_2(or_2451_nl, or_2450_nl, fsm_output(0));
  or_2452_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2048_nl;
  or_2448_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01001")) OR not_tmp_452;
  mux_2045_nl <= MUX_s_1_2_2(or_2448_nl, or_tmp_2304, fsm_output(0));
  or_2446_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101001")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2044_nl <= MUX_s_1_2_2(or_2446_nl, or_tmp_2300, fsm_output(0));
  mux_2046_nl <= MUX_s_1_2_2(mux_2045_nl, mux_2044_nl, fsm_output(4));
  or_2445_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101001")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2042_nl <= MUX_s_1_2_2(or_2445_nl, or_tmp_2298, fsm_output(0));
  or_2443_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101001")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2041_nl <= MUX_s_1_2_2(or_2443_nl, or_tmp_2294, fsm_output(0));
  mux_2043_nl <= MUX_s_1_2_2(mux_2042_nl, mux_2041_nl, fsm_output(4));
  mux_2047_nl <= MUX_s_1_2_2(mux_2046_nl, mux_2043_nl, fsm_output(6));
  mux_2049_nl <= MUX_s_1_2_2(or_2452_nl, mux_2047_nl, fsm_output(2));
  or_2441_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_2439_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (NOT and_763_cse);
  mux_2038_nl <= MUX_s_1_2_2(or_2441_nl, or_2439_nl, fsm_output(0));
  or_2437_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2436_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2037_nl <= MUX_s_1_2_2(or_2437_nl, or_2436_nl, fsm_output(0));
  mux_2039_nl <= MUX_s_1_2_2(mux_2038_nl, mux_2037_nl, fsm_output(4));
  nor_966_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_967_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2036_nl <= MUX_s_1_2_2(nor_966_nl, nor_967_nl, fsm_output(0));
  nand_97_nl <= NOT((fsm_output(4)) AND mux_2036_nl);
  mux_2040_nl <= MUX_s_1_2_2(mux_2039_nl, nand_97_nl, fsm_output(6));
  or_2442_nl <= (fsm_output(2)) OR mux_2040_nl;
  mux_2050_nl <= MUX_s_1_2_2(mux_2049_nl, or_2442_nl, fsm_output(5));
  vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2050_nl) AND (fsm_output(1));
  nor_957_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (NOT and_763_cse));
  nor_958_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_2062_nl <= MUX_s_1_2_2(nor_957_nl, nor_958_nl, fsm_output(0));
  nor_959_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_960_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2061_nl <= MUX_s_1_2_2(nor_959_nl, nor_960_nl, fsm_output(0));
  mux_2063_nl <= MUX_s_1_2_2(mux_2062_nl, mux_2061_nl, fsm_output(4));
  nor_961_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_962_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2059_nl <= MUX_s_1_2_2(nor_961_nl, nor_962_nl, fsm_output(0));
  nor_963_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_964_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2058_nl <= MUX_s_1_2_2(nor_963_nl, nor_964_nl, fsm_output(0));
  mux_2060_nl <= MUX_s_1_2_2(mux_2059_nl, mux_2058_nl, fsm_output(4));
  mux_2064_nl <= MUX_s_1_2_2(mux_2063_nl, mux_2060_nl, fsm_output(6));
  nand_427_nl <= NOT((fsm_output(2)) AND mux_2064_nl);
  or_2462_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR not_tmp_452;
  mux_2055_nl <= MUX_s_1_2_2(or_tmp_2348, or_2462_nl, fsm_output(0));
  or_2459_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2054_nl <= MUX_s_1_2_2(or_tmp_2344, or_2459_nl, fsm_output(0));
  mux_2056_nl <= MUX_s_1_2_2(mux_2055_nl, mux_2054_nl, fsm_output(4));
  or_2456_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2052_nl <= MUX_s_1_2_2(or_tmp_2342, or_2456_nl, fsm_output(0));
  or_2453_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2051_nl <= MUX_s_1_2_2(or_tmp_2338, or_2453_nl, fsm_output(0));
  mux_2053_nl <= MUX_s_1_2_2(mux_2052_nl, mux_2051_nl, fsm_output(4));
  mux_2057_nl <= MUX_s_1_2_2(mux_2056_nl, mux_2053_nl, fsm_output(6));
  or_4100_nl <= (fsm_output(2)) OR mux_2057_nl;
  mux_2065_nl <= MUX_s_1_2_2(nand_427_nl, or_4100_nl, fsm_output(5));
  vec_rsc_0_42_i_we_d_pff <= NOT(mux_2065_nl OR (fsm_output(1)));
  or_2495_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2494_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2078_nl <= MUX_s_1_2_2(or_2495_nl, or_2494_nl, fsm_output(0));
  or_2496_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2078_nl;
  or_2492_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01010")) OR not_tmp_452;
  mux_2075_nl <= MUX_s_1_2_2(or_2492_nl, or_tmp_2348, fsm_output(0));
  or_2490_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101010")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2074_nl <= MUX_s_1_2_2(or_2490_nl, or_tmp_2344, fsm_output(0));
  mux_2076_nl <= MUX_s_1_2_2(mux_2075_nl, mux_2074_nl, fsm_output(4));
  or_2489_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101010")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2072_nl <= MUX_s_1_2_2(or_2489_nl, or_tmp_2342, fsm_output(0));
  or_2487_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101010")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2071_nl <= MUX_s_1_2_2(or_2487_nl, or_tmp_2338, fsm_output(0));
  mux_2073_nl <= MUX_s_1_2_2(mux_2072_nl, mux_2071_nl, fsm_output(4));
  mux_2077_nl <= MUX_s_1_2_2(mux_2076_nl, mux_2073_nl, fsm_output(6));
  mux_2079_nl <= MUX_s_1_2_2(or_2496_nl, mux_2077_nl, fsm_output(2));
  or_2485_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2483_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (NOT and_763_cse);
  mux_2068_nl <= MUX_s_1_2_2(or_2485_nl, or_2483_nl, fsm_output(0));
  or_2481_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2480_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2067_nl <= MUX_s_1_2_2(or_2481_nl, or_2480_nl, fsm_output(0));
  mux_2069_nl <= MUX_s_1_2_2(mux_2068_nl, mux_2067_nl, fsm_output(4));
  nor_955_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_956_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2066_nl <= MUX_s_1_2_2(nor_955_nl, nor_956_nl, fsm_output(0));
  nand_99_nl <= NOT((fsm_output(4)) AND mux_2066_nl);
  mux_2070_nl <= MUX_s_1_2_2(mux_2069_nl, nand_99_nl, fsm_output(6));
  or_2486_nl <= (fsm_output(2)) OR mux_2070_nl;
  mux_2080_nl <= MUX_s_1_2_2(mux_2079_nl, or_2486_nl, fsm_output(5));
  vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2080_nl) AND (fsm_output(1));
  and_585_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101011"))
      AND and_763_cse;
  nor_947_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR not_tmp_330);
  mux_2092_nl <= MUX_s_1_2_2(and_585_nl, nor_947_nl, fsm_output(0));
  nor_948_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_949_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2091_nl <= MUX_s_1_2_2(nor_948_nl, nor_949_nl, fsm_output(0));
  mux_2093_nl <= MUX_s_1_2_2(mux_2092_nl, mux_2091_nl, fsm_output(4));
  nor_950_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_951_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2089_nl <= MUX_s_1_2_2(nor_950_nl, nor_951_nl, fsm_output(0));
  nor_952_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_953_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2088_nl <= MUX_s_1_2_2(nor_952_nl, nor_953_nl, fsm_output(0));
  mux_2090_nl <= MUX_s_1_2_2(mux_2089_nl, mux_2088_nl, fsm_output(4));
  mux_2094_nl <= MUX_s_1_2_2(mux_2093_nl, mux_2090_nl, fsm_output(6));
  nand_426_nl <= NOT((fsm_output(2)) AND mux_2094_nl);
  or_2506_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR not_tmp_452;
  mux_2085_nl <= MUX_s_1_2_2(or_tmp_2392, or_2506_nl, fsm_output(0));
  or_2503_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2084_nl <= MUX_s_1_2_2(or_tmp_2388, or_2503_nl, fsm_output(0));
  mux_2086_nl <= MUX_s_1_2_2(mux_2085_nl, mux_2084_nl, fsm_output(4));
  or_2500_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2082_nl <= MUX_s_1_2_2(or_tmp_2386, or_2500_nl, fsm_output(0));
  or_2497_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2081_nl <= MUX_s_1_2_2(or_tmp_2382, or_2497_nl, fsm_output(0));
  mux_2083_nl <= MUX_s_1_2_2(mux_2082_nl, mux_2081_nl, fsm_output(4));
  mux_2087_nl <= MUX_s_1_2_2(mux_2086_nl, mux_2083_nl, fsm_output(6));
  or_4099_nl <= (fsm_output(2)) OR mux_2087_nl;
  mux_2095_nl <= MUX_s_1_2_2(nand_426_nl, or_4099_nl, fsm_output(5));
  vec_rsc_0_43_i_we_d_pff <= NOT(mux_2095_nl OR (fsm_output(1)));
  or_2539_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2538_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2108_nl <= MUX_s_1_2_2(or_2539_nl, or_2538_nl, fsm_output(0));
  or_2540_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2108_nl;
  or_2536_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01011")) OR not_tmp_452;
  mux_2105_nl <= MUX_s_1_2_2(or_2536_nl, or_tmp_2392, fsm_output(0));
  or_2534_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101011")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2104_nl <= MUX_s_1_2_2(or_2534_nl, or_tmp_2388, fsm_output(0));
  mux_2106_nl <= MUX_s_1_2_2(mux_2105_nl, mux_2104_nl, fsm_output(4));
  or_2533_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101011")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2102_nl <= MUX_s_1_2_2(or_2533_nl, or_tmp_2386, fsm_output(0));
  or_2531_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101011")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2101_nl <= MUX_s_1_2_2(or_2531_nl, or_tmp_2382, fsm_output(0));
  mux_2103_nl <= MUX_s_1_2_2(mux_2102_nl, mux_2101_nl, fsm_output(4));
  mux_2107_nl <= MUX_s_1_2_2(mux_2106_nl, mux_2103_nl, fsm_output(6));
  mux_2109_nl <= MUX_s_1_2_2(or_2540_nl, mux_2107_nl, fsm_output(2));
  or_2529_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  nand_295_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101011"))
      AND and_763_cse);
  mux_2098_nl <= MUX_s_1_2_2(or_2529_nl, nand_295_nl, fsm_output(0));
  or_2525_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2524_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2097_nl <= MUX_s_1_2_2(or_2525_nl, or_2524_nl, fsm_output(0));
  mux_2099_nl <= MUX_s_1_2_2(mux_2098_nl, mux_2097_nl, fsm_output(4));
  nor_945_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_946_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2096_nl <= MUX_s_1_2_2(nor_945_nl, nor_946_nl, fsm_output(0));
  nand_101_nl <= NOT((fsm_output(4)) AND mux_2096_nl);
  mux_2100_nl <= MUX_s_1_2_2(mux_2099_nl, nand_101_nl, fsm_output(6));
  or_2530_nl <= (fsm_output(2)) OR mux_2100_nl;
  mux_2110_nl <= MUX_s_1_2_2(mux_2109_nl, or_2530_nl, fsm_output(5));
  vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2110_nl) AND (fsm_output(1));
  nor_936_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (NOT and_763_cse));
  nor_937_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_2122_nl <= MUX_s_1_2_2(nor_936_nl, nor_937_nl, fsm_output(0));
  nor_938_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_939_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2121_nl <= MUX_s_1_2_2(nor_938_nl, nor_939_nl, fsm_output(0));
  mux_2123_nl <= MUX_s_1_2_2(mux_2122_nl, mux_2121_nl, fsm_output(4));
  nor_940_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_941_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2119_nl <= MUX_s_1_2_2(nor_940_nl, nor_941_nl, fsm_output(0));
  nor_942_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_943_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2118_nl <= MUX_s_1_2_2(nor_942_nl, nor_943_nl, fsm_output(0));
  mux_2120_nl <= MUX_s_1_2_2(mux_2119_nl, mux_2118_nl, fsm_output(4));
  mux_2124_nl <= MUX_s_1_2_2(mux_2123_nl, mux_2120_nl, fsm_output(6));
  nand_425_nl <= NOT((fsm_output(2)) AND mux_2124_nl);
  or_2550_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR not_tmp_452;
  mux_2115_nl <= MUX_s_1_2_2(or_tmp_2436, or_2550_nl, fsm_output(0));
  or_2547_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2114_nl <= MUX_s_1_2_2(or_tmp_2432, or_2547_nl, fsm_output(0));
  mux_2116_nl <= MUX_s_1_2_2(mux_2115_nl, mux_2114_nl, fsm_output(4));
  or_2544_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2112_nl <= MUX_s_1_2_2(or_tmp_2430, or_2544_nl, fsm_output(0));
  or_2541_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2111_nl <= MUX_s_1_2_2(or_tmp_2426, or_2541_nl, fsm_output(0));
  mux_2113_nl <= MUX_s_1_2_2(mux_2112_nl, mux_2111_nl, fsm_output(4));
  mux_2117_nl <= MUX_s_1_2_2(mux_2116_nl, mux_2113_nl, fsm_output(6));
  or_4098_nl <= (fsm_output(2)) OR mux_2117_nl;
  mux_2125_nl <= MUX_s_1_2_2(nand_425_nl, or_4098_nl, fsm_output(5));
  vec_rsc_0_44_i_we_d_pff <= NOT(mux_2125_nl OR (fsm_output(1)));
  or_2583_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2582_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2138_nl <= MUX_s_1_2_2(or_2583_nl, or_2582_nl, fsm_output(0));
  or_2584_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2138_nl;
  or_2580_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01100")) OR not_tmp_452;
  mux_2135_nl <= MUX_s_1_2_2(or_2580_nl, or_tmp_2436, fsm_output(0));
  or_2578_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101100")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2134_nl <= MUX_s_1_2_2(or_2578_nl, or_tmp_2432, fsm_output(0));
  mux_2136_nl <= MUX_s_1_2_2(mux_2135_nl, mux_2134_nl, fsm_output(4));
  or_2577_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101100")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2132_nl <= MUX_s_1_2_2(or_2577_nl, or_tmp_2430, fsm_output(0));
  or_2575_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101100")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2131_nl <= MUX_s_1_2_2(or_2575_nl, or_tmp_2426, fsm_output(0));
  mux_2133_nl <= MUX_s_1_2_2(mux_2132_nl, mux_2131_nl, fsm_output(4));
  mux_2137_nl <= MUX_s_1_2_2(mux_2136_nl, mux_2133_nl, fsm_output(6));
  mux_2139_nl <= MUX_s_1_2_2(or_2584_nl, mux_2137_nl, fsm_output(2));
  or_2573_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2571_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (NOT and_763_cse);
  mux_2128_nl <= MUX_s_1_2_2(or_2573_nl, or_2571_nl, fsm_output(0));
  or_2569_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2568_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2127_nl <= MUX_s_1_2_2(or_2569_nl, or_2568_nl, fsm_output(0));
  mux_2129_nl <= MUX_s_1_2_2(mux_2128_nl, mux_2127_nl, fsm_output(4));
  nor_934_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_935_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2126_nl <= MUX_s_1_2_2(nor_934_nl, nor_935_nl, fsm_output(0));
  nand_103_nl <= NOT((fsm_output(4)) AND mux_2126_nl);
  mux_2130_nl <= MUX_s_1_2_2(mux_2129_nl, nand_103_nl, fsm_output(6));
  or_2574_nl <= (fsm_output(2)) OR mux_2130_nl;
  mux_2140_nl <= MUX_s_1_2_2(mux_2139_nl, or_2574_nl, fsm_output(5));
  vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2140_nl) AND (fsm_output(1));
  and_582_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101101"))
      AND and_763_cse;
  nor_926_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_2152_nl <= MUX_s_1_2_2(and_582_nl, nor_926_nl, fsm_output(0));
  nor_927_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_928_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2151_nl <= MUX_s_1_2_2(nor_927_nl, nor_928_nl, fsm_output(0));
  mux_2153_nl <= MUX_s_1_2_2(mux_2152_nl, mux_2151_nl, fsm_output(4));
  nor_929_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_930_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2149_nl <= MUX_s_1_2_2(nor_929_nl, nor_930_nl, fsm_output(0));
  nor_931_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_932_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2148_nl <= MUX_s_1_2_2(nor_931_nl, nor_932_nl, fsm_output(0));
  mux_2150_nl <= MUX_s_1_2_2(mux_2149_nl, mux_2148_nl, fsm_output(4));
  mux_2154_nl <= MUX_s_1_2_2(mux_2153_nl, mux_2150_nl, fsm_output(6));
  nand_424_nl <= NOT((fsm_output(2)) AND mux_2154_nl);
  or_2594_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR not_tmp_452;
  mux_2145_nl <= MUX_s_1_2_2(or_tmp_2480, or_2594_nl, fsm_output(0));
  or_2591_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2144_nl <= MUX_s_1_2_2(or_tmp_2476, or_2591_nl, fsm_output(0));
  mux_2146_nl <= MUX_s_1_2_2(mux_2145_nl, mux_2144_nl, fsm_output(4));
  or_2588_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2142_nl <= MUX_s_1_2_2(or_tmp_2474, or_2588_nl, fsm_output(0));
  or_2585_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2141_nl <= MUX_s_1_2_2(or_tmp_2470, or_2585_nl, fsm_output(0));
  mux_2143_nl <= MUX_s_1_2_2(mux_2142_nl, mux_2141_nl, fsm_output(4));
  mux_2147_nl <= MUX_s_1_2_2(mux_2146_nl, mux_2143_nl, fsm_output(6));
  or_4097_nl <= (fsm_output(2)) OR mux_2147_nl;
  mux_2155_nl <= MUX_s_1_2_2(nand_424_nl, or_4097_nl, fsm_output(5));
  vec_rsc_0_45_i_we_d_pff <= NOT(mux_2155_nl OR (fsm_output(1)));
  or_2627_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2626_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2168_nl <= MUX_s_1_2_2(or_2627_nl, or_2626_nl, fsm_output(0));
  or_2628_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2168_nl;
  or_2624_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01101")) OR not_tmp_452;
  mux_2165_nl <= MUX_s_1_2_2(or_2624_nl, or_tmp_2480, fsm_output(0));
  or_2622_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101101")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2164_nl <= MUX_s_1_2_2(or_2622_nl, or_tmp_2476, fsm_output(0));
  mux_2166_nl <= MUX_s_1_2_2(mux_2165_nl, mux_2164_nl, fsm_output(4));
  or_2621_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101101")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2162_nl <= MUX_s_1_2_2(or_2621_nl, or_tmp_2474, fsm_output(0));
  or_2619_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101101")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2161_nl <= MUX_s_1_2_2(or_2619_nl, or_tmp_2470, fsm_output(0));
  mux_2163_nl <= MUX_s_1_2_2(mux_2162_nl, mux_2161_nl, fsm_output(4));
  mux_2167_nl <= MUX_s_1_2_2(mux_2166_nl, mux_2163_nl, fsm_output(6));
  mux_2169_nl <= MUX_s_1_2_2(or_2628_nl, mux_2167_nl, fsm_output(2));
  or_2617_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  nand_294_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101101"))
      AND and_763_cse);
  mux_2158_nl <= MUX_s_1_2_2(or_2617_nl, nand_294_nl, fsm_output(0));
  or_2613_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2612_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2157_nl <= MUX_s_1_2_2(or_2613_nl, or_2612_nl, fsm_output(0));
  mux_2159_nl <= MUX_s_1_2_2(mux_2158_nl, mux_2157_nl, fsm_output(4));
  nor_924_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_925_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2156_nl <= MUX_s_1_2_2(nor_924_nl, nor_925_nl, fsm_output(0));
  nand_105_nl <= NOT((fsm_output(4)) AND mux_2156_nl);
  mux_2160_nl <= MUX_s_1_2_2(mux_2159_nl, nand_105_nl, fsm_output(6));
  or_2618_nl <= (fsm_output(2)) OR mux_2160_nl;
  mux_2170_nl <= MUX_s_1_2_2(mux_2169_nl, or_2618_nl, fsm_output(5));
  vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2170_nl) AND (fsm_output(1));
  and_579_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101110"))
      AND and_763_cse;
  and_580_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND and_763_cse;
  mux_2182_nl <= MUX_s_1_2_2(and_579_nl, and_580_nl, fsm_output(0));
  nor_917_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_918_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2181_nl <= MUX_s_1_2_2(nor_917_nl, nor_918_nl, fsm_output(0));
  mux_2183_nl <= MUX_s_1_2_2(mux_2182_nl, mux_2181_nl, fsm_output(4));
  nor_919_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_920_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2179_nl <= MUX_s_1_2_2(nor_919_nl, nor_920_nl, fsm_output(0));
  nor_921_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_922_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2178_nl <= MUX_s_1_2_2(nor_921_nl, nor_922_nl, fsm_output(0));
  mux_2180_nl <= MUX_s_1_2_2(mux_2179_nl, mux_2178_nl, fsm_output(4));
  mux_2184_nl <= MUX_s_1_2_2(mux_2183_nl, mux_2180_nl, fsm_output(6));
  nand_423_nl <= NOT((fsm_output(2)) AND mux_2184_nl);
  or_2638_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR not_tmp_452;
  mux_2175_nl <= MUX_s_1_2_2(or_tmp_2524, or_2638_nl, fsm_output(0));
  or_2635_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2174_nl <= MUX_s_1_2_2(or_tmp_2520, or_2635_nl, fsm_output(0));
  mux_2176_nl <= MUX_s_1_2_2(mux_2175_nl, mux_2174_nl, fsm_output(4));
  or_2632_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2172_nl <= MUX_s_1_2_2(or_tmp_2518, or_2632_nl, fsm_output(0));
  or_2629_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2171_nl <= MUX_s_1_2_2(or_tmp_2514, or_2629_nl, fsm_output(0));
  mux_2173_nl <= MUX_s_1_2_2(mux_2172_nl, mux_2171_nl, fsm_output(4));
  mux_2177_nl <= MUX_s_1_2_2(mux_2176_nl, mux_2173_nl, fsm_output(6));
  or_4096_nl <= (fsm_output(2)) OR mux_2177_nl;
  mux_2185_nl <= MUX_s_1_2_2(nand_423_nl, or_4096_nl, fsm_output(5));
  vec_rsc_0_46_i_we_d_pff <= NOT(mux_2185_nl OR (fsm_output(1)));
  or_2671_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2670_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2198_nl <= MUX_s_1_2_2(or_2671_nl, or_2670_nl, fsm_output(0));
  or_2672_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2198_nl;
  or_2668_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01110")) OR not_tmp_452;
  mux_2195_nl <= MUX_s_1_2_2(or_2668_nl, or_tmp_2524, fsm_output(0));
  or_2666_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101110")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2194_nl <= MUX_s_1_2_2(or_2666_nl, or_tmp_2520, fsm_output(0));
  mux_2196_nl <= MUX_s_1_2_2(mux_2195_nl, mux_2194_nl, fsm_output(4));
  or_2665_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101110")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2192_nl <= MUX_s_1_2_2(or_2665_nl, or_tmp_2518, fsm_output(0));
  or_2663_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101110")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2191_nl <= MUX_s_1_2_2(or_2663_nl, or_tmp_2514, fsm_output(0));
  mux_2193_nl <= MUX_s_1_2_2(mux_2192_nl, mux_2191_nl, fsm_output(4));
  mux_2197_nl <= MUX_s_1_2_2(mux_2196_nl, mux_2193_nl, fsm_output(6));
  mux_2199_nl <= MUX_s_1_2_2(or_2672_nl, mux_2197_nl, fsm_output(2));
  nand_292_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND and_763_cse);
  nand_293_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101110"))
      AND and_763_cse);
  mux_2188_nl <= MUX_s_1_2_2(nand_292_nl, nand_293_nl, fsm_output(0));
  or_2657_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2656_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2187_nl <= MUX_s_1_2_2(or_2657_nl, or_2656_nl, fsm_output(0));
  mux_2189_nl <= MUX_s_1_2_2(mux_2188_nl, mux_2187_nl, fsm_output(4));
  nor_915_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_916_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2186_nl <= MUX_s_1_2_2(nor_915_nl, nor_916_nl, fsm_output(0));
  nand_107_nl <= NOT((fsm_output(4)) AND mux_2186_nl);
  mux_2190_nl <= MUX_s_1_2_2(mux_2189_nl, nand_107_nl, fsm_output(6));
  or_2662_nl <= (fsm_output(2)) OR mux_2190_nl;
  mux_2200_nl <= MUX_s_1_2_2(mux_2199_nl, or_2662_nl, fsm_output(5));
  vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2200_nl) AND (fsm_output(1));
  and_575_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND and_763_cse;
  nor_909_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("101"))
      OR not_tmp_347);
  mux_2212_nl <= MUX_s_1_2_2(and_575_nl, nor_909_nl, fsm_output(0));
  and_576_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_577_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  mux_2211_nl <= MUX_s_1_2_2(and_576_nl, and_577_nl, fsm_output(0));
  mux_2213_nl <= MUX_s_1_2_2(mux_2212_nl, mux_2211_nl, fsm_output(4));
  and_812_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7));
  and_819_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT (fsm_output(3))) AND (fsm_output(7));
  mux_2209_nl <= MUX_s_1_2_2(and_812_nl, and_819_nl, fsm_output(0));
  nor_912_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_913_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2208_nl <= MUX_s_1_2_2(nor_912_nl, nor_913_nl, fsm_output(0));
  mux_2210_nl <= MUX_s_1_2_2(mux_2209_nl, mux_2208_nl, fsm_output(4));
  mux_2214_nl <= MUX_s_1_2_2(mux_2213_nl, mux_2210_nl, fsm_output(6));
  nand_422_nl <= NOT((fsm_output(2)) AND mux_2214_nl);
  or_2682_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("01111"))))
      OR not_tmp_452;
  mux_2205_nl <= MUX_s_1_2_2(or_tmp_2567, or_2682_nl, fsm_output(0));
  nand_287_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2204_nl <= MUX_s_1_2_2(or_tmp_2564, nand_287_nl, fsm_output(0));
  mux_2206_nl <= MUX_s_1_2_2(mux_2205_nl, mux_2204_nl, fsm_output(4));
  nand_477_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2202_nl <= MUX_s_1_2_2(or_tmp_2562, nand_477_nl, fsm_output(0));
  or_2673_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2201_nl <= MUX_s_1_2_2(or_tmp_2558, or_2673_nl, fsm_output(0));
  mux_2203_nl <= MUX_s_1_2_2(mux_2202_nl, mux_2201_nl, fsm_output(4));
  mux_2207_nl <= MUX_s_1_2_2(mux_2206_nl, mux_2203_nl, fsm_output(6));
  or_4095_nl <= (fsm_output(2)) OR mux_2207_nl;
  mux_2215_nl <= MUX_s_1_2_2(nand_422_nl, or_4095_nl, fsm_output(5));
  vec_rsc_0_47_i_we_d_pff <= NOT(mux_2215_nl OR (fsm_output(1)));
  or_2714_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2713_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2228_nl <= MUX_s_1_2_2(or_2714_nl, or_2713_nl, fsm_output(0));
  or_2715_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2228_nl;
  or_2711_nl <= (NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(4
      DOWNTO 0)=STD_LOGIC_VECTOR'("01111")))) OR not_tmp_452;
  mux_2225_nl <= MUX_s_1_2_2(or_2711_nl, or_tmp_2567, fsm_output(0));
  nand_278_nl <= NOT(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("101111")) AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2224_nl <= MUX_s_1_2_2(nand_278_nl, or_tmp_2564, fsm_output(0));
  mux_2226_nl <= MUX_s_1_2_2(mux_2225_nl, mux_2224_nl, fsm_output(4));
  nand_402_nl <= NOT(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("101111")) AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2222_nl <= MUX_s_1_2_2(nand_402_nl, or_tmp_2562, fsm_output(0));
  or_2706_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101111")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2221_nl <= MUX_s_1_2_2(or_2706_nl, or_tmp_2558, fsm_output(0));
  mux_2223_nl <= MUX_s_1_2_2(mux_2222_nl, mux_2221_nl, fsm_output(4));
  mux_2227_nl <= MUX_s_1_2_2(mux_2226_nl, mux_2223_nl, fsm_output(6));
  mux_2229_nl <= MUX_s_1_2_2(or_2715_nl, mux_2227_nl, fsm_output(2));
  or_2704_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)) OR not_tmp_321;
  nand_281_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND and_763_cse);
  mux_2218_nl <= MUX_s_1_2_2(or_2704_nl, nand_281_nl, fsm_output(0));
  nand_282_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("10111"))
      AND COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
      (fsm_output(3)) AND (NOT (fsm_output(7))));
  nand_283_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2217_nl <= MUX_s_1_2_2(nand_282_nl, nand_283_nl, fsm_output(0));
  mux_2219_nl <= MUX_s_1_2_2(mux_2218_nl, mux_2217_nl, fsm_output(4));
  nor_907_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_908_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2216_nl <= MUX_s_1_2_2(nor_907_nl, nor_908_nl, fsm_output(0));
  nand_109_nl <= NOT((fsm_output(4)) AND mux_2216_nl);
  mux_2220_nl <= MUX_s_1_2_2(mux_2219_nl, nand_109_nl, fsm_output(6));
  or_2705_nl <= (fsm_output(2)) OR mux_2220_nl;
  mux_2230_nl <= MUX_s_1_2_2(mux_2229_nl, or_2705_nl, fsm_output(5));
  vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2230_nl) AND (fsm_output(1));
  nor_898_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR not_tmp_523);
  nor_899_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_2242_nl <= MUX_s_1_2_2(nor_898_nl, nor_899_nl, fsm_output(0));
  nor_900_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_901_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2241_nl <= MUX_s_1_2_2(nor_900_nl, nor_901_nl, fsm_output(0));
  mux_2243_nl <= MUX_s_1_2_2(mux_2242_nl, mux_2241_nl, fsm_output(4));
  nor_902_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_903_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2239_nl <= MUX_s_1_2_2(nor_902_nl, nor_903_nl, fsm_output(0));
  nor_904_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_905_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2238_nl <= MUX_s_1_2_2(nor_904_nl, nor_905_nl, fsm_output(0));
  mux_2240_nl <= MUX_s_1_2_2(mux_2239_nl, mux_2238_nl, fsm_output(4));
  mux_2244_nl <= MUX_s_1_2_2(mux_2243_nl, mux_2240_nl, fsm_output(6));
  nand_421_nl <= NOT((fsm_output(2)) AND mux_2244_nl);
  or_2725_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR not_tmp_522;
  mux_2235_nl <= MUX_s_1_2_2(or_tmp_2611, or_2725_nl, fsm_output(0));
  or_2722_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2234_nl <= MUX_s_1_2_2(or_tmp_2607, or_2722_nl, fsm_output(0));
  mux_2236_nl <= MUX_s_1_2_2(mux_2235_nl, mux_2234_nl, fsm_output(4));
  or_2719_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2232_nl <= MUX_s_1_2_2(or_tmp_2605, or_2719_nl, fsm_output(0));
  or_2716_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2231_nl <= MUX_s_1_2_2(or_tmp_2601, or_2716_nl, fsm_output(0));
  mux_2233_nl <= MUX_s_1_2_2(mux_2232_nl, mux_2231_nl, fsm_output(4));
  mux_2237_nl <= MUX_s_1_2_2(mux_2236_nl, mux_2233_nl, fsm_output(6));
  or_4094_nl <= (fsm_output(2)) OR mux_2237_nl;
  mux_2245_nl <= MUX_s_1_2_2(nand_421_nl, or_4094_nl, fsm_output(5));
  vec_rsc_0_48_i_we_d_pff <= NOT(mux_2245_nl OR (fsm_output(1)));
  or_2758_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2757_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2258_nl <= MUX_s_1_2_2(or_2758_nl, or_2757_nl, fsm_output(0));
  or_2759_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2258_nl;
  or_2755_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR not_tmp_522;
  mux_2255_nl <= MUX_s_1_2_2(or_2755_nl, or_tmp_2611, fsm_output(0));
  or_2753_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110000")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2254_nl <= MUX_s_1_2_2(or_2753_nl, or_tmp_2607, fsm_output(0));
  mux_2256_nl <= MUX_s_1_2_2(mux_2255_nl, mux_2254_nl, fsm_output(4));
  or_2752_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110000")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2252_nl <= MUX_s_1_2_2(or_2752_nl, or_tmp_2605, fsm_output(0));
  or_2750_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110000")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2251_nl <= MUX_s_1_2_2(or_2750_nl, or_tmp_2601, fsm_output(0));
  mux_2253_nl <= MUX_s_1_2_2(mux_2252_nl, mux_2251_nl, fsm_output(4));
  mux_2257_nl <= MUX_s_1_2_2(mux_2256_nl, mux_2253_nl, fsm_output(6));
  mux_2259_nl <= MUX_s_1_2_2(or_2759_nl, mux_2257_nl, fsm_output(2));
  or_2748_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2746_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR not_tmp_527;
  mux_2248_nl <= MUX_s_1_2_2(or_2748_nl, or_2746_nl, fsm_output(0));
  or_2744_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2743_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2247_nl <= MUX_s_1_2_2(or_2744_nl, or_2743_nl, fsm_output(0));
  mux_2249_nl <= MUX_s_1_2_2(mux_2248_nl, mux_2247_nl, fsm_output(4));
  nor_896_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_897_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2246_nl <= MUX_s_1_2_2(nor_896_nl, nor_897_nl, fsm_output(0));
  nand_111_nl <= NOT((fsm_output(4)) AND mux_2246_nl);
  mux_2250_nl <= MUX_s_1_2_2(mux_2249_nl, nand_111_nl, fsm_output(6));
  or_2749_nl <= (fsm_output(2)) OR mux_2250_nl;
  mux_2260_nl <= MUX_s_1_2_2(mux_2259_nl, or_2749_nl, fsm_output(5));
  vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2260_nl) AND (fsm_output(1));
  nor_887_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR not_tmp_523);
  nor_888_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_2272_nl <= MUX_s_1_2_2(nor_887_nl, nor_888_nl, fsm_output(0));
  nor_889_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_890_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2271_nl <= MUX_s_1_2_2(nor_889_nl, nor_890_nl, fsm_output(0));
  mux_2273_nl <= MUX_s_1_2_2(mux_2272_nl, mux_2271_nl, fsm_output(4));
  nor_891_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_892_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2269_nl <= MUX_s_1_2_2(nor_891_nl, nor_892_nl, fsm_output(0));
  nor_893_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_894_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2268_nl <= MUX_s_1_2_2(nor_893_nl, nor_894_nl, fsm_output(0));
  mux_2270_nl <= MUX_s_1_2_2(mux_2269_nl, mux_2268_nl, fsm_output(4));
  mux_2274_nl <= MUX_s_1_2_2(mux_2273_nl, mux_2270_nl, fsm_output(6));
  nand_420_nl <= NOT((fsm_output(2)) AND mux_2274_nl);
  or_2769_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR not_tmp_522;
  mux_2265_nl <= MUX_s_1_2_2(or_tmp_2655, or_2769_nl, fsm_output(0));
  or_2766_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2264_nl <= MUX_s_1_2_2(or_tmp_2651, or_2766_nl, fsm_output(0));
  mux_2266_nl <= MUX_s_1_2_2(mux_2265_nl, mux_2264_nl, fsm_output(4));
  or_2763_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2262_nl <= MUX_s_1_2_2(or_tmp_2649, or_2763_nl, fsm_output(0));
  or_2760_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2261_nl <= MUX_s_1_2_2(or_tmp_2645, or_2760_nl, fsm_output(0));
  mux_2263_nl <= MUX_s_1_2_2(mux_2262_nl, mux_2261_nl, fsm_output(4));
  mux_2267_nl <= MUX_s_1_2_2(mux_2266_nl, mux_2263_nl, fsm_output(6));
  or_4093_nl <= (fsm_output(2)) OR mux_2267_nl;
  mux_2275_nl <= MUX_s_1_2_2(nand_420_nl, or_4093_nl, fsm_output(5));
  vec_rsc_0_49_i_we_d_pff <= NOT(mux_2275_nl OR (fsm_output(1)));
  or_2802_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2801_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2288_nl <= MUX_s_1_2_2(or_2802_nl, or_2801_nl, fsm_output(0));
  or_2803_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2288_nl;
  or_2799_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR not_tmp_522;
  mux_2285_nl <= MUX_s_1_2_2(or_2799_nl, or_tmp_2655, fsm_output(0));
  or_2797_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110001")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2284_nl <= MUX_s_1_2_2(or_2797_nl, or_tmp_2651, fsm_output(0));
  mux_2286_nl <= MUX_s_1_2_2(mux_2285_nl, mux_2284_nl, fsm_output(4));
  or_2796_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110001")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2282_nl <= MUX_s_1_2_2(or_2796_nl, or_tmp_2649, fsm_output(0));
  or_2794_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110001")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2281_nl <= MUX_s_1_2_2(or_2794_nl, or_tmp_2645, fsm_output(0));
  mux_2283_nl <= MUX_s_1_2_2(mux_2282_nl, mux_2281_nl, fsm_output(4));
  mux_2287_nl <= MUX_s_1_2_2(mux_2286_nl, mux_2283_nl, fsm_output(6));
  mux_2289_nl <= MUX_s_1_2_2(or_2803_nl, mux_2287_nl, fsm_output(2));
  or_2792_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_2790_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR not_tmp_527;
  mux_2278_nl <= MUX_s_1_2_2(or_2792_nl, or_2790_nl, fsm_output(0));
  or_2788_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2787_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2277_nl <= MUX_s_1_2_2(or_2788_nl, or_2787_nl, fsm_output(0));
  mux_2279_nl <= MUX_s_1_2_2(mux_2278_nl, mux_2277_nl, fsm_output(4));
  nor_885_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_886_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2276_nl <= MUX_s_1_2_2(nor_885_nl, nor_886_nl, fsm_output(0));
  nand_113_nl <= NOT((fsm_output(4)) AND mux_2276_nl);
  mux_2280_nl <= MUX_s_1_2_2(mux_2279_nl, nand_113_nl, fsm_output(6));
  or_2793_nl <= (fsm_output(2)) OR mux_2280_nl;
  mux_2290_nl <= MUX_s_1_2_2(mux_2289_nl, or_2793_nl, fsm_output(5));
  vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2290_nl) AND (fsm_output(1));
  nor_876_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR not_tmp_523);
  nor_877_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR (NOT and_763_cse));
  mux_2302_nl <= MUX_s_1_2_2(nor_876_nl, nor_877_nl, fsm_output(0));
  nor_878_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_879_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2301_nl <= MUX_s_1_2_2(nor_878_nl, nor_879_nl, fsm_output(0));
  mux_2303_nl <= MUX_s_1_2_2(mux_2302_nl, mux_2301_nl, fsm_output(4));
  nor_880_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_881_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2299_nl <= MUX_s_1_2_2(nor_880_nl, nor_881_nl, fsm_output(0));
  nor_882_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_883_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2298_nl <= MUX_s_1_2_2(nor_882_nl, nor_883_nl, fsm_output(0));
  mux_2300_nl <= MUX_s_1_2_2(mux_2299_nl, mux_2298_nl, fsm_output(4));
  mux_2304_nl <= MUX_s_1_2_2(mux_2303_nl, mux_2300_nl, fsm_output(6));
  nand_419_nl <= NOT((fsm_output(2)) AND mux_2304_nl);
  or_2813_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR not_tmp_522;
  mux_2295_nl <= MUX_s_1_2_2(or_tmp_2699, or_2813_nl, fsm_output(0));
  or_2810_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2294_nl <= MUX_s_1_2_2(or_tmp_2695, or_2810_nl, fsm_output(0));
  mux_2296_nl <= MUX_s_1_2_2(mux_2295_nl, mux_2294_nl, fsm_output(4));
  or_2807_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2292_nl <= MUX_s_1_2_2(or_tmp_2693, or_2807_nl, fsm_output(0));
  or_2804_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2291_nl <= MUX_s_1_2_2(or_tmp_2689, or_2804_nl, fsm_output(0));
  mux_2293_nl <= MUX_s_1_2_2(mux_2292_nl, mux_2291_nl, fsm_output(4));
  mux_2297_nl <= MUX_s_1_2_2(mux_2296_nl, mux_2293_nl, fsm_output(6));
  or_4092_nl <= (fsm_output(2)) OR mux_2297_nl;
  mux_2305_nl <= MUX_s_1_2_2(nand_419_nl, or_4092_nl, fsm_output(5));
  vec_rsc_0_50_i_we_d_pff <= NOT(mux_2305_nl OR (fsm_output(1)));
  or_2846_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2845_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2318_nl <= MUX_s_1_2_2(or_2846_nl, or_2845_nl, fsm_output(0));
  or_2847_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2318_nl;
  or_2843_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR not_tmp_522;
  mux_2315_nl <= MUX_s_1_2_2(or_2843_nl, or_tmp_2699, fsm_output(0));
  or_2841_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110010")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2314_nl <= MUX_s_1_2_2(or_2841_nl, or_tmp_2695, fsm_output(0));
  mux_2316_nl <= MUX_s_1_2_2(mux_2315_nl, mux_2314_nl, fsm_output(4));
  or_2840_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110010")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2312_nl <= MUX_s_1_2_2(or_2840_nl, or_tmp_2693, fsm_output(0));
  or_2838_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110010")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2311_nl <= MUX_s_1_2_2(or_2838_nl, or_tmp_2689, fsm_output(0));
  mux_2313_nl <= MUX_s_1_2_2(mux_2312_nl, mux_2311_nl, fsm_output(4));
  mux_2317_nl <= MUX_s_1_2_2(mux_2316_nl, mux_2313_nl, fsm_output(6));
  mux_2319_nl <= MUX_s_1_2_2(or_2847_nl, mux_2317_nl, fsm_output(2));
  or_2836_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2834_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR not_tmp_527;
  mux_2308_nl <= MUX_s_1_2_2(or_2836_nl, or_2834_nl, fsm_output(0));
  or_2832_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2831_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2307_nl <= MUX_s_1_2_2(or_2832_nl, or_2831_nl, fsm_output(0));
  mux_2309_nl <= MUX_s_1_2_2(mux_2308_nl, mux_2307_nl, fsm_output(4));
  nor_874_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_875_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2306_nl <= MUX_s_1_2_2(nor_874_nl, nor_875_nl, fsm_output(0));
  nand_115_nl <= NOT((fsm_output(4)) AND mux_2306_nl);
  mux_2310_nl <= MUX_s_1_2_2(mux_2309_nl, nand_115_nl, fsm_output(6));
  or_2837_nl <= (fsm_output(2)) OR mux_2310_nl;
  mux_2320_nl <= MUX_s_1_2_2(mux_2319_nl, or_2837_nl, fsm_output(5));
  vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2320_nl) AND (fsm_output(1));
  nor_865_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR not_tmp_523);
  nor_866_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR not_tmp_330);
  mux_2332_nl <= MUX_s_1_2_2(nor_865_nl, nor_866_nl, fsm_output(0));
  nor_867_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_868_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2331_nl <= MUX_s_1_2_2(nor_867_nl, nor_868_nl, fsm_output(0));
  mux_2333_nl <= MUX_s_1_2_2(mux_2332_nl, mux_2331_nl, fsm_output(4));
  nor_869_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_870_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2329_nl <= MUX_s_1_2_2(nor_869_nl, nor_870_nl, fsm_output(0));
  nor_871_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_872_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2328_nl <= MUX_s_1_2_2(nor_871_nl, nor_872_nl, fsm_output(0));
  mux_2330_nl <= MUX_s_1_2_2(mux_2329_nl, mux_2328_nl, fsm_output(4));
  mux_2334_nl <= MUX_s_1_2_2(mux_2333_nl, mux_2330_nl, fsm_output(6));
  nand_418_nl <= NOT((fsm_output(2)) AND mux_2334_nl);
  or_2857_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR not_tmp_522;
  mux_2325_nl <= MUX_s_1_2_2(or_tmp_2743, or_2857_nl, fsm_output(0));
  or_2854_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2324_nl <= MUX_s_1_2_2(or_tmp_2739, or_2854_nl, fsm_output(0));
  mux_2326_nl <= MUX_s_1_2_2(mux_2325_nl, mux_2324_nl, fsm_output(4));
  or_2851_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2322_nl <= MUX_s_1_2_2(or_tmp_2737, or_2851_nl, fsm_output(0));
  or_2848_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2321_nl <= MUX_s_1_2_2(or_tmp_2733, or_2848_nl, fsm_output(0));
  mux_2323_nl <= MUX_s_1_2_2(mux_2322_nl, mux_2321_nl, fsm_output(4));
  mux_2327_nl <= MUX_s_1_2_2(mux_2326_nl, mux_2323_nl, fsm_output(6));
  or_4091_nl <= (fsm_output(2)) OR mux_2327_nl;
  mux_2335_nl <= MUX_s_1_2_2(nand_418_nl, or_4091_nl, fsm_output(5));
  vec_rsc_0_51_i_we_d_pff <= NOT(mux_2335_nl OR (fsm_output(1)));
  or_2890_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2889_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2348_nl <= MUX_s_1_2_2(or_2890_nl, or_2889_nl, fsm_output(0));
  or_2891_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2348_nl;
  or_2887_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR not_tmp_522;
  mux_2345_nl <= MUX_s_1_2_2(or_2887_nl, or_tmp_2743, fsm_output(0));
  or_2885_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110011")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2344_nl <= MUX_s_1_2_2(or_2885_nl, or_tmp_2739, fsm_output(0));
  mux_2346_nl <= MUX_s_1_2_2(mux_2345_nl, mux_2344_nl, fsm_output(4));
  or_2884_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110011")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2342_nl <= MUX_s_1_2_2(or_2884_nl, or_tmp_2737, fsm_output(0));
  or_2882_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110011")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2341_nl <= MUX_s_1_2_2(or_2882_nl, or_tmp_2733, fsm_output(0));
  mux_2343_nl <= MUX_s_1_2_2(mux_2342_nl, mux_2341_nl, fsm_output(4));
  mux_2347_nl <= MUX_s_1_2_2(mux_2346_nl, mux_2343_nl, fsm_output(6));
  mux_2349_nl <= MUX_s_1_2_2(or_2891_nl, mux_2347_nl, fsm_output(2));
  or_2880_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_2878_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR not_tmp_527;
  mux_2338_nl <= MUX_s_1_2_2(or_2880_nl, or_2878_nl, fsm_output(0));
  or_2876_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2875_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2337_nl <= MUX_s_1_2_2(or_2876_nl, or_2875_nl, fsm_output(0));
  mux_2339_nl <= MUX_s_1_2_2(mux_2338_nl, mux_2337_nl, fsm_output(4));
  nor_863_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_864_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2336_nl <= MUX_s_1_2_2(nor_863_nl, nor_864_nl, fsm_output(0));
  nand_117_nl <= NOT((fsm_output(4)) AND mux_2336_nl);
  mux_2340_nl <= MUX_s_1_2_2(mux_2339_nl, nand_117_nl, fsm_output(6));
  or_2881_nl <= (fsm_output(2)) OR mux_2340_nl;
  mux_2350_nl <= MUX_s_1_2_2(mux_2349_nl, or_2881_nl, fsm_output(5));
  vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2350_nl) AND (fsm_output(1));
  nor_854_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR not_tmp_523);
  nor_855_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_2362_nl <= MUX_s_1_2_2(nor_854_nl, nor_855_nl, fsm_output(0));
  nor_856_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_857_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2361_nl <= MUX_s_1_2_2(nor_856_nl, nor_857_nl, fsm_output(0));
  mux_2363_nl <= MUX_s_1_2_2(mux_2362_nl, mux_2361_nl, fsm_output(4));
  nor_858_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_859_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2359_nl <= MUX_s_1_2_2(nor_858_nl, nor_859_nl, fsm_output(0));
  nor_860_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_861_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2358_nl <= MUX_s_1_2_2(nor_860_nl, nor_861_nl, fsm_output(0));
  mux_2360_nl <= MUX_s_1_2_2(mux_2359_nl, mux_2358_nl, fsm_output(4));
  mux_2364_nl <= MUX_s_1_2_2(mux_2363_nl, mux_2360_nl, fsm_output(6));
  nand_417_nl <= NOT((fsm_output(2)) AND mux_2364_nl);
  or_2901_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR not_tmp_522;
  mux_2355_nl <= MUX_s_1_2_2(or_tmp_2787, or_2901_nl, fsm_output(0));
  or_2898_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2354_nl <= MUX_s_1_2_2(or_tmp_2783, or_2898_nl, fsm_output(0));
  mux_2356_nl <= MUX_s_1_2_2(mux_2355_nl, mux_2354_nl, fsm_output(4));
  or_2895_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2352_nl <= MUX_s_1_2_2(or_tmp_2781, or_2895_nl, fsm_output(0));
  or_2892_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2351_nl <= MUX_s_1_2_2(or_tmp_2777, or_2892_nl, fsm_output(0));
  mux_2353_nl <= MUX_s_1_2_2(mux_2352_nl, mux_2351_nl, fsm_output(4));
  mux_2357_nl <= MUX_s_1_2_2(mux_2356_nl, mux_2353_nl, fsm_output(6));
  or_4090_nl <= (fsm_output(2)) OR mux_2357_nl;
  mux_2365_nl <= MUX_s_1_2_2(nand_417_nl, or_4090_nl, fsm_output(5));
  vec_rsc_0_52_i_we_d_pff <= NOT(mux_2365_nl OR (fsm_output(1)));
  or_2934_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2933_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2378_nl <= MUX_s_1_2_2(or_2934_nl, or_2933_nl, fsm_output(0));
  or_2935_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2378_nl;
  or_2931_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR not_tmp_522;
  mux_2375_nl <= MUX_s_1_2_2(or_2931_nl, or_tmp_2787, fsm_output(0));
  or_2929_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110100")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2374_nl <= MUX_s_1_2_2(or_2929_nl, or_tmp_2783, fsm_output(0));
  mux_2376_nl <= MUX_s_1_2_2(mux_2375_nl, mux_2374_nl, fsm_output(4));
  or_2928_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110100")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2372_nl <= MUX_s_1_2_2(or_2928_nl, or_tmp_2781, fsm_output(0));
  or_2926_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110100")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2371_nl <= MUX_s_1_2_2(or_2926_nl, or_tmp_2777, fsm_output(0));
  mux_2373_nl <= MUX_s_1_2_2(mux_2372_nl, mux_2371_nl, fsm_output(4));
  mux_2377_nl <= MUX_s_1_2_2(mux_2376_nl, mux_2373_nl, fsm_output(6));
  mux_2379_nl <= MUX_s_1_2_2(or_2935_nl, mux_2377_nl, fsm_output(2));
  or_2924_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_2922_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR not_tmp_544;
  mux_2368_nl <= MUX_s_1_2_2(or_2924_nl, or_2922_nl, fsm_output(0));
  or_2920_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2919_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2367_nl <= MUX_s_1_2_2(or_2920_nl, or_2919_nl, fsm_output(0));
  mux_2369_nl <= MUX_s_1_2_2(mux_2368_nl, mux_2367_nl, fsm_output(4));
  nor_852_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_853_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2366_nl <= MUX_s_1_2_2(nor_852_nl, nor_853_nl, fsm_output(0));
  nand_119_nl <= NOT((fsm_output(4)) AND mux_2366_nl);
  mux_2370_nl <= MUX_s_1_2_2(mux_2369_nl, nand_119_nl, fsm_output(6));
  or_2925_nl <= (fsm_output(2)) OR mux_2370_nl;
  mux_2380_nl <= MUX_s_1_2_2(mux_2379_nl, or_2925_nl, fsm_output(5));
  vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2380_nl) AND (fsm_output(1));
  nor_843_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR not_tmp_523);
  nor_844_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_2392_nl <= MUX_s_1_2_2(nor_843_nl, nor_844_nl, fsm_output(0));
  nor_845_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_846_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2391_nl <= MUX_s_1_2_2(nor_845_nl, nor_846_nl, fsm_output(0));
  mux_2393_nl <= MUX_s_1_2_2(mux_2392_nl, mux_2391_nl, fsm_output(4));
  nor_847_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_848_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2389_nl <= MUX_s_1_2_2(nor_847_nl, nor_848_nl, fsm_output(0));
  nor_849_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_850_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2388_nl <= MUX_s_1_2_2(nor_849_nl, nor_850_nl, fsm_output(0));
  mux_2390_nl <= MUX_s_1_2_2(mux_2389_nl, mux_2388_nl, fsm_output(4));
  mux_2394_nl <= MUX_s_1_2_2(mux_2393_nl, mux_2390_nl, fsm_output(6));
  nand_416_nl <= NOT((fsm_output(2)) AND mux_2394_nl);
  or_2945_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR not_tmp_522;
  mux_2385_nl <= MUX_s_1_2_2(or_tmp_2831, or_2945_nl, fsm_output(0));
  or_2942_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2384_nl <= MUX_s_1_2_2(or_tmp_2827, or_2942_nl, fsm_output(0));
  mux_2386_nl <= MUX_s_1_2_2(mux_2385_nl, mux_2384_nl, fsm_output(4));
  or_2939_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2382_nl <= MUX_s_1_2_2(or_tmp_2825, or_2939_nl, fsm_output(0));
  or_2936_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2381_nl <= MUX_s_1_2_2(or_tmp_2821, or_2936_nl, fsm_output(0));
  mux_2383_nl <= MUX_s_1_2_2(mux_2382_nl, mux_2381_nl, fsm_output(4));
  mux_2387_nl <= MUX_s_1_2_2(mux_2386_nl, mux_2383_nl, fsm_output(6));
  or_4089_nl <= (fsm_output(2)) OR mux_2387_nl;
  mux_2395_nl <= MUX_s_1_2_2(nand_416_nl, or_4089_nl, fsm_output(5));
  vec_rsc_0_53_i_we_d_pff <= NOT(mux_2395_nl OR (fsm_output(1)));
  or_2978_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_2977_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2408_nl <= MUX_s_1_2_2(or_2978_nl, or_2977_nl, fsm_output(0));
  or_2979_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2408_nl;
  or_2975_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR not_tmp_522;
  mux_2405_nl <= MUX_s_1_2_2(or_2975_nl, or_tmp_2831, fsm_output(0));
  or_2973_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110101")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2404_nl <= MUX_s_1_2_2(or_2973_nl, or_tmp_2827, fsm_output(0));
  mux_2406_nl <= MUX_s_1_2_2(mux_2405_nl, mux_2404_nl, fsm_output(4));
  or_2972_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110101")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2402_nl <= MUX_s_1_2_2(or_2972_nl, or_tmp_2825, fsm_output(0));
  or_2970_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110101")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2401_nl <= MUX_s_1_2_2(or_2970_nl, or_tmp_2821, fsm_output(0));
  mux_2403_nl <= MUX_s_1_2_2(mux_2402_nl, mux_2401_nl, fsm_output(4));
  mux_2407_nl <= MUX_s_1_2_2(mux_2406_nl, mux_2403_nl, fsm_output(6));
  mux_2409_nl <= MUX_s_1_2_2(or_2979_nl, mux_2407_nl, fsm_output(2));
  or_2968_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_2966_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR not_tmp_549;
  mux_2398_nl <= MUX_s_1_2_2(or_2968_nl, or_2966_nl, fsm_output(0));
  or_2964_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2963_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2397_nl <= MUX_s_1_2_2(or_2964_nl, or_2963_nl, fsm_output(0));
  mux_2399_nl <= MUX_s_1_2_2(mux_2398_nl, mux_2397_nl, fsm_output(4));
  nor_841_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_842_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2396_nl <= MUX_s_1_2_2(nor_841_nl, nor_842_nl, fsm_output(0));
  nand_121_nl <= NOT((fsm_output(4)) AND mux_2396_nl);
  mux_2400_nl <= MUX_s_1_2_2(mux_2399_nl, nand_121_nl, fsm_output(6));
  or_2969_nl <= (fsm_output(2)) OR mux_2400_nl;
  mux_2410_nl <= MUX_s_1_2_2(mux_2409_nl, or_2969_nl, fsm_output(5));
  vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2410_nl) AND (fsm_output(1));
  nor_833_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR not_tmp_523);
  and_567_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND and_763_cse;
  mux_2422_nl <= MUX_s_1_2_2(nor_833_nl, and_567_nl, fsm_output(0));
  nor_834_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_835_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2421_nl <= MUX_s_1_2_2(nor_834_nl, nor_835_nl, fsm_output(0));
  mux_2423_nl <= MUX_s_1_2_2(mux_2422_nl, mux_2421_nl, fsm_output(4));
  nor_836_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_837_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2419_nl <= MUX_s_1_2_2(nor_836_nl, nor_837_nl, fsm_output(0));
  nor_838_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_839_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2418_nl <= MUX_s_1_2_2(nor_838_nl, nor_839_nl, fsm_output(0));
  mux_2420_nl <= MUX_s_1_2_2(mux_2419_nl, mux_2418_nl, fsm_output(4));
  mux_2424_nl <= MUX_s_1_2_2(mux_2423_nl, mux_2420_nl, fsm_output(6));
  nand_415_nl <= NOT((fsm_output(2)) AND mux_2424_nl);
  or_2989_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR not_tmp_522;
  mux_2415_nl <= MUX_s_1_2_2(or_tmp_2875, or_2989_nl, fsm_output(0));
  or_2986_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2414_nl <= MUX_s_1_2_2(or_tmp_2871, or_2986_nl, fsm_output(0));
  mux_2416_nl <= MUX_s_1_2_2(mux_2415_nl, mux_2414_nl, fsm_output(4));
  or_2983_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2412_nl <= MUX_s_1_2_2(or_tmp_2869, or_2983_nl, fsm_output(0));
  or_2980_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2411_nl <= MUX_s_1_2_2(or_tmp_2865, or_2980_nl, fsm_output(0));
  mux_2413_nl <= MUX_s_1_2_2(mux_2412_nl, mux_2411_nl, fsm_output(4));
  mux_2417_nl <= MUX_s_1_2_2(mux_2416_nl, mux_2413_nl, fsm_output(6));
  or_4088_nl <= (fsm_output(2)) OR mux_2417_nl;
  mux_2425_nl <= MUX_s_1_2_2(nand_415_nl, or_4088_nl, fsm_output(5));
  vec_rsc_0_54_i_we_d_pff <= NOT(mux_2425_nl OR (fsm_output(1)));
  or_3022_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3021_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2438_nl <= MUX_s_1_2_2(or_3022_nl, or_3021_nl, fsm_output(0));
  or_3023_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2438_nl;
  or_3019_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR not_tmp_522;
  mux_2435_nl <= MUX_s_1_2_2(or_3019_nl, or_tmp_2875, fsm_output(0));
  or_3017_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110110")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2434_nl <= MUX_s_1_2_2(or_3017_nl, or_tmp_2871, fsm_output(0));
  mux_2436_nl <= MUX_s_1_2_2(mux_2435_nl, mux_2434_nl, fsm_output(4));
  or_3016_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110110")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2432_nl <= MUX_s_1_2_2(or_3016_nl, or_tmp_2869, fsm_output(0));
  or_3014_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110110")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2431_nl <= MUX_s_1_2_2(or_3014_nl, or_tmp_2865, fsm_output(0));
  mux_2433_nl <= MUX_s_1_2_2(mux_2432_nl, mux_2431_nl, fsm_output(4));
  mux_2437_nl <= MUX_s_1_2_2(mux_2436_nl, mux_2433_nl, fsm_output(6));
  mux_2439_nl <= MUX_s_1_2_2(or_3023_nl, mux_2437_nl, fsm_output(2));
  nand_271_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND and_763_cse);
  or_3010_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR not_tmp_544;
  mux_2428_nl <= MUX_s_1_2_2(nand_271_nl, or_3010_nl, fsm_output(0));
  or_3008_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_3007_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2427_nl <= MUX_s_1_2_2(or_3008_nl, or_3007_nl, fsm_output(0));
  mux_2429_nl <= MUX_s_1_2_2(mux_2428_nl, mux_2427_nl, fsm_output(4));
  nor_831_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_832_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2426_nl <= MUX_s_1_2_2(nor_831_nl, nor_832_nl, fsm_output(0));
  nand_123_nl <= NOT((fsm_output(4)) AND mux_2426_nl);
  mux_2430_nl <= MUX_s_1_2_2(mux_2429_nl, nand_123_nl, fsm_output(6));
  or_3013_nl <= (fsm_output(2)) OR mux_2430_nl;
  mux_2440_nl <= MUX_s_1_2_2(mux_2439_nl, or_3013_nl, fsm_output(5));
  vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2440_nl) AND (fsm_output(1));
  nor_824_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))))
      OR not_tmp_523);
  nor_825_nl <= NOT((NOT (COMP_LOOP_acc_13_psp_sva(3))) OR (COMP_LOOP_acc_13_psp_sva(1))
      OR not_tmp_414);
  mux_2452_nl <= MUX_s_1_2_2(nor_824_nl, nor_825_nl, fsm_output(0));
  and_564_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_565_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  mux_2451_nl <= MUX_s_1_2_2(and_564_nl, and_565_nl, fsm_output(0));
  mux_2453_nl <= MUX_s_1_2_2(mux_2452_nl, mux_2451_nl, fsm_output(4));
  and_813_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7));
  and_820_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT (fsm_output(3))) AND (fsm_output(7));
  mux_2449_nl <= MUX_s_1_2_2(and_813_nl, and_820_nl, fsm_output(0));
  nor_828_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_829_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2448_nl <= MUX_s_1_2_2(nor_828_nl, nor_829_nl, fsm_output(0));
  mux_2450_nl <= MUX_s_1_2_2(mux_2449_nl, mux_2448_nl, fsm_output(4));
  mux_2454_nl <= MUX_s_1_2_2(mux_2453_nl, mux_2450_nl, fsm_output(6));
  nand_414_nl <= NOT((fsm_output(2)) AND mux_2454_nl);
  or_3033_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))))
      OR not_tmp_522;
  mux_2445_nl <= MUX_s_1_2_2(or_tmp_2919, or_3033_nl, fsm_output(0));
  nand_267_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2444_nl <= MUX_s_1_2_2(or_tmp_2915, nand_267_nl, fsm_output(0));
  mux_2446_nl <= MUX_s_1_2_2(mux_2445_nl, mux_2444_nl, fsm_output(4));
  nand_476_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2442_nl <= MUX_s_1_2_2(or_tmp_2913, nand_476_nl, fsm_output(0));
  or_3024_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2441_nl <= MUX_s_1_2_2(or_tmp_2909, or_3024_nl, fsm_output(0));
  mux_2443_nl <= MUX_s_1_2_2(mux_2442_nl, mux_2441_nl, fsm_output(4));
  mux_2447_nl <= MUX_s_1_2_2(mux_2446_nl, mux_2443_nl, fsm_output(6));
  or_4087_nl <= (fsm_output(2)) OR mux_2447_nl;
  mux_2455_nl <= MUX_s_1_2_2(nand_414_nl, or_4087_nl, fsm_output(5));
  vec_rsc_0_55_i_we_d_pff <= NOT(mux_2455_nl OR (fsm_output(1)));
  or_3066_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3065_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2468_nl <= MUX_s_1_2_2(or_3066_nl, or_3065_nl, fsm_output(0));
  or_3067_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2468_nl;
  or_3063_nl <= (NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0111")))) OR not_tmp_522;
  mux_2465_nl <= MUX_s_1_2_2(or_3063_nl, or_tmp_2919, fsm_output(0));
  nand_258_nl <= NOT(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("110111")) AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2464_nl <= MUX_s_1_2_2(nand_258_nl, or_tmp_2915, fsm_output(0));
  mux_2466_nl <= MUX_s_1_2_2(mux_2465_nl, mux_2464_nl, fsm_output(4));
  nand_400_nl <= NOT(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("110111")) AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2462_nl <= MUX_s_1_2_2(nand_400_nl, or_tmp_2913, fsm_output(0));
  or_3058_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110111")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2461_nl <= MUX_s_1_2_2(or_3058_nl, or_tmp_2909, fsm_output(0));
  mux_2463_nl <= MUX_s_1_2_2(mux_2462_nl, mux_2461_nl, fsm_output(4));
  mux_2467_nl <= MUX_s_1_2_2(mux_2466_nl, mux_2463_nl, fsm_output(6));
  mux_2469_nl <= MUX_s_1_2_2(or_3067_nl, mux_2467_nl, fsm_output(2));
  or_3056_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)) OR not_tmp_321;
  or_3054_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      OR not_tmp_549;
  mux_2458_nl <= MUX_s_1_2_2(or_3056_nl, or_3054_nl, fsm_output(0));
  nand_261_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11011"))
      AND COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
      (fsm_output(3)) AND (NOT (fsm_output(7))));
  nand_262_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2457_nl <= MUX_s_1_2_2(nand_261_nl, nand_262_nl, fsm_output(0));
  mux_2459_nl <= MUX_s_1_2_2(mux_2458_nl, mux_2457_nl, fsm_output(4));
  nor_822_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_823_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110111"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2456_nl <= MUX_s_1_2_2(nor_822_nl, nor_823_nl, fsm_output(0));
  nand_125_nl <= NOT((fsm_output(4)) AND mux_2456_nl);
  mux_2460_nl <= MUX_s_1_2_2(mux_2459_nl, nand_125_nl, fsm_output(6));
  or_3057_nl <= (fsm_output(2)) OR mux_2460_nl;
  mux_2470_nl <= MUX_s_1_2_2(mux_2469_nl, or_3057_nl, fsm_output(5));
  vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2470_nl) AND (fsm_output(1));
  nor_813_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR not_tmp_560);
  nor_814_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_763_cse));
  mux_2482_nl <= MUX_s_1_2_2(nor_813_nl, nor_814_nl, fsm_output(0));
  nor_815_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_816_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2481_nl <= MUX_s_1_2_2(nor_815_nl, nor_816_nl, fsm_output(0));
  mux_2483_nl <= MUX_s_1_2_2(mux_2482_nl, mux_2481_nl, fsm_output(4));
  nor_817_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_818_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2479_nl <= MUX_s_1_2_2(nor_817_nl, nor_818_nl, fsm_output(0));
  nor_819_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_820_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2478_nl <= MUX_s_1_2_2(nor_819_nl, nor_820_nl, fsm_output(0));
  mux_2480_nl <= MUX_s_1_2_2(mux_2479_nl, mux_2478_nl, fsm_output(4));
  mux_2484_nl <= MUX_s_1_2_2(mux_2483_nl, mux_2480_nl, fsm_output(6));
  nand_413_nl <= NOT((fsm_output(2)) AND mux_2484_nl);
  or_3077_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR not_tmp_559;
  mux_2475_nl <= MUX_s_1_2_2(or_tmp_2963, or_3077_nl, fsm_output(0));
  or_3074_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2474_nl <= MUX_s_1_2_2(or_tmp_2959, or_3074_nl, fsm_output(0));
  mux_2476_nl <= MUX_s_1_2_2(mux_2475_nl, mux_2474_nl, fsm_output(4));
  or_3071_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2472_nl <= MUX_s_1_2_2(or_tmp_2957, or_3071_nl, fsm_output(0));
  or_3068_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2471_nl <= MUX_s_1_2_2(or_tmp_2953, or_3068_nl, fsm_output(0));
  mux_2473_nl <= MUX_s_1_2_2(mux_2472_nl, mux_2471_nl, fsm_output(4));
  mux_2477_nl <= MUX_s_1_2_2(mux_2476_nl, mux_2473_nl, fsm_output(6));
  or_4086_nl <= (fsm_output(2)) OR mux_2477_nl;
  mux_2485_nl <= MUX_s_1_2_2(nand_413_nl, or_4086_nl, fsm_output(5));
  vec_rsc_0_56_i_we_d_pff <= NOT(mux_2485_nl OR (fsm_output(1)));
  or_3110_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3109_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2498_nl <= MUX_s_1_2_2(or_3110_nl, or_3109_nl, fsm_output(0));
  or_3111_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2498_nl;
  or_3107_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR not_tmp_559;
  mux_2495_nl <= MUX_s_1_2_2(or_3107_nl, or_tmp_2963, fsm_output(0));
  or_3105_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111000")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2494_nl <= MUX_s_1_2_2(or_3105_nl, or_tmp_2959, fsm_output(0));
  mux_2496_nl <= MUX_s_1_2_2(mux_2495_nl, mux_2494_nl, fsm_output(4));
  or_3104_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111000")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2492_nl <= MUX_s_1_2_2(or_3104_nl, or_tmp_2957, fsm_output(0));
  or_3102_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111000")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2491_nl <= MUX_s_1_2_2(or_3102_nl, or_tmp_2953, fsm_output(0));
  mux_2493_nl <= MUX_s_1_2_2(mux_2492_nl, mux_2491_nl, fsm_output(4));
  mux_2497_nl <= MUX_s_1_2_2(mux_2496_nl, mux_2493_nl, fsm_output(6));
  mux_2499_nl <= MUX_s_1_2_2(or_3111_nl, mux_2497_nl, fsm_output(2));
  or_3100_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT and_763_cse);
  or_3098_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR not_tmp_527;
  mux_2488_nl <= MUX_s_1_2_2(or_3100_nl, or_3098_nl, fsm_output(0));
  or_3096_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_3095_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2487_nl <= MUX_s_1_2_2(or_3096_nl, or_3095_nl, fsm_output(0));
  mux_2489_nl <= MUX_s_1_2_2(mux_2488_nl, mux_2487_nl, fsm_output(4));
  nor_811_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_812_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2486_nl <= MUX_s_1_2_2(nor_811_nl, nor_812_nl, fsm_output(0));
  nand_127_nl <= NOT((fsm_output(4)) AND mux_2486_nl);
  mux_2490_nl <= MUX_s_1_2_2(mux_2489_nl, nand_127_nl, fsm_output(6));
  or_3101_nl <= (fsm_output(2)) OR mux_2490_nl;
  mux_2500_nl <= MUX_s_1_2_2(mux_2499_nl, or_3101_nl, fsm_output(5));
  vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2500_nl) AND (fsm_output(1));
  nor_802_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR not_tmp_560);
  nor_803_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(1)) OR not_tmp_321);
  mux_2512_nl <= MUX_s_1_2_2(nor_802_nl, nor_803_nl, fsm_output(0));
  nor_804_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_805_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2511_nl <= MUX_s_1_2_2(nor_804_nl, nor_805_nl, fsm_output(0));
  mux_2513_nl <= MUX_s_1_2_2(mux_2512_nl, mux_2511_nl, fsm_output(4));
  nor_806_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_807_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2509_nl <= MUX_s_1_2_2(nor_806_nl, nor_807_nl, fsm_output(0));
  nor_808_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_809_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2508_nl <= MUX_s_1_2_2(nor_808_nl, nor_809_nl, fsm_output(0));
  mux_2510_nl <= MUX_s_1_2_2(mux_2509_nl, mux_2508_nl, fsm_output(4));
  mux_2514_nl <= MUX_s_1_2_2(mux_2513_nl, mux_2510_nl, fsm_output(6));
  nand_412_nl <= NOT((fsm_output(2)) AND mux_2514_nl);
  or_3121_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_565;
  mux_2505_nl <= MUX_s_1_2_2(or_tmp_3007, or_3121_nl, fsm_output(0));
  or_3118_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2504_nl <= MUX_s_1_2_2(or_tmp_3003, or_3118_nl, fsm_output(0));
  mux_2506_nl <= MUX_s_1_2_2(mux_2505_nl, mux_2504_nl, fsm_output(4));
  or_3115_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2502_nl <= MUX_s_1_2_2(or_tmp_3001, or_3115_nl, fsm_output(0));
  or_3112_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2501_nl <= MUX_s_1_2_2(or_tmp_2997, or_3112_nl, fsm_output(0));
  mux_2503_nl <= MUX_s_1_2_2(mux_2502_nl, mux_2501_nl, fsm_output(4));
  mux_2507_nl <= MUX_s_1_2_2(mux_2506_nl, mux_2503_nl, fsm_output(6));
  or_4085_nl <= (fsm_output(2)) OR mux_2507_nl;
  mux_2515_nl <= MUX_s_1_2_2(nand_412_nl, or_4085_nl, fsm_output(5));
  vec_rsc_0_57_i_we_d_pff <= NOT(mux_2515_nl OR (fsm_output(1)));
  or_3154_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3153_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2528_nl <= MUX_s_1_2_2(or_3154_nl, or_3153_nl, fsm_output(0));
  or_3155_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2528_nl;
  or_3151_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_565;
  mux_2525_nl <= MUX_s_1_2_2(or_3151_nl, or_tmp_3007, fsm_output(0));
  or_3149_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111001")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2524_nl <= MUX_s_1_2_2(or_3149_nl, or_tmp_3003, fsm_output(0));
  mux_2526_nl <= MUX_s_1_2_2(mux_2525_nl, mux_2524_nl, fsm_output(4));
  or_3148_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111001")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2522_nl <= MUX_s_1_2_2(or_3148_nl, or_tmp_3001, fsm_output(0));
  or_3146_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111001")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2521_nl <= MUX_s_1_2_2(or_3146_nl, or_tmp_2997, fsm_output(0));
  mux_2523_nl <= MUX_s_1_2_2(mux_2522_nl, mux_2521_nl, fsm_output(4));
  mux_2527_nl <= MUX_s_1_2_2(mux_2526_nl, mux_2523_nl, fsm_output(6));
  mux_2529_nl <= MUX_s_1_2_2(or_3155_nl, mux_2527_nl, fsm_output(2));
  or_3144_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm) OR not_tmp_321;
  or_3142_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR not_tmp_527;
  mux_2518_nl <= MUX_s_1_2_2(or_3144_nl, or_3142_nl, fsm_output(0));
  or_3140_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_3139_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2517_nl <= MUX_s_1_2_2(or_3140_nl, or_3139_nl, fsm_output(0));
  mux_2519_nl <= MUX_s_1_2_2(mux_2518_nl, mux_2517_nl, fsm_output(4));
  nor_800_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_801_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2516_nl <= MUX_s_1_2_2(nor_800_nl, nor_801_nl, fsm_output(0));
  nand_129_nl <= NOT((fsm_output(4)) AND mux_2516_nl);
  mux_2520_nl <= MUX_s_1_2_2(mux_2519_nl, nand_129_nl, fsm_output(6));
  or_3145_nl <= (fsm_output(2)) OR mux_2520_nl;
  mux_2530_nl <= MUX_s_1_2_2(mux_2529_nl, or_3145_nl, fsm_output(5));
  vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2530_nl) AND (fsm_output(1));
  nor_792_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR not_tmp_570);
  and_560_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND and_763_cse;
  mux_2542_nl <= MUX_s_1_2_2(nor_792_nl, and_560_nl, fsm_output(0));
  nor_793_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_794_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2541_nl <= MUX_s_1_2_2(nor_793_nl, nor_794_nl, fsm_output(0));
  mux_2543_nl <= MUX_s_1_2_2(mux_2542_nl, mux_2541_nl, fsm_output(4));
  nor_795_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_796_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2539_nl <= MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output(0));
  nor_797_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_798_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2538_nl <= MUX_s_1_2_2(nor_797_nl, nor_798_nl, fsm_output(0));
  mux_2540_nl <= MUX_s_1_2_2(mux_2539_nl, mux_2538_nl, fsm_output(4));
  mux_2544_nl <= MUX_s_1_2_2(mux_2543_nl, mux_2540_nl, fsm_output(6));
  nand_411_nl <= NOT((fsm_output(2)) AND mux_2544_nl);
  or_3165_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR not_tmp_559;
  mux_2535_nl <= MUX_s_1_2_2(or_tmp_3051, or_3165_nl, fsm_output(0));
  or_3162_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2534_nl <= MUX_s_1_2_2(or_tmp_3047, or_3162_nl, fsm_output(0));
  mux_2536_nl <= MUX_s_1_2_2(mux_2535_nl, mux_2534_nl, fsm_output(4));
  or_3159_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2532_nl <= MUX_s_1_2_2(or_tmp_3045, or_3159_nl, fsm_output(0));
  or_3156_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2531_nl <= MUX_s_1_2_2(or_tmp_3041, or_3156_nl, fsm_output(0));
  mux_2533_nl <= MUX_s_1_2_2(mux_2532_nl, mux_2531_nl, fsm_output(4));
  mux_2537_nl <= MUX_s_1_2_2(mux_2536_nl, mux_2533_nl, fsm_output(6));
  or_4084_nl <= (fsm_output(2)) OR mux_2537_nl;
  mux_2545_nl <= MUX_s_1_2_2(nand_411_nl, or_4084_nl, fsm_output(5));
  vec_rsc_0_58_i_we_d_pff <= NOT(mux_2545_nl OR (fsm_output(1)));
  or_3198_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3197_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2558_nl <= MUX_s_1_2_2(or_3198_nl, or_3197_nl, fsm_output(0));
  or_3199_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2558_nl;
  or_3195_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR not_tmp_559;
  mux_2555_nl <= MUX_s_1_2_2(or_3195_nl, or_tmp_3051, fsm_output(0));
  or_3193_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111010")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2554_nl <= MUX_s_1_2_2(or_3193_nl, or_tmp_3047, fsm_output(0));
  mux_2556_nl <= MUX_s_1_2_2(mux_2555_nl, mux_2554_nl, fsm_output(4));
  or_3192_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111010")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2552_nl <= MUX_s_1_2_2(or_3192_nl, or_tmp_3045, fsm_output(0));
  or_3190_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111010")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2551_nl <= MUX_s_1_2_2(or_3190_nl, or_tmp_3041, fsm_output(0));
  mux_2553_nl <= MUX_s_1_2_2(mux_2552_nl, mux_2551_nl, fsm_output(4));
  mux_2557_nl <= MUX_s_1_2_2(mux_2556_nl, mux_2553_nl, fsm_output(6));
  mux_2559_nl <= MUX_s_1_2_2(or_3199_nl, mux_2557_nl, fsm_output(2));
  nand_252_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND and_763_cse);
  or_3186_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR not_tmp_527;
  mux_2548_nl <= MUX_s_1_2_2(nand_252_nl, or_3186_nl, fsm_output(0));
  or_3184_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_3183_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2547_nl <= MUX_s_1_2_2(or_3184_nl, or_3183_nl, fsm_output(0));
  mux_2549_nl <= MUX_s_1_2_2(mux_2548_nl, mux_2547_nl, fsm_output(4));
  nor_790_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_791_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2546_nl <= MUX_s_1_2_2(nor_790_nl, nor_791_nl, fsm_output(0));
  nand_131_nl <= NOT((fsm_output(4)) AND mux_2546_nl);
  mux_2550_nl <= MUX_s_1_2_2(mux_2549_nl, nand_131_nl, fsm_output(6));
  or_3189_nl <= (fsm_output(2)) OR mux_2550_nl;
  mux_2560_nl <= MUX_s_1_2_2(mux_2559_nl, or_3189_nl, fsm_output(5));
  vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2560_nl) AND (fsm_output(1));
  nor_783_nl <= NOT((NOT (COMP_LOOP_acc_10_cse_10_1_5_sva(0))) OR (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      OR not_tmp_570);
  nor_784_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))))
      OR not_tmp_330);
  mux_2572_nl <= MUX_s_1_2_2(nor_783_nl, nor_784_nl, fsm_output(0));
  and_557_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_558_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  mux_2571_nl <= MUX_s_1_2_2(and_557_nl, and_558_nl, fsm_output(0));
  mux_2573_nl <= MUX_s_1_2_2(mux_2572_nl, mux_2571_nl, fsm_output(4));
  and_814_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7));
  and_821_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT (fsm_output(3))) AND (fsm_output(7));
  mux_2569_nl <= MUX_s_1_2_2(and_814_nl, and_821_nl, fsm_output(0));
  nor_787_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_788_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2568_nl <= MUX_s_1_2_2(nor_787_nl, nor_788_nl, fsm_output(0));
  mux_2570_nl <= MUX_s_1_2_2(mux_2569_nl, mux_2568_nl, fsm_output(4));
  mux_2574_nl <= MUX_s_1_2_2(mux_2573_nl, mux_2570_nl, fsm_output(6));
  nand_410_nl <= NOT((fsm_output(2)) AND mux_2574_nl);
  or_3208_nl <= (COMP_LOOP_acc_1_cse_6_sva(2)) OR not_tmp_575;
  mux_2565_nl <= MUX_s_1_2_2(or_tmp_3094, or_3208_nl, fsm_output(0));
  nand_247_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2564_nl <= MUX_s_1_2_2(or_tmp_3091, nand_247_nl, fsm_output(0));
  mux_2566_nl <= MUX_s_1_2_2(mux_2565_nl, mux_2564_nl, fsm_output(4));
  nand_475_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2562_nl <= MUX_s_1_2_2(or_tmp_3089, nand_475_nl, fsm_output(0));
  or_3200_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2561_nl <= MUX_s_1_2_2(or_tmp_3085, or_3200_nl, fsm_output(0));
  mux_2563_nl <= MUX_s_1_2_2(mux_2562_nl, mux_2561_nl, fsm_output(4));
  mux_2567_nl <= MUX_s_1_2_2(mux_2566_nl, mux_2563_nl, fsm_output(6));
  or_4083_nl <= (fsm_output(2)) OR mux_2567_nl;
  mux_2575_nl <= MUX_s_1_2_2(nand_410_nl, or_4083_nl, fsm_output(5));
  vec_rsc_0_59_i_we_d_pff <= NOT(mux_2575_nl OR (fsm_output(1)));
  or_3241_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3240_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2588_nl <= MUX_s_1_2_2(or_3241_nl, or_3240_nl, fsm_output(0));
  or_3242_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2588_nl;
  or_3238_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR (COMP_LOOP_acc_1_cse_6_sva(2))
      OR not_tmp_575;
  mux_2585_nl <= MUX_s_1_2_2(or_3238_nl, or_tmp_3094, fsm_output(0));
  nand_238_nl <= NOT(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111011")) AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2584_nl <= MUX_s_1_2_2(nand_238_nl, or_tmp_3091, fsm_output(0));
  mux_2586_nl <= MUX_s_1_2_2(mux_2585_nl, mux_2584_nl, fsm_output(4));
  nand_398_nl <= NOT(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111011")) AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2582_nl <= MUX_s_1_2_2(nand_398_nl, or_tmp_3089, fsm_output(0));
  or_3233_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111011")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2581_nl <= MUX_s_1_2_2(or_3233_nl, or_tmp_3085, fsm_output(0));
  mux_2583_nl <= MUX_s_1_2_2(mux_2582_nl, mux_2581_nl, fsm_output(4));
  mux_2587_nl <= MUX_s_1_2_2(mux_2586_nl, mux_2583_nl, fsm_output(6));
  mux_2589_nl <= MUX_s_1_2_2(or_3242_nl, mux_2587_nl, fsm_output(2));
  or_3231_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)) OR not_tmp_321;
  or_3229_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))))
      OR not_tmp_527;
  mux_2578_nl <= MUX_s_1_2_2(or_3231_nl, or_3229_nl, fsm_output(0));
  nand_242_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11101"))
      AND COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
      (fsm_output(3)) AND (NOT (fsm_output(7))));
  nand_243_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2577_nl <= MUX_s_1_2_2(nand_242_nl, nand_243_nl, fsm_output(0));
  mux_2579_nl <= MUX_s_1_2_2(mux_2578_nl, mux_2577_nl, fsm_output(4));
  nor_781_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_782_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111011"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2576_nl <= MUX_s_1_2_2(nor_781_nl, nor_782_nl, fsm_output(0));
  nand_133_nl <= NOT((fsm_output(4)) AND mux_2576_nl);
  mux_2580_nl <= MUX_s_1_2_2(mux_2579_nl, nand_133_nl, fsm_output(6));
  or_3232_nl <= (fsm_output(2)) OR mux_2580_nl;
  mux_2590_nl <= MUX_s_1_2_2(mux_2589_nl, or_3232_nl, fsm_output(5));
  vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2590_nl) AND (fsm_output(1));
  nor_773_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR not_tmp_560);
  and_555_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("00"))
      AND and_763_cse;
  mux_2602_nl <= MUX_s_1_2_2(nor_773_nl, and_555_nl, fsm_output(0));
  nor_774_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  nor_775_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7)));
  mux_2601_nl <= MUX_s_1_2_2(nor_774_nl, nor_775_nl, fsm_output(0));
  mux_2603_nl <= MUX_s_1_2_2(mux_2602_nl, mux_2601_nl, fsm_output(4));
  nor_776_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  nor_777_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (NOT (fsm_output(7))));
  mux_2599_nl <= MUX_s_1_2_2(nor_776_nl, nor_777_nl, fsm_output(0));
  nor_778_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_779_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2598_nl <= MUX_s_1_2_2(nor_778_nl, nor_779_nl, fsm_output(0));
  mux_2600_nl <= MUX_s_1_2_2(mux_2599_nl, mux_2598_nl, fsm_output(4));
  mux_2604_nl <= MUX_s_1_2_2(mux_2603_nl, mux_2600_nl, fsm_output(6));
  nand_409_nl <= NOT((fsm_output(2)) AND mux_2604_nl);
  or_3252_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR not_tmp_559;
  mux_2595_nl <= MUX_s_1_2_2(or_tmp_3138, or_3252_nl, fsm_output(0));
  or_3249_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2594_nl <= MUX_s_1_2_2(or_tmp_3134, or_3249_nl, fsm_output(0));
  mux_2596_nl <= MUX_s_1_2_2(mux_2595_nl, mux_2594_nl, fsm_output(4));
  or_3246_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2592_nl <= MUX_s_1_2_2(or_tmp_3132, or_3246_nl, fsm_output(0));
  or_3243_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2591_nl <= MUX_s_1_2_2(or_tmp_3128, or_3243_nl, fsm_output(0));
  mux_2593_nl <= MUX_s_1_2_2(mux_2592_nl, mux_2591_nl, fsm_output(4));
  mux_2597_nl <= MUX_s_1_2_2(mux_2596_nl, mux_2593_nl, fsm_output(6));
  or_4082_nl <= (fsm_output(2)) OR mux_2597_nl;
  mux_2605_nl <= MUX_s_1_2_2(nand_409_nl, or_4082_nl, fsm_output(5));
  vec_rsc_0_60_i_we_d_pff <= NOT(mux_2605_nl OR (fsm_output(1)));
  or_3285_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3284_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2618_nl <= MUX_s_1_2_2(or_3285_nl, or_3284_nl, fsm_output(0));
  or_3286_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2618_nl;
  or_3282_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR not_tmp_559;
  mux_2615_nl <= MUX_s_1_2_2(or_3282_nl, or_tmp_3138, fsm_output(0));
  or_3280_nl <= (NOT COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111100")) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2614_nl <= MUX_s_1_2_2(or_3280_nl, or_tmp_3134, fsm_output(0));
  mux_2616_nl <= MUX_s_1_2_2(mux_2615_nl, mux_2614_nl, fsm_output(4));
  or_3279_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111100")) OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  mux_2612_nl <= MUX_s_1_2_2(or_3279_nl, or_tmp_3132, fsm_output(0));
  or_3277_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111100")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2611_nl <= MUX_s_1_2_2(or_3277_nl, or_tmp_3128, fsm_output(0));
  mux_2613_nl <= MUX_s_1_2_2(mux_2612_nl, mux_2611_nl, fsm_output(4));
  mux_2617_nl <= MUX_s_1_2_2(mux_2616_nl, mux_2613_nl, fsm_output(6));
  mux_2619_nl <= MUX_s_1_2_2(or_3286_nl, mux_2617_nl, fsm_output(2));
  nand_237_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND and_763_cse);
  or_3273_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR not_tmp_544;
  mux_2608_nl <= MUX_s_1_2_2(nand_237_nl, or_3273_nl, fsm_output(0));
  or_3271_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (NOT COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm) OR (VEC_LOOP_j_10_0_sva_9_0(0))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_3270_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (NOT (fsm_output(3))) OR (fsm_output(7));
  mux_2607_nl <= MUX_s_1_2_2(or_3271_nl, or_3270_nl, fsm_output(0));
  mux_2609_nl <= MUX_s_1_2_2(mux_2608_nl, mux_2607_nl, fsm_output(4));
  nor_771_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_772_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2606_nl <= MUX_s_1_2_2(nor_771_nl, nor_772_nl, fsm_output(0));
  nand_135_nl <= NOT((fsm_output(4)) AND mux_2606_nl);
  mux_2610_nl <= MUX_s_1_2_2(mux_2609_nl, nand_135_nl, fsm_output(6));
  or_3276_nl <= (fsm_output(2)) OR mux_2610_nl;
  mux_2620_nl <= MUX_s_1_2_2(mux_2619_nl, or_3276_nl, fsm_output(5));
  vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2620_nl) AND (fsm_output(1));
  nor_764_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR not_tmp_560);
  nor_765_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (VEC_LOOP_j_10_0_sva_9_0(1))))) OR not_tmp_321);
  mux_2632_nl <= MUX_s_1_2_2(nor_764_nl, nor_765_nl, fsm_output(0));
  and_552_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_553_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  mux_2631_nl <= MUX_s_1_2_2(and_552_nl, and_553_nl, fsm_output(0));
  mux_2633_nl <= MUX_s_1_2_2(mux_2632_nl, mux_2631_nl, fsm_output(4));
  and_815_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7));
  and_822_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT (fsm_output(3))) AND (fsm_output(7));
  mux_2629_nl <= MUX_s_1_2_2(and_815_nl, and_822_nl, fsm_output(0));
  nor_768_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_769_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2628_nl <= MUX_s_1_2_2(nor_768_nl, nor_769_nl, fsm_output(0));
  mux_2630_nl <= MUX_s_1_2_2(mux_2629_nl, mux_2628_nl, fsm_output(4));
  mux_2634_nl <= MUX_s_1_2_2(mux_2633_nl, mux_2630_nl, fsm_output(6));
  nand_408_nl <= NOT((fsm_output(2)) AND mux_2634_nl);
  or_3296_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_565;
  mux_2625_nl <= MUX_s_1_2_2(or_tmp_3182, or_3296_nl, fsm_output(0));
  nand_232_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2624_nl <= MUX_s_1_2_2(or_tmp_3178, nand_232_nl, fsm_output(0));
  mux_2626_nl <= MUX_s_1_2_2(mux_2625_nl, mux_2624_nl, fsm_output(4));
  nand_474_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2622_nl <= MUX_s_1_2_2(or_tmp_3176, nand_474_nl, fsm_output(0));
  or_3287_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2621_nl <= MUX_s_1_2_2(or_tmp_3172, or_3287_nl, fsm_output(0));
  mux_2623_nl <= MUX_s_1_2_2(mux_2622_nl, mux_2621_nl, fsm_output(4));
  mux_2627_nl <= MUX_s_1_2_2(mux_2626_nl, mux_2623_nl, fsm_output(6));
  or_4081_nl <= (fsm_output(2)) OR mux_2627_nl;
  mux_2635_nl <= MUX_s_1_2_2(nand_408_nl, or_4081_nl, fsm_output(5));
  vec_rsc_0_61_i_we_d_pff <= NOT(mux_2635_nl OR (fsm_output(1)));
  or_3328_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3327_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2648_nl <= MUX_s_1_2_2(or_3328_nl, or_3327_nl, fsm_output(0));
  or_3329_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2648_nl;
  or_3325_nl <= (NOT COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 1)/=STD_LOGIC_VECTOR'("10")) OR not_tmp_565;
  mux_2645_nl <= MUX_s_1_2_2(or_3325_nl, or_tmp_3182, fsm_output(0));
  nand_223_nl <= NOT(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111101")) AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2644_nl <= MUX_s_1_2_2(nand_223_nl, or_tmp_3178, fsm_output(0));
  mux_2646_nl <= MUX_s_1_2_2(mux_2645_nl, mux_2644_nl, fsm_output(4));
  nand_396_nl <= NOT(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111101")) AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2642_nl <= MUX_s_1_2_2(nand_396_nl, or_tmp_3176, fsm_output(0));
  or_3320_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111101")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2641_nl <= MUX_s_1_2_2(or_3320_nl, or_tmp_3172, fsm_output(0));
  mux_2643_nl <= MUX_s_1_2_2(mux_2642_nl, mux_2641_nl, fsm_output(4));
  mux_2647_nl <= MUX_s_1_2_2(mux_2646_nl, mux_2643_nl, fsm_output(6));
  mux_2649_nl <= MUX_s_1_2_2(or_3329_nl, mux_2647_nl, fsm_output(2));
  or_3318_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)) OR not_tmp_321;
  or_3316_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) OR (NOT((COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      AND (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      AND (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(4))
      AND (fsm_output(3)) AND (fsm_output(7))));
  mux_2638_nl <= MUX_s_1_2_2(or_3318_nl, or_3316_nl, fsm_output(0));
  nand_227_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
      (fsm_output(3)) AND (NOT (fsm_output(7))));
  nand_228_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2637_nl <= MUX_s_1_2_2(nand_227_nl, nand_228_nl, fsm_output(0));
  mux_2639_nl <= MUX_s_1_2_2(mux_2638_nl, mux_2637_nl, fsm_output(4));
  nor_762_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_763_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111101"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2636_nl <= MUX_s_1_2_2(nor_762_nl, nor_763_nl, fsm_output(0));
  nand_137_nl <= NOT((fsm_output(4)) AND mux_2636_nl);
  mux_2640_nl <= MUX_s_1_2_2(mux_2639_nl, nand_137_nl, fsm_output(6));
  or_3319_nl <= (fsm_output(2)) OR mux_2640_nl;
  mux_2650_nl <= MUX_s_1_2_2(mux_2649_nl, or_3319_nl, fsm_output(5));
  vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2650_nl) AND (fsm_output(1));
  nor_756_nl <= NOT((COMP_LOOP_acc_10_cse_10_1_5_sva(0)) OR (NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5
      DOWNTO 1)=STD_LOGIC_VECTOR'("11111")) AND (fsm_output(3)) AND (fsm_output(7)))));
  and_548_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"))
      AND and_763_cse;
  mux_2662_nl <= MUX_s_1_2_2(nor_756_nl, and_548_nl, fsm_output(0));
  and_549_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_550_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  mux_2661_nl <= MUX_s_1_2_2(and_549_nl, and_550_nl, fsm_output(0));
  mux_2663_nl <= MUX_s_1_2_2(mux_2662_nl, mux_2661_nl, fsm_output(4));
  and_816_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7));
  and_823_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0))) AND (NOT (fsm_output(3))) AND (fsm_output(7));
  mux_2659_nl <= MUX_s_1_2_2(and_816_nl, and_823_nl, fsm_output(0));
  nor_759_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_760_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11111"))
      OR (VEC_LOOP_j_10_0_sva_9_0(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2658_nl <= MUX_s_1_2_2(nor_759_nl, nor_760_nl, fsm_output(0));
  mux_2660_nl <= MUX_s_1_2_2(mux_2659_nl, mux_2658_nl, fsm_output(4));
  mux_2664_nl <= MUX_s_1_2_2(mux_2663_nl, mux_2660_nl, fsm_output(6));
  nand_407_nl <= NOT((fsm_output(2)) AND mux_2664_nl);
  or_3339_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR not_tmp_559;
  mux_2655_nl <= MUX_s_1_2_2(or_tmp_3225, or_3339_nl, fsm_output(0));
  nand_218_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2654_nl <= MUX_s_1_2_2(or_tmp_3221, nand_218_nl, fsm_output(0));
  mux_2656_nl <= MUX_s_1_2_2(mux_2655_nl, mux_2654_nl, fsm_output(4));
  nand_473_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2652_nl <= MUX_s_1_2_2(or_tmp_3219, nand_473_nl, fsm_output(0));
  or_3330_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2651_nl <= MUX_s_1_2_2(or_tmp_3215, or_3330_nl, fsm_output(0));
  mux_2653_nl <= MUX_s_1_2_2(mux_2652_nl, mux_2651_nl, fsm_output(4));
  mux_2657_nl <= MUX_s_1_2_2(mux_2656_nl, mux_2653_nl, fsm_output(6));
  or_4080_nl <= (fsm_output(2)) OR mux_2657_nl;
  mux_2665_nl <= MUX_s_1_2_2(nand_407_nl, or_4080_nl, fsm_output(5));
  vec_rsc_0_62_i_we_d_pff <= NOT(mux_2665_nl OR (fsm_output(1)));
  or_3371_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  or_3370_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(7));
  mux_2678_nl <= MUX_s_1_2_2(or_3371_nl, or_3370_nl, fsm_output(0));
  or_3372_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2678_nl;
  or_3368_nl <= (NOT(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("110")))) OR not_tmp_559;
  mux_2675_nl <= MUX_s_1_2_2(or_3368_nl, or_tmp_3225, fsm_output(0));
  nand_210_nl <= NOT(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111110")) AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2674_nl <= MUX_s_1_2_2(nand_210_nl, or_tmp_3221, fsm_output(0));
  mux_2676_nl <= MUX_s_1_2_2(mux_2675_nl, mux_2674_nl, fsm_output(4));
  nand_394_nl <= NOT(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111110")) AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2672_nl <= MUX_s_1_2_2(nand_394_nl, or_tmp_3219, fsm_output(0));
  or_3363_nl <= (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111110")) OR (fsm_output(3)) OR (fsm_output(7));
  mux_2671_nl <= MUX_s_1_2_2(or_3363_nl, or_tmp_3215, fsm_output(0));
  mux_2673_nl <= MUX_s_1_2_2(mux_2672_nl, mux_2671_nl, fsm_output(4));
  mux_2677_nl <= MUX_s_1_2_2(mux_2676_nl, mux_2673_nl, fsm_output(6));
  mux_2679_nl <= MUX_s_1_2_2(or_3372_nl, mux_2677_nl, fsm_output(2));
  nand_212_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND and_763_cse);
  or_3359_nl <= (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(1))) OR (NOT (COMP_LOOP_acc_10_cse_10_1_7_sva(3)))
      OR (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) OR not_tmp_544;
  mux_2668_nl <= MUX_s_1_2_2(nand_212_nl, or_3359_nl, fsm_output(0));
  nand_213_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm AND (NOT (VEC_LOOP_j_10_0_sva_9_0(0)))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  nand_214_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2667_nl <= MUX_s_1_2_2(nand_213_nl, nand_214_nl, fsm_output(0));
  mux_2669_nl <= MUX_s_1_2_2(mux_2668_nl, mux_2667_nl, fsm_output(4));
  nor_754_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (fsm_output(3)) OR (fsm_output(7)));
  nor_755_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111110"))
      OR (fsm_output(3)) OR (fsm_output(7)));
  mux_2666_nl <= MUX_s_1_2_2(nor_754_nl, nor_755_nl, fsm_output(0));
  nand_139_nl <= NOT((fsm_output(4)) AND mux_2666_nl);
  mux_2670_nl <= MUX_s_1_2_2(mux_2669_nl, nand_139_nl, fsm_output(6));
  or_3362_nl <= (fsm_output(2)) OR mux_2670_nl;
  mux_2680_nl <= MUX_s_1_2_2(mux_2679_nl, or_3362_nl, fsm_output(5));
  vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2680_nl) AND (fsm_output(1));
  and_539_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)) AND (fsm_output(7));
  and_540_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)) AND (fsm_output(7));
  mux_2692_nl <= MUX_s_1_2_2(and_539_nl, and_540_nl, fsm_output(0));
  and_541_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_542_nl <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7)));
  mux_2691_nl <= MUX_s_1_2_2(and_541_nl, and_542_nl, fsm_output(0));
  mux_2693_nl <= MUX_s_1_2_2(mux_2692_nl, mux_2691_nl, fsm_output(4));
  and_817_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7));
  and_824_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT (fsm_output(3))) AND (fsm_output(7));
  mux_2689_nl <= MUX_s_1_2_2(and_817_nl, and_824_nl, fsm_output(0));
  and_543_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7)));
  and_544_nl <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7)));
  mux_2688_nl <= MUX_s_1_2_2(and_543_nl, and_544_nl, fsm_output(0));
  mux_2690_nl <= MUX_s_1_2_2(mux_2689_nl, mux_2688_nl, fsm_output(4));
  mux_2694_nl <= MUX_s_1_2_2(mux_2693_nl, mux_2690_nl, fsm_output(6));
  nand_406_nl <= NOT((fsm_output(2)) AND mux_2694_nl);
  mux_2685_nl <= MUX_s_1_2_2(nor_tmp_307, nor_tmp_306, fsm_output(0));
  nand_203_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2684_nl <= MUX_s_1_2_2(or_tmp_3264, nand_203_nl, fsm_output(0));
  mux_2686_nl <= MUX_s_1_2_2((NOT mux_2685_nl), mux_2684_nl, fsm_output(4));
  nand_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2682_nl <= MUX_s_1_2_2(or_tmp_3262, nand_nl, fsm_output(0));
  nand_205_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7))));
  mux_2681_nl <= MUX_s_1_2_2(or_tmp_3258, nand_205_nl, fsm_output(0));
  mux_2683_nl <= MUX_s_1_2_2(mux_2682_nl, mux_2681_nl, fsm_output(4));
  mux_2687_nl <= MUX_s_1_2_2(mux_2686_nl, mux_2683_nl, fsm_output(6));
  or_4079_nl <= (fsm_output(2)) OR mux_2687_nl;
  mux_2695_nl <= MUX_s_1_2_2(nand_406_nl, or_4079_nl, fsm_output(5));
  vec_rsc_0_63_i_we_d_pff <= NOT(mux_2695_nl OR (fsm_output(1)));
  nand_192_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7))));
  nand_193_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7))));
  mux_2708_nl <= MUX_s_1_2_2(nand_192_nl, nand_193_nl, fsm_output(0));
  or_3405_nl <= (fsm_output(6)) OR (fsm_output(4)) OR mux_2708_nl;
  and_535_nl <= COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm AND nor_tmp_306;
  mux_2705_nl <= MUX_s_1_2_2(and_535_nl, nor_tmp_307, fsm_output(0));
  nand_194_nl <= NOT(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111111")) AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2704_nl <= MUX_s_1_2_2(nand_194_nl, or_tmp_3264, fsm_output(0));
  mux_2706_nl <= MUX_s_1_2_2((NOT mux_2705_nl), mux_2704_nl, fsm_output(4));
  nand_392_nl <= NOT(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111111")) AND (NOT (fsm_output(3))) AND (fsm_output(7)));
  mux_2702_nl <= MUX_s_1_2_2(nand_392_nl, or_tmp_3262, fsm_output(0));
  nand_196_nl <= NOT(COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm AND CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(5
      DOWNTO 0)=STD_LOGIC_VECTOR'("111111")) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7))));
  mux_2701_nl <= MUX_s_1_2_2(nand_196_nl, or_tmp_3258, fsm_output(0));
  mux_2703_nl <= MUX_s_1_2_2(mux_2702_nl, mux_2701_nl, fsm_output(4));
  mux_2707_nl <= MUX_s_1_2_2(mux_2706_nl, mux_2703_nl, fsm_output(6));
  mux_2709_nl <= MUX_s_1_2_2(or_3405_nl, mux_2707_nl, fsm_output(2));
  or_4002_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)) OR not_tmp_321;
  nand_198_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)) AND (fsm_output(7)));
  mux_2698_nl <= MUX_s_1_2_2(or_4002_nl, nand_198_nl, fsm_output(0));
  nand_199_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111"))
      AND COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
      (fsm_output(3)) AND (NOT (fsm_output(7))));
  nand_200_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_3_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)) AND (NOT (fsm_output(7))));
  mux_2697_nl <= MUX_s_1_2_2(nand_199_nl, nand_200_nl, fsm_output(0));
  mux_2699_nl <= MUX_s_1_2_2(mux_2698_nl, mux_2697_nl, fsm_output(4));
  and_536_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7)));
  and_537_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3))) AND (NOT (fsm_output(7)));
  mux_2696_nl <= MUX_s_1_2_2(and_536_nl, and_537_nl, fsm_output(0));
  nand_141_nl <= NOT((fsm_output(4)) AND mux_2696_nl);
  mux_2700_nl <= MUX_s_1_2_2(mux_2699_nl, nand_141_nl, fsm_output(6));
  or_3396_nl <= (fsm_output(2)) OR mux_2700_nl;
  mux_2710_nl <= MUX_s_1_2_2(mux_2709_nl, or_3396_nl, fsm_output(5));
  vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d <= (NOT mux_2710_nl) AND (fsm_output(1));
  twiddle_rsc_0_0_i_radr_d_pff <= MUX1HOT_v_4_7_2((z_out_8(6 DOWNTO 3)), (z_out_7(9
      DOWNTO 6)), (z_out_7(8 DOWNTO 5)), (COMP_LOOP_5_tmp_mul_idiv_sva(7 DOWNTO 4)),
      (COMP_LOOP_2_tmp_mul_idiv_sva(9 DOWNTO 6)), (COMP_LOOP_3_tmp_lshift_ncse_sva(8
      DOWNTO 5)), (COMP_LOOP_2_tmp_lshift_ncse_sva(9 DOWNTO 6)), STD_LOGIC_VECTOR'(
      and_dcpl_74 & COMP_LOOP_or_110_rgt & and_dcpl_258 & and_dcpl_260 & and_dcpl_261
      & and_dcpl_263 & and_dcpl_265));
  nor_746_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)));
  nor_743_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(3))));
  nor_744_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (NOT (fsm_output(3))));
  mux_2715_nl <= MUX_s_1_2_2(nor_743_nl, nor_744_nl, fsm_output(0));
  nor_745_nl <= NOT(CONV_SL_1_1(z_out_8(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR
      (fsm_output(3)));
  mux_2714_nl <= MUX_s_1_2_2(nor_745_nl, nor_746_cse, fsm_output(0));
  mux_2716_nl <= MUX_s_1_2_2(mux_2715_nl, mux_2714_nl, fsm_output(1));
  nor_747_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR (fsm_output(3)));
  mux_2712_nl <= MUX_s_1_2_2(nor_747_nl, nor_746_cse, fsm_output(0));
  nor_749_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(3)));
  nor_750_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000000"))
      OR (fsm_output(3)));
  mux_2711_nl <= MUX_s_1_2_2(nor_749_nl, nor_750_nl, fsm_output(0));
  mux_2713_nl <= MUX_s_1_2_2(mux_2712_nl, mux_2711_nl, fsm_output(1));
  mux_2717_nl <= MUX_s_1_2_2(mux_2716_nl, mux_2713_nl, fsm_output(2));
  twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2717_nl AND and_dcpl_268;
  twiddle_rsc_0_1_i_radr_d_pff <= z_out_7(9 DOWNTO 6);
  nor_740_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_739_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("00000"))
      OR nand_191_cse);
  mux_2719_nl <= MUX_s_1_2_2(nor_739_nl, nor_740_cse, fsm_output(0));
  nor_742_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000001"))
      OR (fsm_output(3)));
  mux_2718_nl <= MUX_s_1_2_2(nor_740_cse, nor_742_nl, fsm_output(0));
  mux_2720_nl <= MUX_s_1_2_2(mux_2719_nl, mux_2718_nl, fsm_output(1));
  twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2720_nl AND and_dcpl_268;
  twiddle_rsc_0_2_i_radr_d_pff <= MUX_v_4_2_2((z_out_7(9 DOWNTO 6)), (z_out_7(8 DOWNTO
      5)), COMP_LOOP_tmp_or_43_cse);
  nor_735_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(3)));
  nor_734_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00001"))
      OR (fsm_output(3)));
  nor_733_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2723_nl <= MUX_s_1_2_2(nor_734_cse, nor_735_cse, fsm_output(0));
  mux_2724_nl <= MUX_s_1_2_2(nor_733_nl, mux_2723_nl, fsm_output(2));
  nor_736_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2721_nl <= MUX_s_1_2_2(nor_735_cse, nor_734_cse, fsm_output(0));
  mux_2722_nl <= MUX_s_1_2_2(nor_736_nl, mux_2721_nl, fsm_output(2));
  mux_2725_nl <= MUX_s_1_2_2(mux_2724_nl, mux_2722_nl, fsm_output(1));
  twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2725_nl AND and_dcpl_268;
  nor_730_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_729_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_190_cse);
  mux_2727_nl <= MUX_s_1_2_2(nor_729_nl, nor_730_cse, fsm_output(0));
  nor_732_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000011"))
      OR (fsm_output(3)));
  mux_2726_nl <= MUX_s_1_2_2(nor_730_cse, nor_732_nl, fsm_output(0));
  mux_2728_nl <= MUX_s_1_2_2(mux_2727_nl, mux_2726_nl, fsm_output(1));
  twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2728_nl AND and_dcpl_268;
  twiddle_rsc_0_4_i_radr_d_pff <= MUX1HOT_v_4_6_2((z_out_7(9 DOWNTO 6)), (z_out_7(8
      DOWNTO 5)), (COMP_LOOP_5_tmp_mul_idiv_sva(7 DOWNTO 4)), (COMP_LOOP_2_tmp_mul_idiv_sva(9
      DOWNTO 6)), (COMP_LOOP_3_tmp_lshift_ncse_sva(8 DOWNTO 5)), (COMP_LOOP_2_tmp_lshift_ncse_sva(9
      DOWNTO 6)), STD_LOGIC_VECTOR'( COMP_LOOP_or_110_rgt & and_dcpl_258 & and_dcpl_260
      & and_dcpl_261 & and_dcpl_263 & and_dcpl_265));
  nor_722_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(3))));
  nor_723_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT (fsm_output(3))));
  mux_2732_nl <= MUX_s_1_2_2(nor_722_nl, nor_723_nl, fsm_output(0));
  nor_724_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(3)));
  nor_725_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)));
  mux_2731_nl <= MUX_s_1_2_2(nor_724_nl, nor_725_nl, fsm_output(0));
  mux_2733_nl <= MUX_s_1_2_2(mux_2732_nl, mux_2731_nl, fsm_output(2));
  nor_726_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  nor_727_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(3)));
  nor_728_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000100"))
      OR (fsm_output(3)));
  mux_2729_nl <= MUX_s_1_2_2(nor_727_nl, nor_728_nl, fsm_output(0));
  mux_2730_nl <= MUX_s_1_2_2(nor_726_nl, mux_2729_nl, fsm_output(2));
  mux_2734_nl <= MUX_s_1_2_2(mux_2733_nl, mux_2730_nl, fsm_output(1));
  twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2734_nl AND and_dcpl_268;
  nor_719_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_718_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("00010"))
      OR nand_191_cse);
  mux_2736_nl <= MUX_s_1_2_2(nor_718_nl, nor_719_cse, fsm_output(0));
  nor_721_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000101"))
      OR (fsm_output(3)));
  mux_2735_nl <= MUX_s_1_2_2(nor_719_cse, nor_721_nl, fsm_output(0));
  mux_2737_nl <= MUX_s_1_2_2(mux_2736_nl, mux_2735_nl, fsm_output(1));
  twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2737_nl AND and_dcpl_268;
  nor_714_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(3)));
  nor_713_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00011"))
      OR (fsm_output(3)));
  nor_712_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2740_nl <= MUX_s_1_2_2(nor_713_cse, nor_714_cse, fsm_output(0));
  mux_2741_nl <= MUX_s_1_2_2(nor_712_nl, mux_2740_nl, fsm_output(2));
  nor_715_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2738_nl <= MUX_s_1_2_2(nor_714_cse, nor_713_cse, fsm_output(0));
  mux_2739_nl <= MUX_s_1_2_2(nor_715_nl, mux_2738_nl, fsm_output(2));
  mux_2742_nl <= MUX_s_1_2_2(mux_2741_nl, mux_2739_nl, fsm_output(1));
  twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2742_nl AND and_dcpl_268;
  nor_709_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_708_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000"))
      OR nand_188_cse);
  mux_2744_nl <= MUX_s_1_2_2(nor_708_nl, nor_709_cse, fsm_output(0));
  nor_711_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("000111"))
      OR (fsm_output(3)));
  mux_2743_nl <= MUX_s_1_2_2(nor_709_cse, nor_711_nl, fsm_output(0));
  mux_2745_nl <= MUX_s_1_2_2(mux_2744_nl, mux_2743_nl, fsm_output(1));
  twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2745_nl AND and_dcpl_268;
  nor_703_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)));
  nor_700_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(3))));
  nor_701_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (NOT (fsm_output(3))));
  mux_2750_nl <= MUX_s_1_2_2(nor_700_nl, nor_701_nl, fsm_output(0));
  nor_702_nl <= NOT(CONV_SL_1_1(z_out_8(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR
      (fsm_output(3)));
  mux_2749_nl <= MUX_s_1_2_2(nor_702_nl, nor_703_cse, fsm_output(0));
  mux_2751_nl <= MUX_s_1_2_2(mux_2750_nl, mux_2749_nl, fsm_output(1));
  nor_704_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00100"))
      OR (fsm_output(3)));
  mux_2747_nl <= MUX_s_1_2_2(nor_704_nl, nor_703_cse, fsm_output(0));
  nor_706_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(3)));
  nor_707_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001000"))
      OR (fsm_output(3)));
  mux_2746_nl <= MUX_s_1_2_2(nor_706_nl, nor_707_nl, fsm_output(0));
  mux_2748_nl <= MUX_s_1_2_2(mux_2747_nl, mux_2746_nl, fsm_output(1));
  mux_2752_nl <= MUX_s_1_2_2(mux_2751_nl, mux_2748_nl, fsm_output(2));
  twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2752_nl AND and_dcpl_268;
  nor_697_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_696_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("00100"))
      OR nand_191_cse);
  mux_2754_nl <= MUX_s_1_2_2(nor_696_nl, nor_697_cse, fsm_output(0));
  nor_699_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001001"))
      OR (fsm_output(3)));
  mux_2753_nl <= MUX_s_1_2_2(nor_697_cse, nor_699_nl, fsm_output(0));
  mux_2755_nl <= MUX_s_1_2_2(mux_2754_nl, mux_2753_nl, fsm_output(1));
  twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2755_nl AND and_dcpl_268;
  nor_692_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(3)));
  nor_691_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00101"))
      OR (fsm_output(3)));
  nor_690_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2758_nl <= MUX_s_1_2_2(nor_691_cse, nor_692_cse, fsm_output(0));
  mux_2759_nl <= MUX_s_1_2_2(nor_690_nl, mux_2758_nl, fsm_output(2));
  nor_693_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2756_nl <= MUX_s_1_2_2(nor_692_cse, nor_691_cse, fsm_output(0));
  mux_2757_nl <= MUX_s_1_2_2(nor_693_nl, mux_2756_nl, fsm_output(2));
  mux_2760_nl <= MUX_s_1_2_2(mux_2759_nl, mux_2757_nl, fsm_output(1));
  twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2760_nl AND and_dcpl_268;
  nor_687_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_686_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("0010"))
      OR nand_190_cse);
  mux_2762_nl <= MUX_s_1_2_2(nor_686_nl, nor_687_cse, fsm_output(0));
  nor_689_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001011"))
      OR (fsm_output(3)));
  mux_2761_nl <= MUX_s_1_2_2(nor_687_cse, nor_689_nl, fsm_output(0));
  mux_2763_nl <= MUX_s_1_2_2(mux_2762_nl, mux_2761_nl, fsm_output(1));
  twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2763_nl AND and_dcpl_268;
  nor_679_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(3))));
  nor_680_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT (fsm_output(3))));
  mux_2767_nl <= MUX_s_1_2_2(nor_679_nl, nor_680_nl, fsm_output(0));
  nor_681_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(3)));
  nor_682_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)));
  mux_2766_nl <= MUX_s_1_2_2(nor_681_nl, nor_682_nl, fsm_output(0));
  mux_2768_nl <= MUX_s_1_2_2(mux_2767_nl, mux_2766_nl, fsm_output(2));
  nor_683_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  nor_684_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(3)));
  nor_685_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001100"))
      OR (fsm_output(3)));
  mux_2764_nl <= MUX_s_1_2_2(nor_684_nl, nor_685_nl, fsm_output(0));
  mux_2765_nl <= MUX_s_1_2_2(nor_683_nl, mux_2764_nl, fsm_output(2));
  mux_2769_nl <= MUX_s_1_2_2(mux_2768_nl, mux_2765_nl, fsm_output(1));
  twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2769_nl AND and_dcpl_268;
  nor_676_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_675_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("00110"))
      OR nand_191_cse);
  mux_2771_nl <= MUX_s_1_2_2(nor_675_nl, nor_676_cse, fsm_output(0));
  nor_678_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001101"))
      OR (fsm_output(3)));
  mux_2770_nl <= MUX_s_1_2_2(nor_676_cse, nor_678_nl, fsm_output(0));
  mux_2772_nl <= MUX_s_1_2_2(mux_2771_nl, mux_2770_nl, fsm_output(1));
  twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2772_nl AND and_dcpl_268;
  nor_671_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(3)));
  nor_670_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00111"))
      OR (fsm_output(3)));
  nor_669_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2775_nl <= MUX_s_1_2_2(nor_670_cse, nor_671_cse, fsm_output(0));
  mux_2776_nl <= MUX_s_1_2_2(nor_669_nl, mux_2775_nl, fsm_output(2));
  nor_672_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2773_nl <= MUX_s_1_2_2(nor_671_cse, nor_670_cse, fsm_output(0));
  mux_2774_nl <= MUX_s_1_2_2(nor_672_nl, mux_2773_nl, fsm_output(2));
  mux_2777_nl <= MUX_s_1_2_2(mux_2776_nl, mux_2774_nl, fsm_output(1));
  twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2777_nl AND and_dcpl_268;
  nor_666_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_665_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00"))
      OR nand_184_cse);
  mux_2779_nl <= MUX_s_1_2_2(nor_665_nl, nor_666_cse, fsm_output(0));
  nor_668_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("001111"))
      OR (fsm_output(3)));
  mux_2778_nl <= MUX_s_1_2_2(nor_666_cse, nor_668_nl, fsm_output(0));
  mux_2780_nl <= MUX_s_1_2_2(mux_2779_nl, mux_2778_nl, fsm_output(1));
  twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2780_nl AND and_dcpl_268;
  nor_660_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)));
  nor_657_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(3))));
  nor_658_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (NOT (fsm_output(3))));
  mux_2785_nl <= MUX_s_1_2_2(nor_657_nl, nor_658_nl, fsm_output(0));
  nor_659_nl <= NOT(CONV_SL_1_1(z_out_8(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR
      (fsm_output(3)));
  mux_2784_nl <= MUX_s_1_2_2(nor_659_nl, nor_660_cse, fsm_output(0));
  mux_2786_nl <= MUX_s_1_2_2(mux_2785_nl, mux_2784_nl, fsm_output(1));
  nor_661_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR (fsm_output(3)));
  mux_2782_nl <= MUX_s_1_2_2(nor_661_nl, nor_660_cse, fsm_output(0));
  nor_663_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(3)));
  nor_664_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010000"))
      OR (fsm_output(3)));
  mux_2781_nl <= MUX_s_1_2_2(nor_663_nl, nor_664_nl, fsm_output(0));
  mux_2783_nl <= MUX_s_1_2_2(mux_2782_nl, mux_2781_nl, fsm_output(1));
  mux_2787_nl <= MUX_s_1_2_2(mux_2786_nl, mux_2783_nl, fsm_output(2));
  twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2787_nl AND and_dcpl_268;
  nor_654_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_653_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("01000"))
      OR nand_191_cse);
  mux_2789_nl <= MUX_s_1_2_2(nor_653_nl, nor_654_cse, fsm_output(0));
  nor_656_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010001"))
      OR (fsm_output(3)));
  mux_2788_nl <= MUX_s_1_2_2(nor_654_cse, nor_656_nl, fsm_output(0));
  mux_2790_nl <= MUX_s_1_2_2(mux_2789_nl, mux_2788_nl, fsm_output(1));
  twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2790_nl AND and_dcpl_268;
  nor_649_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(3)));
  nor_648_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01001"))
      OR (fsm_output(3)));
  nor_647_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2793_nl <= MUX_s_1_2_2(nor_648_cse, nor_649_cse, fsm_output(0));
  mux_2794_nl <= MUX_s_1_2_2(nor_647_nl, mux_2793_nl, fsm_output(2));
  nor_650_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2791_nl <= MUX_s_1_2_2(nor_649_cse, nor_648_cse, fsm_output(0));
  mux_2792_nl <= MUX_s_1_2_2(nor_650_nl, mux_2791_nl, fsm_output(2));
  mux_2795_nl <= MUX_s_1_2_2(mux_2794_nl, mux_2792_nl, fsm_output(1));
  twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2795_nl AND and_dcpl_268;
  nor_644_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_643_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_190_cse);
  mux_2797_nl <= MUX_s_1_2_2(nor_643_nl, nor_644_cse, fsm_output(0));
  nor_646_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010011"))
      OR (fsm_output(3)));
  mux_2796_nl <= MUX_s_1_2_2(nor_644_cse, nor_646_nl, fsm_output(0));
  mux_2798_nl <= MUX_s_1_2_2(mux_2797_nl, mux_2796_nl, fsm_output(1));
  twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2798_nl AND and_dcpl_268;
  nor_636_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(3))));
  nor_637_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (NOT (fsm_output(3))));
  mux_2802_nl <= MUX_s_1_2_2(nor_636_nl, nor_637_nl, fsm_output(0));
  nor_638_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(3)));
  nor_639_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)));
  mux_2801_nl <= MUX_s_1_2_2(nor_638_nl, nor_639_nl, fsm_output(0));
  mux_2803_nl <= MUX_s_1_2_2(mux_2802_nl, mux_2801_nl, fsm_output(2));
  nor_640_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  nor_641_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(3)));
  nor_642_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010100"))
      OR (fsm_output(3)));
  mux_2799_nl <= MUX_s_1_2_2(nor_641_nl, nor_642_nl, fsm_output(0));
  mux_2800_nl <= MUX_s_1_2_2(nor_640_nl, mux_2799_nl, fsm_output(2));
  mux_2804_nl <= MUX_s_1_2_2(mux_2803_nl, mux_2800_nl, fsm_output(1));
  twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2804_nl AND and_dcpl_268;
  nor_633_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_632_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("01010"))
      OR nand_191_cse);
  mux_2806_nl <= MUX_s_1_2_2(nor_632_nl, nor_633_cse, fsm_output(0));
  nor_635_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010101"))
      OR (fsm_output(3)));
  mux_2805_nl <= MUX_s_1_2_2(nor_633_cse, nor_635_nl, fsm_output(0));
  mux_2807_nl <= MUX_s_1_2_2(mux_2806_nl, mux_2805_nl, fsm_output(1));
  twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2807_nl AND and_dcpl_268;
  nor_628_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(3)));
  nor_627_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01011"))
      OR (fsm_output(3)));
  nor_626_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2810_nl <= MUX_s_1_2_2(nor_627_cse, nor_628_cse, fsm_output(0));
  mux_2811_nl <= MUX_s_1_2_2(nor_626_nl, mux_2810_nl, fsm_output(2));
  nor_629_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2808_nl <= MUX_s_1_2_2(nor_628_cse, nor_627_cse, fsm_output(0));
  mux_2809_nl <= MUX_s_1_2_2(nor_629_nl, mux_2808_nl, fsm_output(2));
  mux_2812_nl <= MUX_s_1_2_2(mux_2811_nl, mux_2809_nl, fsm_output(1));
  twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2812_nl AND and_dcpl_268;
  nor_623_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_622_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("010"))
      OR nand_188_cse);
  mux_2814_nl <= MUX_s_1_2_2(nor_622_nl, nor_623_cse, fsm_output(0));
  nor_625_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("010111"))
      OR (fsm_output(3)));
  mux_2813_nl <= MUX_s_1_2_2(nor_623_cse, nor_625_nl, fsm_output(0));
  mux_2815_nl <= MUX_s_1_2_2(mux_2814_nl, mux_2813_nl, fsm_output(1));
  twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2815_nl AND and_dcpl_268;
  nor_617_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)));
  nor_614_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(3))));
  nor_615_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (NOT (fsm_output(3))));
  mux_2820_nl <= MUX_s_1_2_2(nor_614_nl, nor_615_nl, fsm_output(0));
  nor_616_nl <= NOT(CONV_SL_1_1(z_out_8(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR
      (fsm_output(3)));
  mux_2819_nl <= MUX_s_1_2_2(nor_616_nl, nor_617_cse, fsm_output(0));
  mux_2821_nl <= MUX_s_1_2_2(mux_2820_nl, mux_2819_nl, fsm_output(1));
  nor_618_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01100"))
      OR (fsm_output(3)));
  mux_2817_nl <= MUX_s_1_2_2(nor_618_nl, nor_617_cse, fsm_output(0));
  nor_620_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(3)));
  nor_621_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011000"))
      OR (fsm_output(3)));
  mux_2816_nl <= MUX_s_1_2_2(nor_620_nl, nor_621_nl, fsm_output(0));
  mux_2818_nl <= MUX_s_1_2_2(mux_2817_nl, mux_2816_nl, fsm_output(1));
  mux_2822_nl <= MUX_s_1_2_2(mux_2821_nl, mux_2818_nl, fsm_output(2));
  twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2822_nl AND and_dcpl_268;
  nor_611_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_610_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("01100"))
      OR nand_191_cse);
  mux_2824_nl <= MUX_s_1_2_2(nor_610_nl, nor_611_cse, fsm_output(0));
  nor_613_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011001"))
      OR (fsm_output(3)));
  mux_2823_nl <= MUX_s_1_2_2(nor_611_cse, nor_613_nl, fsm_output(0));
  mux_2825_nl <= MUX_s_1_2_2(mux_2824_nl, mux_2823_nl, fsm_output(1));
  twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2825_nl AND and_dcpl_268;
  nor_606_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(3)));
  nor_605_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01101"))
      OR (fsm_output(3)));
  nor_604_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2828_nl <= MUX_s_1_2_2(nor_605_cse, nor_606_cse, fsm_output(0));
  mux_2829_nl <= MUX_s_1_2_2(nor_604_nl, mux_2828_nl, fsm_output(2));
  nor_607_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2826_nl <= MUX_s_1_2_2(nor_606_cse, nor_605_cse, fsm_output(0));
  mux_2827_nl <= MUX_s_1_2_2(nor_607_nl, mux_2826_nl, fsm_output(2));
  mux_2830_nl <= MUX_s_1_2_2(mux_2829_nl, mux_2827_nl, fsm_output(1));
  twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2830_nl AND and_dcpl_268;
  nor_601_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_600_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("0110"))
      OR nand_190_cse);
  mux_2832_nl <= MUX_s_1_2_2(nor_600_nl, nor_601_cse, fsm_output(0));
  nor_603_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011011"))
      OR (fsm_output(3)));
  mux_2831_nl <= MUX_s_1_2_2(nor_601_cse, nor_603_nl, fsm_output(0));
  mux_2833_nl <= MUX_s_1_2_2(mux_2832_nl, mux_2831_nl, fsm_output(1));
  twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2833_nl AND and_dcpl_268;
  nor_593_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(3))));
  nor_594_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (NOT (fsm_output(3))));
  mux_2837_nl <= MUX_s_1_2_2(nor_593_nl, nor_594_nl, fsm_output(0));
  nor_595_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(3)));
  nor_596_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)));
  mux_2836_nl <= MUX_s_1_2_2(nor_595_nl, nor_596_nl, fsm_output(0));
  mux_2838_nl <= MUX_s_1_2_2(mux_2837_nl, mux_2836_nl, fsm_output(2));
  nor_597_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  nor_598_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(3)));
  nor_599_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011100"))
      OR (fsm_output(3)));
  mux_2834_nl <= MUX_s_1_2_2(nor_598_nl, nor_599_nl, fsm_output(0));
  mux_2835_nl <= MUX_s_1_2_2(nor_597_nl, mux_2834_nl, fsm_output(2));
  mux_2839_nl <= MUX_s_1_2_2(mux_2838_nl, mux_2835_nl, fsm_output(1));
  twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2839_nl AND and_dcpl_268;
  nor_590_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_589_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("01110"))
      OR nand_191_cse);
  mux_2841_nl <= MUX_s_1_2_2(nor_589_nl, nor_590_cse, fsm_output(0));
  nor_592_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011101"))
      OR (fsm_output(3)));
  mux_2840_nl <= MUX_s_1_2_2(nor_590_cse, nor_592_nl, fsm_output(0));
  mux_2842_nl <= MUX_s_1_2_2(mux_2841_nl, mux_2840_nl, fsm_output(1));
  twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2842_nl AND and_dcpl_268;
  nor_585_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(3)));
  nor_584_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01111"))
      OR (fsm_output(3)));
  nor_583_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2845_nl <= MUX_s_1_2_2(nor_584_cse, nor_585_cse, fsm_output(0));
  mux_2846_nl <= MUX_s_1_2_2(nor_583_nl, mux_2845_nl, fsm_output(2));
  nor_586_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2843_nl <= MUX_s_1_2_2(nor_585_cse, nor_584_cse, fsm_output(0));
  mux_2844_nl <= MUX_s_1_2_2(nor_586_nl, mux_2843_nl, fsm_output(2));
  mux_2847_nl <= MUX_s_1_2_2(mux_2846_nl, mux_2844_nl, fsm_output(1));
  twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2847_nl AND and_dcpl_268;
  and_533_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("011111")) AND
      CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  nor_581_nl <= NOT((fsm_output(2)) OR (z_out_7(5)) OR (NOT(CONV_SL_1_1(z_out_7(4
      DOWNTO 0)=STD_LOGIC_VECTOR'("11111")) AND (fsm_output(3)))));
  mux_2849_nl <= MUX_s_1_2_2(nor_581_nl, and_533_cse, fsm_output(0));
  nor_582_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("011111"))
      OR (fsm_output(3)));
  mux_2848_nl <= MUX_s_1_2_2(and_533_cse, nor_582_nl, fsm_output(0));
  mux_2850_nl <= MUX_s_1_2_2(mux_2849_nl, mux_2848_nl, fsm_output(1));
  twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2850_nl AND and_dcpl_268;
  nor_576_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)));
  nor_573_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR nand_174_cse);
  nor_574_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000"))
      OR nand_175_cse);
  mux_2855_nl <= MUX_s_1_2_2(nor_573_nl, nor_574_nl, fsm_output(0));
  nor_575_nl <= NOT(CONV_SL_1_1(z_out_8(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR
      (fsm_output(3)));
  mux_2854_nl <= MUX_s_1_2_2(nor_575_nl, nor_576_cse, fsm_output(0));
  mux_2856_nl <= MUX_s_1_2_2(mux_2855_nl, mux_2854_nl, fsm_output(1));
  nor_577_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10000"))
      OR (fsm_output(3)));
  mux_2852_nl <= MUX_s_1_2_2(nor_577_nl, nor_576_cse, fsm_output(0));
  nor_579_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(3)));
  nor_580_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100000"))
      OR (fsm_output(3)));
  mux_2851_nl <= MUX_s_1_2_2(nor_579_nl, nor_580_nl, fsm_output(0));
  mux_2853_nl <= MUX_s_1_2_2(mux_2852_nl, mux_2851_nl, fsm_output(1));
  mux_2857_nl <= MUX_s_1_2_2(mux_2856_nl, mux_2853_nl, fsm_output(2));
  twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2857_nl AND and_dcpl_268;
  nor_570_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_569_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("10000"))
      OR nand_191_cse);
  mux_2859_nl <= MUX_s_1_2_2(nor_569_nl, nor_570_cse, fsm_output(0));
  nor_572_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100001"))
      OR (fsm_output(3)));
  mux_2858_nl <= MUX_s_1_2_2(nor_570_cse, nor_572_nl, fsm_output(0));
  mux_2860_nl <= MUX_s_1_2_2(mux_2859_nl, mux_2858_nl, fsm_output(1));
  twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2860_nl AND and_dcpl_268;
  nor_565_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(3)));
  nor_564_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10001"))
      OR (fsm_output(3)));
  nor_563_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2863_nl <= MUX_s_1_2_2(nor_564_cse, nor_565_cse, fsm_output(0));
  mux_2864_nl <= MUX_s_1_2_2(nor_563_nl, mux_2863_nl, fsm_output(2));
  nor_566_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2861_nl <= MUX_s_1_2_2(nor_565_cse, nor_564_cse, fsm_output(0));
  mux_2862_nl <= MUX_s_1_2_2(nor_566_nl, mux_2861_nl, fsm_output(2));
  mux_2865_nl <= MUX_s_1_2_2(mux_2864_nl, mux_2862_nl, fsm_output(1));
  twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2865_nl AND and_dcpl_268;
  nor_560_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_559_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("1000"))
      OR nand_190_cse);
  mux_2867_nl <= MUX_s_1_2_2(nor_559_nl, nor_560_cse, fsm_output(0));
  nor_562_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100011"))
      OR (fsm_output(3)));
  mux_2866_nl <= MUX_s_1_2_2(nor_560_cse, nor_562_nl, fsm_output(0));
  mux_2868_nl <= MUX_s_1_2_2(mux_2867_nl, mux_2866_nl, fsm_output(1));
  twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2868_nl AND and_dcpl_268;
  nor_552_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(3))));
  nor_553_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (NOT (fsm_output(3))));
  mux_2872_nl <= MUX_s_1_2_2(nor_552_nl, nor_553_nl, fsm_output(0));
  nor_554_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(3)));
  nor_555_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)));
  mux_2871_nl <= MUX_s_1_2_2(nor_554_nl, nor_555_nl, fsm_output(0));
  mux_2873_nl <= MUX_s_1_2_2(mux_2872_nl, mux_2871_nl, fsm_output(2));
  nor_556_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  nor_557_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(3)));
  nor_558_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"))
      OR (fsm_output(3)));
  mux_2869_nl <= MUX_s_1_2_2(nor_557_nl, nor_558_nl, fsm_output(0));
  mux_2870_nl <= MUX_s_1_2_2(nor_556_nl, mux_2869_nl, fsm_output(2));
  mux_2874_nl <= MUX_s_1_2_2(mux_2873_nl, mux_2870_nl, fsm_output(1));
  twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2874_nl AND and_dcpl_268;
  nor_549_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_548_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("10010"))
      OR nand_191_cse);
  mux_2876_nl <= MUX_s_1_2_2(nor_548_nl, nor_549_cse, fsm_output(0));
  nor_551_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100101"))
      OR (fsm_output(3)));
  mux_2875_nl <= MUX_s_1_2_2(nor_549_cse, nor_551_nl, fsm_output(0));
  mux_2877_nl <= MUX_s_1_2_2(mux_2876_nl, mux_2875_nl, fsm_output(1));
  twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2877_nl AND and_dcpl_268;
  nor_544_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(3)));
  nor_543_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10011"))
      OR (fsm_output(3)));
  nor_542_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2880_nl <= MUX_s_1_2_2(nor_543_cse, nor_544_cse, fsm_output(0));
  mux_2881_nl <= MUX_s_1_2_2(nor_542_nl, mux_2880_nl, fsm_output(2));
  nor_545_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2878_nl <= MUX_s_1_2_2(nor_544_cse, nor_543_cse, fsm_output(0));
  mux_2879_nl <= MUX_s_1_2_2(nor_545_nl, mux_2878_nl, fsm_output(2));
  mux_2882_nl <= MUX_s_1_2_2(mux_2881_nl, mux_2879_nl, fsm_output(1));
  twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2882_nl AND and_dcpl_268;
  nor_539_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_538_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("100"))
      OR nand_188_cse);
  mux_2884_nl <= MUX_s_1_2_2(nor_538_nl, nor_539_cse, fsm_output(0));
  nor_541_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100111"))
      OR (fsm_output(3)));
  mux_2883_nl <= MUX_s_1_2_2(nor_539_cse, nor_541_nl, fsm_output(0));
  mux_2885_nl <= MUX_s_1_2_2(mux_2884_nl, mux_2883_nl, fsm_output(1));
  twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2885_nl AND and_dcpl_268;
  nor_533_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)));
  nor_530_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR nand_174_cse);
  nor_531_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("01000"))
      OR nand_175_cse);
  mux_2890_nl <= MUX_s_1_2_2(nor_530_nl, nor_531_nl, fsm_output(0));
  nor_532_nl <= NOT(CONV_SL_1_1(z_out_8(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR
      (fsm_output(3)));
  mux_2889_nl <= MUX_s_1_2_2(nor_532_nl, nor_533_cse, fsm_output(0));
  mux_2891_nl <= MUX_s_1_2_2(mux_2890_nl, mux_2889_nl, fsm_output(1));
  nor_534_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10100"))
      OR (fsm_output(3)));
  mux_2887_nl <= MUX_s_1_2_2(nor_534_nl, nor_533_cse, fsm_output(0));
  nor_536_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(3)));
  nor_537_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101000"))
      OR (fsm_output(3)));
  mux_2886_nl <= MUX_s_1_2_2(nor_536_nl, nor_537_nl, fsm_output(0));
  mux_2888_nl <= MUX_s_1_2_2(mux_2887_nl, mux_2886_nl, fsm_output(1));
  mux_2892_nl <= MUX_s_1_2_2(mux_2891_nl, mux_2888_nl, fsm_output(2));
  twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2892_nl AND and_dcpl_268;
  nor_527_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_526_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("10100"))
      OR nand_191_cse);
  mux_2894_nl <= MUX_s_1_2_2(nor_526_nl, nor_527_cse, fsm_output(0));
  nor_529_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101001"))
      OR (fsm_output(3)));
  mux_2893_nl <= MUX_s_1_2_2(nor_527_cse, nor_529_nl, fsm_output(0));
  mux_2895_nl <= MUX_s_1_2_2(mux_2894_nl, mux_2893_nl, fsm_output(1));
  twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2895_nl AND and_dcpl_268;
  nor_522_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(3)));
  nor_521_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10101"))
      OR (fsm_output(3)));
  nor_520_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2898_nl <= MUX_s_1_2_2(nor_521_cse, nor_522_cse, fsm_output(0));
  mux_2899_nl <= MUX_s_1_2_2(nor_520_nl, mux_2898_nl, fsm_output(2));
  nor_523_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2896_nl <= MUX_s_1_2_2(nor_522_cse, nor_521_cse, fsm_output(0));
  mux_2897_nl <= MUX_s_1_2_2(nor_523_nl, mux_2896_nl, fsm_output(2));
  mux_2900_nl <= MUX_s_1_2_2(mux_2899_nl, mux_2897_nl, fsm_output(1));
  twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2900_nl AND and_dcpl_268;
  nor_517_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_516_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("1010"))
      OR nand_190_cse);
  mux_2902_nl <= MUX_s_1_2_2(nor_516_nl, nor_517_cse, fsm_output(0));
  nor_519_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101011"))
      OR (fsm_output(3)));
  mux_2901_nl <= MUX_s_1_2_2(nor_517_cse, nor_519_nl, fsm_output(0));
  mux_2903_nl <= MUX_s_1_2_2(mux_2902_nl, mux_2901_nl, fsm_output(1));
  twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2903_nl AND and_dcpl_268;
  nor_509_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(3))));
  nor_510_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (NOT (fsm_output(3))));
  mux_2907_nl <= MUX_s_1_2_2(nor_509_nl, nor_510_nl, fsm_output(0));
  nor_511_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(3)));
  nor_512_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)));
  mux_2906_nl <= MUX_s_1_2_2(nor_511_nl, nor_512_nl, fsm_output(0));
  mux_2908_nl <= MUX_s_1_2_2(mux_2907_nl, mux_2906_nl, fsm_output(2));
  nor_513_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  nor_514_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(3)));
  nor_515_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101100"))
      OR (fsm_output(3)));
  mux_2904_nl <= MUX_s_1_2_2(nor_514_nl, nor_515_nl, fsm_output(0));
  mux_2905_nl <= MUX_s_1_2_2(nor_513_nl, mux_2904_nl, fsm_output(2));
  mux_2909_nl <= MUX_s_1_2_2(mux_2908_nl, mux_2905_nl, fsm_output(1));
  twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2909_nl AND and_dcpl_268;
  nor_506_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_505_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("10110"))
      OR nand_191_cse);
  mux_2911_nl <= MUX_s_1_2_2(nor_505_nl, nor_506_cse, fsm_output(0));
  nor_508_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101101"))
      OR (fsm_output(3)));
  mux_2910_nl <= MUX_s_1_2_2(nor_506_cse, nor_508_nl, fsm_output(0));
  mux_2912_nl <= MUX_s_1_2_2(mux_2911_nl, mux_2910_nl, fsm_output(1));
  twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2912_nl AND and_dcpl_268;
  nor_501_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(3)));
  nor_500_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("10111"))
      OR (fsm_output(3)));
  nor_499_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2915_nl <= MUX_s_1_2_2(nor_500_cse, nor_501_cse, fsm_output(0));
  mux_2916_nl <= MUX_s_1_2_2(nor_499_nl, mux_2915_nl, fsm_output(2));
  nor_502_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2913_nl <= MUX_s_1_2_2(nor_501_cse, nor_500_cse, fsm_output(0));
  mux_2914_nl <= MUX_s_1_2_2(nor_502_nl, mux_2913_nl, fsm_output(2));
  mux_2917_nl <= MUX_s_1_2_2(mux_2916_nl, mux_2914_nl, fsm_output(1));
  twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2917_nl AND and_dcpl_268;
  and_531_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("101111")) AND
      CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  nor_497_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10"))
      OR nand_184_cse);
  mux_2919_nl <= MUX_s_1_2_2(nor_497_nl, and_531_cse, fsm_output(0));
  nor_498_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("101111"))
      OR (fsm_output(3)));
  mux_2918_nl <= MUX_s_1_2_2(and_531_cse, nor_498_nl, fsm_output(0));
  mux_2920_nl <= MUX_s_1_2_2(mux_2919_nl, mux_2918_nl, fsm_output(1));
  twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2920_nl AND and_dcpl_268;
  nor_492_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)));
  nor_489_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)))));
  nor_490_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(3)))));
  mux_2925_nl <= MUX_s_1_2_2(nor_489_nl, nor_490_nl, fsm_output(0));
  nor_491_nl <= NOT(CONV_SL_1_1(z_out_8(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR
      (fsm_output(3)));
  mux_2924_nl <= MUX_s_1_2_2(nor_491_nl, nor_492_cse, fsm_output(0));
  mux_2926_nl <= MUX_s_1_2_2(mux_2925_nl, mux_2924_nl, fsm_output(1));
  nor_493_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11000"))
      OR (fsm_output(3)));
  mux_2922_nl <= MUX_s_1_2_2(nor_493_nl, nor_492_cse, fsm_output(0));
  nor_495_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(3)));
  nor_496_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110000"))
      OR (fsm_output(3)));
  mux_2921_nl <= MUX_s_1_2_2(nor_495_nl, nor_496_nl, fsm_output(0));
  mux_2923_nl <= MUX_s_1_2_2(mux_2922_nl, mux_2921_nl, fsm_output(1));
  mux_2927_nl <= MUX_s_1_2_2(mux_2926_nl, mux_2923_nl, fsm_output(2));
  twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2927_nl AND and_dcpl_268;
  nor_486_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_485_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("11000"))
      OR nand_191_cse);
  mux_2929_nl <= MUX_s_1_2_2(nor_485_nl, nor_486_cse, fsm_output(0));
  nor_488_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110001"))
      OR (fsm_output(3)));
  mux_2928_nl <= MUX_s_1_2_2(nor_486_cse, nor_488_nl, fsm_output(0));
  mux_2930_nl <= MUX_s_1_2_2(mux_2929_nl, mux_2928_nl, fsm_output(1));
  twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2930_nl AND and_dcpl_268;
  nor_481_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(3)));
  nor_480_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11001"))
      OR (fsm_output(3)));
  nor_479_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2933_nl <= MUX_s_1_2_2(nor_480_cse, nor_481_cse, fsm_output(0));
  mux_2934_nl <= MUX_s_1_2_2(nor_479_nl, mux_2933_nl, fsm_output(2));
  nor_482_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2931_nl <= MUX_s_1_2_2(nor_481_cse, nor_480_cse, fsm_output(0));
  mux_2932_nl <= MUX_s_1_2_2(nor_482_nl, mux_2931_nl, fsm_output(2));
  mux_2935_nl <= MUX_s_1_2_2(mux_2934_nl, mux_2932_nl, fsm_output(1));
  twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2935_nl AND and_dcpl_268;
  nor_476_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_475_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("1100"))
      OR nand_190_cse);
  mux_2937_nl <= MUX_s_1_2_2(nor_475_nl, nor_476_cse, fsm_output(0));
  nor_478_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110011"))
      OR (fsm_output(3)));
  mux_2936_nl <= MUX_s_1_2_2(nor_476_cse, nor_478_nl, fsm_output(0));
  mux_2938_nl <= MUX_s_1_2_2(mux_2937_nl, mux_2936_nl, fsm_output(1));
  twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2938_nl AND and_dcpl_268;
  nor_468_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(3))));
  nor_469_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (NOT (fsm_output(3))));
  mux_2942_nl <= MUX_s_1_2_2(nor_468_nl, nor_469_nl, fsm_output(0));
  nor_470_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(3)));
  nor_471_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)));
  mux_2941_nl <= MUX_s_1_2_2(nor_470_nl, nor_471_nl, fsm_output(0));
  mux_2943_nl <= MUX_s_1_2_2(mux_2942_nl, mux_2941_nl, fsm_output(2));
  nor_472_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  nor_473_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(3)));
  nor_474_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110100"))
      OR (fsm_output(3)));
  mux_2939_nl <= MUX_s_1_2_2(nor_473_nl, nor_474_nl, fsm_output(0));
  mux_2940_nl <= MUX_s_1_2_2(nor_472_nl, mux_2939_nl, fsm_output(2));
  mux_2944_nl <= MUX_s_1_2_2(mux_2943_nl, mux_2940_nl, fsm_output(1));
  twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2944_nl AND and_dcpl_268;
  nor_465_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_464_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("11010"))
      OR nand_191_cse);
  mux_2946_nl <= MUX_s_1_2_2(nor_464_nl, nor_465_cse, fsm_output(0));
  nor_467_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110101"))
      OR (fsm_output(3)));
  mux_2945_nl <= MUX_s_1_2_2(nor_465_cse, nor_467_nl, fsm_output(0));
  mux_2947_nl <= MUX_s_1_2_2(mux_2946_nl, mux_2945_nl, fsm_output(1));
  twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2947_nl AND and_dcpl_268;
  nor_460_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(3)));
  nor_459_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11011"))
      OR (fsm_output(3)));
  nor_458_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2950_nl <= MUX_s_1_2_2(nor_459_cse, nor_460_cse, fsm_output(0));
  mux_2951_nl <= MUX_s_1_2_2(nor_458_nl, mux_2950_nl, fsm_output(2));
  nor_461_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2948_nl <= MUX_s_1_2_2(nor_460_cse, nor_459_cse, fsm_output(0));
  mux_2949_nl <= MUX_s_1_2_2(nor_461_nl, mux_2948_nl, fsm_output(2));
  mux_2952_nl <= MUX_s_1_2_2(mux_2951_nl, mux_2949_nl, fsm_output(1));
  twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2952_nl AND and_dcpl_268;
  and_529_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("110111")) AND
      CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  nor_456_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("110"))
      OR nand_188_cse);
  mux_2954_nl <= MUX_s_1_2_2(nor_456_nl, and_529_cse, fsm_output(0));
  nor_457_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("110111"))
      OR (fsm_output(3)));
  mux_2953_nl <= MUX_s_1_2_2(and_529_cse, nor_457_nl, fsm_output(0));
  mux_2955_nl <= MUX_s_1_2_2(mux_2954_nl, mux_2953_nl, fsm_output(1));
  twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2955_nl AND and_dcpl_268;
  nor_451_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)));
  nor_449_nl <= NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)))));
  nor_450_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 3)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(3)))));
  mux_2960_nl <= MUX_s_1_2_2(nor_449_nl, nor_450_nl, fsm_output(0));
  and_528_nl <= CONV_SL_1_1(z_out_8(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (NOT
      (fsm_output(3)));
  mux_2959_nl <= MUX_s_1_2_2(and_528_nl, nor_451_cse, fsm_output(0));
  mux_2961_nl <= MUX_s_1_2_2(mux_2960_nl, mux_2959_nl, fsm_output(1));
  nor_452_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11100"))
      OR (fsm_output(3)));
  mux_2957_nl <= MUX_s_1_2_2(nor_452_nl, nor_451_cse, fsm_output(0));
  nor_454_nl <= NOT(CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(3)));
  nor_455_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111000"))
      OR (fsm_output(3)));
  mux_2956_nl <= MUX_s_1_2_2(nor_454_nl, nor_455_nl, fsm_output(0));
  mux_2958_nl <= MUX_s_1_2_2(mux_2957_nl, mux_2956_nl, fsm_output(1));
  mux_2962_nl <= MUX_s_1_2_2(mux_2961_nl, mux_2958_nl, fsm_output(2));
  twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2962_nl AND and_dcpl_268;
  nor_446_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")));
  nor_445_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("11100"))
      OR nand_191_cse);
  mux_2964_nl <= MUX_s_1_2_2(nor_445_nl, nor_446_cse, fsm_output(0));
  nor_448_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111001"))
      OR (fsm_output(3)));
  mux_2963_nl <= MUX_s_1_2_2(nor_446_cse, nor_448_nl, fsm_output(0));
  mux_2965_nl <= MUX_s_1_2_2(mux_2964_nl, mux_2963_nl, fsm_output(1));
  twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2965_nl AND and_dcpl_268;
  nor_441_cse <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(3)));
  nor_440_cse <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11101"))
      OR (fsm_output(3)));
  nor_439_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(3))));
  mux_2968_nl <= MUX_s_1_2_2(nor_440_cse, nor_441_cse, fsm_output(0));
  mux_2969_nl <= MUX_s_1_2_2(nor_439_nl, mux_2968_nl, fsm_output(2));
  nor_442_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  mux_2966_nl <= MUX_s_1_2_2(nor_441_cse, nor_440_cse, fsm_output(0));
  mux_2967_nl <= MUX_s_1_2_2(nor_442_nl, mux_2966_nl, fsm_output(2));
  mux_2970_nl <= MUX_s_1_2_2(mux_2969_nl, mux_2967_nl, fsm_output(1));
  twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2970_nl AND and_dcpl_268;
  and_526_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111011")) AND
      CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  nor_437_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 2)/=STD_LOGIC_VECTOR'("1110"))
      OR nand_190_cse);
  mux_2972_nl <= MUX_s_1_2_2(nor_437_nl, and_526_cse, fsm_output(0));
  nor_438_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111011"))
      OR (fsm_output(3)));
  mux_2971_nl <= MUX_s_1_2_2(and_526_cse, nor_438_nl, fsm_output(0));
  mux_2973_nl <= MUX_s_1_2_2(mux_2972_nl, mux_2971_nl, fsm_output(1));
  twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2973_nl AND and_dcpl_268;
  and_789_nl <= CONV_SL_1_1(COMP_LOOP_3_tmp_lshift_ncse_sva(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11110"))
      AND (fsm_output(3));
  and_810_nl <= CONV_SL_1_1(COMP_LOOP_2_tmp_lshift_ncse_sva(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111100"))
      AND (fsm_output(3));
  mux_2977_nl <= MUX_s_1_2_2(and_789_nl, and_810_nl, fsm_output(0));
  nor_433_nl <= NOT(CONV_SL_1_1(z_out_7(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("11110"))
      OR (fsm_output(3)));
  nor_434_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)));
  mux_2976_nl <= MUX_s_1_2_2(nor_433_nl, nor_434_nl, fsm_output(0));
  mux_2978_nl <= MUX_s_1_2_2(mux_2977_nl, mux_2976_nl, fsm_output(2));
  nor_435_nl <= NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(3)));
  and_525_nl <= CONV_SL_1_1(COMP_LOOP_5_tmp_mul_idiv_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(3)));
  nor_436_nl <= NOT(CONV_SL_1_1(COMP_LOOP_2_tmp_mul_idiv_sva(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100"))
      OR (fsm_output(3)));
  mux_2974_nl <= MUX_s_1_2_2(and_525_nl, nor_436_nl, fsm_output(0));
  mux_2975_nl <= MUX_s_1_2_2(nor_435_nl, mux_2974_nl, fsm_output(2));
  mux_2979_nl <= MUX_s_1_2_2(mux_2978_nl, mux_2975_nl, fsm_output(1));
  twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2979_nl AND and_dcpl_268;
  and_523_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101")) AND
      CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  nor_429_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("11110"))
      OR nand_191_cse);
  mux_2981_nl <= MUX_s_1_2_2(nor_429_nl, and_523_cse, fsm_output(0));
  nor_430_nl <= NOT((fsm_output(2)) OR CONV_SL_1_1(z_out_7(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111101"))
      OR (fsm_output(3)));
  mux_2980_nl <= MUX_s_1_2_2(and_523_cse, nor_430_nl, fsm_output(0));
  mux_2982_nl <= MUX_s_1_2_2(mux_2981_nl, mux_2980_nl, fsm_output(1));
  twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2982_nl AND and_dcpl_268;
  and_519_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110")) AND
      (NOT (fsm_output(3)));
  and_518_cse <= CONV_SL_1_1(z_out_7(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111")) AND
      (NOT (fsm_output(3)));
  and_790_nl <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110")) AND
      (NOT (fsm_output(0))) AND (fsm_output(3));
  mux_2985_nl <= MUX_s_1_2_2(and_518_cse, and_519_cse, fsm_output(0));
  mux_2986_nl <= MUX_s_1_2_2(and_790_nl, mux_2985_nl, fsm_output(2));
  and_520_nl <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111110")) AND
      (fsm_output(0)) AND (NOT (fsm_output(3)));
  mux_2983_nl <= MUX_s_1_2_2(and_519_cse, and_518_cse, fsm_output(0));
  mux_2984_nl <= MUX_s_1_2_2(and_520_nl, mux_2983_nl, fsm_output(2));
  mux_2987_nl <= MUX_s_1_2_2(mux_2986_nl, mux_2984_nl, fsm_output(1));
  twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2987_nl AND and_dcpl_268;
  and_515_cse <= CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111")) AND
      CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("01"));
  nor_427_nl <= NOT((fsm_output(2)) OR (NOT(CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (fsm_output(3)))));
  mux_2989_nl <= MUX_s_1_2_2(nor_427_nl, and_515_cse, fsm_output(0));
  and_517_nl <= (NOT (fsm_output(2))) AND CONV_SL_1_1(z_out_7(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111111"))
      AND (NOT (fsm_output(3)));
  mux_2988_nl <= MUX_s_1_2_2(and_515_cse, and_517_nl, fsm_output(0));
  mux_2990_nl <= MUX_s_1_2_2(mux_2989_nl, mux_2988_nl, fsm_output(1));
  twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d <= mux_2990_nl AND and_dcpl_268;
  nor_1716_cse <= NOT((fsm_output(7)) OR (fsm_output(5)));
  nor_1715_cse <= NOT((fsm_output(3)) OR (fsm_output(6)));
  and_dcpl_477 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_488 <= (NOT (fsm_output(4))) AND (fsm_output(0)) AND (NOT (fsm_output(3)))
      AND (fsm_output(6)) AND and_dcpl_477 AND (fsm_output(7)) AND (fsm_output(5));
  and_dcpl_501 <= NOT(CONV_SL_1_1(fsm_output/=STD_LOGIC_VECTOR'("00000010")));
  and_dcpl_503 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_509 <= (NOT (fsm_output(7))) AND (fsm_output(5));
  and_dcpl_513 <= and_dcpl_503 AND and_dcpl_509;
  and_dcpl_514 <= (fsm_output(3)) AND (NOT (fsm_output(6)));
  and_903_cse <= and_dcpl_80 AND and_dcpl_514 AND and_dcpl_513;
  and_dcpl_519 <= (fsm_output(3)) AND (fsm_output(6));
  and_907_cse <= and_dcpl_80 AND and_dcpl_519 AND nor_1744_cse AND nor_1716_cse;
  and_910_cse <= and_dcpl_80 AND (NOT (fsm_output(3))) AND (fsm_output(6)) AND and_dcpl_513;
  and_dcpl_526 <= nor_1744_cse AND (fsm_output(7)) AND (NOT (fsm_output(5)));
  and_914_cse <= and_dcpl_80 AND nor_1715_cse AND and_dcpl_526;
  and_918_cse <= and_dcpl_58 AND and_dcpl_514 AND and_dcpl_503 AND (fsm_output(7))
      AND (fsm_output(5));
  and_920_cse <= and_dcpl_58 AND and_dcpl_519 AND and_dcpl_526;
  and_dcpl_570 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01")) AND
      nor_1716_cse;
  and_dcpl_573 <= and_dcpl_58 AND nor_1715_cse;
  and_dcpl_574 <= and_dcpl_573 AND and_dcpl_570;
  and_dcpl_576 <= (NOT (fsm_output(4))) AND (fsm_output(0)) AND nor_1715_cse;
  and_dcpl_577 <= and_dcpl_576 AND and_dcpl_570;
  and_dcpl_579 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10")) AND
      nor_1716_cse;
  and_dcpl_580 <= and_dcpl_576 AND and_dcpl_579;
  and_dcpl_582 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND
      nor_1716_cse;
  and_dcpl_583 <= and_dcpl_573 AND and_dcpl_582;
  and_dcpl_588 <= and_dcpl_58 AND (fsm_output(3)) AND (NOT (fsm_output(6))) AND (NOT
      (fsm_output(2))) AND (NOT (fsm_output(1))) AND nor_1716_cse;
  and_dcpl_589 <= and_dcpl_573 AND and_dcpl_579;
  and_dcpl_590 <= and_dcpl_576 AND and_dcpl_582;
  and_dcpl_599 <= nor_1744_cse AND nor_1716_cse;
  and_dcpl_602 <= and_dcpl_80 AND nor_1715_cse AND and_dcpl_599;
  and_dcpl_605 <= and_dcpl_503 AND (NOT (fsm_output(7))) AND (fsm_output(5));
  and_dcpl_608 <= and_dcpl_58 AND and_dcpl_514 AND and_dcpl_605;
  and_dcpl_611 <= and_dcpl_58 AND (fsm_output(3)) AND (fsm_output(6)) AND and_dcpl_599;
  and_dcpl_612 <= (NOT (fsm_output(3))) AND (fsm_output(6));
  and_dcpl_614 <= and_dcpl_58 AND and_dcpl_612 AND and_dcpl_605;
  and_dcpl_615 <= (fsm_output(7)) AND (NOT (fsm_output(5)));
  and_dcpl_617 <= and_dcpl_573 AND nor_1744_cse AND and_dcpl_615;
  and_dcpl_618 <= and_dcpl_503 AND and_dcpl_615;
  and_dcpl_619 <= and_dcpl_80 AND and_dcpl_514;
  and_dcpl_620 <= and_dcpl_619 AND and_dcpl_618;
  and_dcpl_623 <= and_dcpl_619 AND nor_1744_cse AND (fsm_output(7)) AND (fsm_output(5));
  and_dcpl_625 <= and_dcpl_80 AND and_dcpl_612 AND and_dcpl_618;
  and_dcpl_632 <= and_dcpl_573 AND and_dcpl_503 AND nor_1716_cse;
  and_dcpl_636 <= and_dcpl_573 AND nor_1744_cse AND and_dcpl_509;
  COMP_LOOP_or_65_itm <= (and_dcpl_58 AND nor_1715_cse AND nor_1744_cse AND and_dcpl_509)
      OR and_903_cse OR and_907_cse OR and_910_cse OR and_914_cse OR and_918_cse
      OR and_920_cse;
  COMP_LOOP_tmp_or_83_itm <= and_dcpl_589 OR and_dcpl_590;
  COMP_LOOP_tmp_or_54_ssc <= and_dcpl_580 OR and_dcpl_583 OR and_dcpl_588;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((and_dcpl_60 AND and_dcpl_57) OR STAGE_LOOP_i_3_0_sva_mx0c1) = '1' )
          THEN
        STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "1010"), z_out_4,
            STAGE_LOOP_i_3_0_sva_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_1423_nl, mux_789_nl, fsm_output(5))) = '1' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_vec_rsc_triosy_0_63_obj_ld_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        COMP_LOOP_1_tmp_mul_idiv_sva_2_0 <= STD_LOGIC_VECTOR'( "000");
        COMP_LOOP_nor_326_itm <= '0';
        COMP_LOOP_nor_319_itm <= '0';
        COMP_LOOP_3_tmp_mul_idiv_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
      ELSE
        reg_vec_rsc_triosy_0_63_obj_ld_cse <= and_dcpl_65 AND (NOT (fsm_output(0)))
            AND (NOT (fsm_output(4))) AND (fsm_output(6)) AND (fsm_output(2)) AND
            (NOT (fsm_output(1))) AND (fsm_output(5)) AND (NOT (z_out_2(4)));
        reg_ensig_cgo_cse <= mux_2997_rmff;
        COMP_LOOP_1_tmp_mul_idiv_sva_2_0 <= z_out_8(2 DOWNTO 0);
        COMP_LOOP_nor_326_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_319_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
        COMP_LOOP_3_tmp_mul_idiv_sva_4_0 <= z_out_7(4 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      tmp_21_sva_2 <= MUX_v_64_2_2(twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_58_i_q_d,
          and_dcpl_263);
      tmp_21_sva_6 <= twiddle_rsc_0_6_i_q_d;
      tmp_21_sva_11 <= MUX_v_64_2_2(twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_30_i_q_d,
          and_dcpl_263);
      tmp_21_sva_13 <= MUX_v_64_2_2(twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_34_i_q_d,
          and_dcpl_263);
      tmp_21_sva_14 <= MUX_v_64_2_2(twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_38_i_q_d,
          and_dcpl_263);
      tmp_21_sva_15 <= MUX_v_64_2_2(twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_42_i_q_d,
          and_dcpl_263);
      tmp_21_sva_17 <= MUX_v_64_2_2(twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_46_i_q_d,
          and_dcpl_263);
      tmp_21_sva_18 <= MUX_v_64_2_2(twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_50_i_q_d,
          and_dcpl_263);
      tmp_21_sva_19 <= MUX_v_64_2_2(twiddle_rsc_0_19_i_q_d, twiddle_rsc_0_54_i_q_d,
          and_dcpl_263);
      tmp_21_sva_21 <= MUX_v_64_2_2(twiddle_rsc_0_21_i_q_d, twiddle_rsc_0_6_i_q_d,
          and_dcpl_263);
      tmp_21_sva_22 <= MUX_v_64_2_2(twiddle_rsc_0_22_i_q_d, twiddle_rsc_0_62_i_q_d,
          and_dcpl_263);
      tmp_21_sva_23 <= MUX_v_64_2_2(twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_10_i_q_d,
          and_dcpl_263);
      tmp_21_sva_25 <= MUX_v_64_2_2(twiddle_rsc_0_25_i_q_d, twiddle_rsc_0_14_i_q_d,
          and_dcpl_263);
      tmp_21_sva_26 <= MUX_v_64_2_2(twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_18_i_q_d,
          and_dcpl_263);
      tmp_21_sva_30 <= twiddle_rsc_0_30_i_q_d;
      tmp_21_sva_34 <= twiddle_rsc_0_34_i_q_d;
      tmp_21_sva_38 <= twiddle_rsc_0_38_i_q_d;
      tmp_21_sva_42 <= twiddle_rsc_0_42_i_q_d;
      tmp_21_sva_46 <= twiddle_rsc_0_46_i_q_d;
      tmp_21_sva_50 <= twiddle_rsc_0_50_i_q_d;
      tmp_21_sva_54 <= twiddle_rsc_0_54_i_q_d;
      tmp_21_sva_58 <= twiddle_rsc_0_58_i_q_d;
      tmp_21_sva_62 <= twiddle_rsc_0_62_i_q_d;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_j_10_0_sva_9_0 <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (VEC_LOOP_j_10_0_sva_9_0_mx0c0 OR (and_dcpl_108 AND and_dcpl_97)) =
          '1' ) THEN
        VEC_LOOP_j_10_0_sva_9_0 <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"),
            (z_out_3(9 DOWNTO 0)), VEC_LOOP_j_not_1_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_422_nl, mux_tmp_720, fsm_output(5))) = '1' ) THEN
        STAGE_LOOP_lshift_psp_sva <= z_out;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(or_4159_nl, nand_493_nl, fsm_output(7))) = '1' ) THEN
        COMP_LOOP_k_10_3_sva_6_0 <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), reg_COMP_LOOP_k_10_3_ftd,
            nand_480_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva <= COMP_LOOP_1_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_psp_sva <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_5_tmp_mul_idiv_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_5_tmp_mul_idiv_sva <= z_out_7(7 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm <= z_out_3(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_1_tmp_acc_cse_sva <= z_out_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1518_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_760_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_761_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_509_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_510_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_258_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_6_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_260_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_261_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_262_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_10_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_264_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_12_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_13_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_14_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_268_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_522_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_270_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_18_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_272_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_20_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_21_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_22_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_23_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_24_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_25_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_26_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_27_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_28_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_29_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_30_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_284_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_285_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_286_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_34_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_288_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_36_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_37_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_38_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_39_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_40_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_41_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_42_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_43_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_44_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_45_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_46_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_47_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_48_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_49_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_50_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_51_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_52_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_53_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_54_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_55_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_56_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_57_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_58_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_59_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_60_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_61_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_62_itm <= '0';
      ELSIF ( mux_3025_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
        COMP_LOOP_COMP_LOOP_and_1518_itm <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva_1(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
            CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva_1(4 DOWNTO 2)=STD_LOGIC_VECTOR'("000"));
        COMP_LOOP_COMP_LOOP_and_760_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000101"));
        COMP_LOOP_COMP_LOOP_and_761_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000110"));
        COMP_LOOP_COMP_LOOP_and_509_itm <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva_1(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT(CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva_1(4
            DOWNTO 2)/=STD_LOGIC_VECTOR'("000")) OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_510_itm <= CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva_1(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
            CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva_1(4 DOWNTO 2)=STD_LOGIC_VECTOR'("000"));
        COMP_LOOP_COMP_LOOP_and_258_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000111"));
        COMP_LOOP_COMP_LOOP_and_6_itm <= CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO
            0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("000"));
        COMP_LOOP_COMP_LOOP_and_260_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001001"));
        COMP_LOOP_COMP_LOOP_and_261_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001010"));
        COMP_LOOP_COMP_LOOP_and_262_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001011"));
        COMP_LOOP_COMP_LOOP_and_10_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(0)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(2))));
        COMP_LOOP_COMP_LOOP_and_264_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001101"));
        COMP_LOOP_COMP_LOOP_and_12_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(0)) AND (VEC_LOOP_j_10_0_sva_9_0(2))
            AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_13_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(0)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_14_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(0)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("00"));
        COMP_LOOP_COMP_LOOP_and_268_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010001"));
        COMP_LOOP_COMP_LOOP_and_522_itm <= (COMP_LOOP_acc_11_psp_sva_1(3)) AND (COMP_LOOP_acc_11_psp_sva_1(0))
            AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT((COMP_LOOP_acc_11_psp_sva_1(4))
            OR (COMP_LOOP_acc_11_psp_sva_1(2)) OR (COMP_LOOP_acc_11_psp_sva_1(1))));
        COMP_LOOP_COMP_LOOP_and_270_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
        COMP_LOOP_COMP_LOOP_and_18_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(1)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2))
            OR (COMP_LOOP_acc_psp_sva_mx0w0(0)) OR (VEC_LOOP_j_10_0_sva_9_0(2))));
        COMP_LOOP_COMP_LOOP_and_272_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
        COMP_LOOP_COMP_LOOP_and_20_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(1)) AND (VEC_LOOP_j_10_0_sva_9_0(2))
            AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2))
            OR (COMP_LOOP_acc_psp_sva_mx0w0(0)) OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_21_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(1)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2))
            OR (COMP_LOOP_acc_psp_sva_mx0w0(0)) OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_22_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(1)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2))
            OR (COMP_LOOP_acc_psp_sva_mx0w0(0))));
        COMP_LOOP_COMP_LOOP_and_23_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2))
            OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))));
        COMP_LOOP_COMP_LOOP_and_24_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
            (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
        COMP_LOOP_COMP_LOOP_and_25_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(1)) AND
            (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2)) OR (VEC_LOOP_j_10_0_sva_9_0(2))
            OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_26_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2))
            OR (VEC_LOOP_j_10_0_sva_9_0(2))));
        COMP_LOOP_COMP_LOOP_and_27_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(2)) AND
            (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))));
        COMP_LOOP_COMP_LOOP_and_28_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(2)) AND
            (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2))
            OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_29_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(2))
            OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_30_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (NOT (COMP_LOOP_acc_psp_sva_mx0w0(2)));
        COMP_LOOP_COMP_LOOP_and_284_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100001"));
        COMP_LOOP_COMP_LOOP_and_285_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100010"));
        COMP_LOOP_COMP_LOOP_and_286_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100011"));
        COMP_LOOP_COMP_LOOP_and_34_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(2))));
        COMP_LOOP_COMP_LOOP_and_288_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100101"));
        COMP_LOOP_COMP_LOOP_and_36_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (VEC_LOOP_j_10_0_sva_9_0(2))
            AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_37_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT(CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_38_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("00"));
        COMP_LOOP_COMP_LOOP_and_39_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (COMP_LOOP_acc_psp_sva_mx0w0(0))
            AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))));
        COMP_LOOP_COMP_LOOP_and_40_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (COMP_LOOP_acc_psp_sva_mx0w0(0))
            AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1))
            OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
        COMP_LOOP_COMP_LOOP_and_41_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (COMP_LOOP_acc_psp_sva_mx0w0(0))
            AND (VEC_LOOP_j_10_0_sva_9_0(1)) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1))
            OR (VEC_LOOP_j_10_0_sva_9_0(2)) OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_42_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (COMP_LOOP_acc_psp_sva_mx0w0(0))
            AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
            AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1)) OR (VEC_LOOP_j_10_0_sva_9_0(2))));
        COMP_LOOP_COMP_LOOP_and_43_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (COMP_LOOP_acc_psp_sva_mx0w0(0))
            AND (VEC_LOOP_j_10_0_sva_9_0(2)) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1))
            OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))));
        COMP_LOOP_COMP_LOOP_and_44_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (COMP_LOOP_acc_psp_sva_mx0w0(0))
            AND (VEC_LOOP_j_10_0_sva_9_0(2)) AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
            (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1)) OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_45_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (COMP_LOOP_acc_psp_sva_mx0w0(0))
            AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
            AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(1)) OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_46_itm <= (COMP_LOOP_acc_psp_sva_mx0w0(2)) AND (COMP_LOOP_acc_psp_sva_mx0w0(0))
            AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
            AND (NOT (COMP_LOOP_acc_psp_sva_mx0w0(1)));
        COMP_LOOP_COMP_LOOP_and_47_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0))
            OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))));
        COMP_LOOP_COMP_LOOP_and_48_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(0)) AND
            (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
        COMP_LOOP_COMP_LOOP_and_49_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(1)) AND
            (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0)) OR (VEC_LOOP_j_10_0_sva_9_0(2))
            OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_50_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0))
            OR (VEC_LOOP_j_10_0_sva_9_0(2))));
        COMP_LOOP_COMP_LOOP_and_51_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(2)) AND
            (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0)) OR CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(1
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))));
        COMP_LOOP_COMP_LOOP_and_52_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (VEC_LOOP_j_10_0_sva_9_0(2)) AND
            (VEC_LOOP_j_10_0_sva_9_0(0)) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0))
            OR (VEC_LOOP_j_10_0_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_53_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT((COMP_LOOP_acc_psp_sva_mx0w0(0))
            OR (VEC_LOOP_j_10_0_sva_9_0(0))));
        COMP_LOOP_COMP_LOOP_and_54_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (NOT (COMP_LOOP_acc_psp_sva_mx0w0(0)));
        COMP_LOOP_COMP_LOOP_and_55_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("000"));
        COMP_LOOP_COMP_LOOP_and_56_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("001"));
        COMP_LOOP_COMP_LOOP_and_57_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("010"));
        COMP_LOOP_COMP_LOOP_and_58_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("011"));
        COMP_LOOP_COMP_LOOP_and_59_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("100"));
        COMP_LOOP_COMP_LOOP_and_60_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("101"));
        COMP_LOOP_COMP_LOOP_and_61_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("110"));
        COMP_LOOP_COMP_LOOP_and_62_itm <= CONV_SL_1_1(COMP_LOOP_acc_psp_sva_mx0w0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND CONV_SL_1_1(VEC_LOOP_j_10_0_sva_9_0(2
            DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_73_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_74_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_75_itm <= '0';
      ELSIF ( COMP_LOOP_or_121_cse = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_73_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_73_nl,
            COMP_LOOP_COMP_LOOP_and_824_nl, and_dcpl_258);
        COMP_LOOP_COMP_LOOP_and_74_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_74_nl,
            COMP_LOOP_COMP_LOOP_and_851_nl, and_dcpl_258);
        COMP_LOOP_COMP_LOOP_and_75_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_75_nl,
            COMP_LOOP_COMP_LOOP_and_858_nl, and_dcpl_258);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_100_itm <= '0';
      ELSIF ( (NOT(mux_3037_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_100_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_100_nl,
            COMP_LOOP_COMP_LOOP_and_323_nl, COMP_LOOP_COMP_LOOP_and_1073_nl, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_261 & and_dcpl_370));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_101_itm <= '0';
      ELSIF ( (mux_3039_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_101_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_101_nl,
            COMP_LOOP_COMP_LOOP_and_348_nl, COMP_LOOP_COMP_LOOP_and_1075_nl, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_259 & and_403_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_102_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_109_itm <= '0';
      ELSIF ( COMP_LOOP_or_126_cse = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_102_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_102_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_78_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse, COMP_LOOP_COMP_LOOP_and_1076_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_112));
        COMP_LOOP_COMP_LOOP_and_109_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_109_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse, COMP_LOOP_COMP_LOOP_and_1094_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_112));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_103_itm <= '0';
      ELSIF ( (NOT(mux_3046_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_103_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_103_nl,
            COMP_LOOP_COMP_LOOP_and_350_nl, COMP_LOOP_COMP_LOOP_and_1079_nl, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_261 & and_dcpl_375));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_104_itm <= '0';
      ELSIF ( (NOT(mux_3047_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_104_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_104_nl,
            COMP_LOOP_COMP_LOOP_and_354_nl, COMP_LOOP_COMP_LOOP_and_1080_nl, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_77 & and_409_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_105_itm <= '0';
      ELSIF ( (NOT(mux_3048_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_105_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_105_nl,
            COMP_LOOP_COMP_LOOP_and_362_nl, COMP_LOOP_COMP_LOOP_and_1082_nl, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_77 & and_dcpl_375));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_106_itm <= '0';
      ELSIF ( (NOT(mux_3053_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_106_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_106_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_79_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse, COMP_LOOP_COMP_LOOP_and_1087_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_411_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_107_itm <= '0';
      ELSIF ( (mux_3059_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_107_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_107_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_cse, COMP_LOOP_COMP_LOOP_and_1088_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_382));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_108_itm <= '0';
      ELSIF ( (NOT(mux_3063_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_108_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_108_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse, COMP_LOOP_COMP_LOOP_and_1090_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_384));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_110_itm <= '0';
      ELSIF ( (mux_3064_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_110_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_110_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_23_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse, COMP_LOOP_COMP_LOOP_and_1103_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_375));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_115_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_117_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_122_itm <= '0';
      ELSIF ( COMP_LOOP_or_135_cse = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_115_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_115_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_27_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_88_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_cse, COMP_LOOP_COMP_LOOP_and_1328_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_86));
        COMP_LOOP_COMP_LOOP_and_117_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_117_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_29_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_90_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_28_cse, COMP_LOOP_COMP_LOOP_and_1332_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_86));
        COMP_LOOP_COMP_LOOP_and_122_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_122_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_33_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_94_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_32_cse, COMP_LOOP_COMP_LOOP_and_1355_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_86));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_116_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_tmp_3003, mux_3073_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_116_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_116_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_28_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_89_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_27_cse, COMP_LOOP_COMP_LOOP_and_1331_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_90));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_118_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3081_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_COMP_LOOP_and_118_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_118_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_30_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_91_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_29_cse, COMP_LOOP_COMP_LOOP_and_1334_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_384));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_119_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3085_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_COMP_LOOP_and_119_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_119_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_244_cse,
            COMP_LOOP_COMP_LOOP_and_1339_nl, STD_LOGIC_VECTOR'( and_dcpl_74 & COMP_LOOP_or_110_rgt
            & and_dcpl_261 & and_dcpl_265));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_120_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3092_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_COMP_LOOP_and_120_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_120_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_31_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_92_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_30_cse, COMP_LOOP_COMP_LOOP_and_1340_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_387));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_121_itm <= '0';
      ELSIF ( (MUX_s_1_2_2((NOT mux_3097_nl), (fsm_output(7)), fsm_output(6))) =
          '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_121_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_121_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_32_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_93_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_31_cse, COMP_LOOP_COMP_LOOP_and_1342_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_370));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_123_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_tmp_3003, mux_742_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_123_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_123_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_95_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_33_cse, COMP_LOOP_COMP_LOOP_and_1356_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_382));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_124_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3102_nl, (fsm_output(7)), fsm_output(6))) = '1' )
          THEN
        COMP_LOOP_COMP_LOOP_and_124_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_124_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_96_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_cse, COMP_LOOP_COMP_LOOP_and_1358_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_115));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_125_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3107_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_COMP_LOOP_and_125_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_125_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_97_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_cse, COMP_LOOP_COMP_LOOP_and_1362_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_388));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3111_nl, and_705_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_14_psp_sva <= COMP_LOOP_acc_14_psp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_3115_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_4_sva <= COMP_LOOP_acc_1_cse_4_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( and_dcpl_390 = '0' ) THEN
        COMP_LOOP_acc_11_psp_sva <= COMP_LOOP_acc_11_psp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( and_dcpl_392 = '0' ) THEN
        COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_3123_nl AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_2_sva <= COMP_LOOP_2_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(mux_3124_nl AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_3_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_5_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_5_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_281_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_nor_281_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_282_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_nor_282_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_284_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_nor_284_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_288_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_nor_288_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_296_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_nor_296_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_333_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_333_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_334_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_334_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_335_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_335_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_336_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_336_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_337_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_337_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_338_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_338_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_339_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_339_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_340_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_340_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_341_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_341_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_342_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_342_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_343_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_343_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_344_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_344_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_345_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_345_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_311_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_nor_311_itm <= NOT(CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_347_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_347_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_349_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_349_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_351_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_351_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_352_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_352_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_353_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_353_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_355_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_355_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_356_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_356_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_357_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_357_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_358_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_358_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_359_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_359_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_360_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_360_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_361_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_361_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_363_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_363_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_364_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_364_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_365_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_365_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_366_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_366_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_367_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_367_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_368_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_368_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_369_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_369_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_370_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_370_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_371_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_371_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_372_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_372_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_373_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_373_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_374_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_374_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_375_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_375_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_376_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_376_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_377_itm <= '0';
      ELSIF ( and_dcpl_396 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_377_itm <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_315_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_315_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_289_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_289_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_313_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_313_itm <= NOT((COMP_LOOP_2_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_2_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_2_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_3_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_3126_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_3_sva <= COMP_LOOP_3_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_3128_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm <= COMP_LOOP_acc_12_nl(8);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_9_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_9_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_505_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_nor_505_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_506_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_nor_506_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_569_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_569_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_508_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_nor_508_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_571_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_571_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_572_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_572_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_573_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_573_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_512_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_nor_512_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_575_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_575_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_576_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_576_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_577_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_577_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_578_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_578_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_579_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_579_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_580_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_580_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_581_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_581_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_520_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_nor_520_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_584_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_584_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_585_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_585_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_586_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_586_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_587_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_587_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_588_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_588_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_589_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_589_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_590_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_590_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_591_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_591_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_592_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_592_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_593_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_593_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_594_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_594_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_595_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_595_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_596_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_596_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_597_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_597_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_535_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_nor_535_itm <= NOT(CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_599_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_599_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_600_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_600_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_601_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_601_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_602_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_602_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_603_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_603_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_604_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_604_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_605_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_605_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_606_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_606_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_607_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_607_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_608_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_608_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_609_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_609_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_610_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_610_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_611_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_611_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_612_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_612_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_613_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_613_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_614_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_614_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_615_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_615_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_616_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_616_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_617_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_617_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_618_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_618_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_619_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_619_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_620_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_620_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_621_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_621_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_622_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_622_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_623_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_623_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_624_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_624_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_625_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_625_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_626_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_626_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_627_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_627_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_628_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_628_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_629_itm <= '0';
      ELSIF ( and_dcpl_399 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_629_itm <= CONV_SL_1_1(COMP_LOOP_3_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_521_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_521_itm <= NOT((COMP_LOOP_3_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_3_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_3_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_3130_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_4_sva <= COMP_LOOP_4_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_3132_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_5_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_13_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_13_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_729_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_nor_729_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_730_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_nor_730_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_821_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_821_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_732_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_nor_732_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_823_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_823_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_825_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_825_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_736_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_nor_736_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_827_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_827_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_828_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_828_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_829_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_829_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_830_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_830_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_831_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_831_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_832_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_832_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_833_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_833_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_744_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_nor_744_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_835_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_835_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_836_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_836_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_837_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_837_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_838_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_838_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_839_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_839_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_840_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_840_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_841_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_841_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_842_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_842_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_843_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_843_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_844_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_844_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_845_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_845_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_846_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_846_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_847_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_847_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_848_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_848_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_849_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_849_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_759_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_nor_759_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_852_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_852_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_853_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_853_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_854_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_854_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_855_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_855_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_856_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_856_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_857_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_857_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_859_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_859_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_860_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_860_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_861_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_861_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_862_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_862_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_863_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_863_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_864_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_864_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_865_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_865_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_866_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_866_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_867_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_867_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_868_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_868_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_869_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_869_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_870_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_870_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_871_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_871_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_872_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_872_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_873_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_873_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_874_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_874_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_875_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_875_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_876_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_876_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_877_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_877_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_878_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_878_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_879_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_879_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_880_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_880_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_881_itm <= '0';
      ELSIF ( and_dcpl_402 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_881_itm <= CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_767_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_767_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_760_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_760_itm <= NOT(CONV_SL_1_1(COMP_LOOP_4_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_734_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_734_itm <= NOT((COMP_LOOP_4_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_4_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_4_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (MUX_s_1_2_2(mux_3140_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0(9
            DOWNTO 2)) + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & '1'), 8));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_5_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3143_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_acc_10_cse_10_1_5_sva <= COMP_LOOP_5_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_3146_nl, (fsm_output(7)), fsm_output(5))) = '1' ) THEN
        COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_6_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_17_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_nor_17_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_953_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_nor_953_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_954_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_nor_954_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_956_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_nor_956_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1077_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1077_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_960_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_nor_960_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1081_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1081_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1083_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1083_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1084_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1084_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1085_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1085_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_968_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_nor_968_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1089_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1089_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1091_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1091_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1092_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1092_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1093_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1093_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1095_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1095_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1096_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1096_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1097_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1097_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1098_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1098_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1099_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1099_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1100_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1100_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1101_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1101_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_983_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_nor_983_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1105_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1105_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1107_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1107_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1108_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1108_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1109_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1109_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1111_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1111_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1112_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1112_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1113_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1113_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1114_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1114_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1115_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1115_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1116_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1116_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1117_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1117_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1119_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1119_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1120_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1120_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1121_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1121_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1122_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1122_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1123_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1123_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1124_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1124_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1125_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1125_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1126_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1126_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111000"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1127_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1127_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111001"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1128_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1128_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111010"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1129_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1129_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1130_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1130_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111100"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1131_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1131_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1132_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1132_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1133_itm <= '0';
      ELSIF ( and_dcpl_403 = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_1133_itm <= CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_970_itm <= '0';
      ELSIF ( and_dcpl_404 = '0' ) THEN
        COMP_LOOP_nor_970_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_969_itm <= '0';
      ELSIF ( (NOT(mux_3152_nl AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_nor_969_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_984_itm <= '0';
      ELSIF ( and_dcpl_406 = '0' ) THEN
        COMP_LOOP_nor_984_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_964_itm <= '0';
      ELSIF ( and_dcpl_406 = '0' ) THEN
        COMP_LOOP_nor_964_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_961_itm <= '0';
      ELSIF ( and_dcpl_406 = '0' ) THEN
        COMP_LOOP_nor_961_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_955_itm <= '0';
      ELSIF ( and_dcpl_407 = '0' ) THEN
        COMP_LOOP_nor_955_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(5
            DOWNTO 2)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_962_itm <= '0';
      ELSIF ( (NOT(mux_3160_nl AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_nor_962_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_957_itm <= '0';
      ELSIF ( (NOT((mux_221_cse XOR (fsm_output(5))) AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_nor_957_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_976_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_976_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_958_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_958_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_998_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_998_itm <= NOT(CONV_SL_1_1(COMP_LOOP_5_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_972_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_972_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_987_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_987_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_985_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_985_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_nor_140_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_nor_140_itm <= COMP_LOOP_tmp_nor_140_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_nor_141_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_nor_141_itm <= COMP_LOOP_tmp_nor_141_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_166_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_166_itm <= CONV_SL_1_1(z_out_7(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
            AND COMP_LOOP_tmp_nor_76_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_nor_143_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_nor_143_itm <= COMP_LOOP_tmp_nor_77_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_168_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_168_itm <= (z_out_7(2)) AND (z_out_7(0))
            AND COMP_LOOP_tmp_nor_78_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_169_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_169_itm <= CONV_SL_1_1(z_out_7(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
            AND COMP_LOOP_tmp_nor_79_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_170_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_170_itm <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_nor_146_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_nor_146_itm <= COMP_LOOP_tmp_nor_80_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_172_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_172_itm <= (z_out_7(3)) AND (z_out_7(0))
            AND COMP_LOOP_tmp_nor_81_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_173_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_173_itm <= (z_out_7(3)) AND (z_out_7(1))
            AND COMP_LOOP_tmp_nor_82_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_itm <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_175_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_175_itm <= CONV_SL_1_1(z_out_7(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
            AND COMP_LOOP_tmp_nor_83_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_176_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_176_itm <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_177_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_177_itm <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_178_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_178_itm <= CONV_SL_1_1(z_out_7(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_991_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_991_itm <= NOT((COMP_LOOP_5_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_5_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_5_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3163_nl, (fsm_output(7)), fsm_output(6))) = '1' )
          THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "101")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_tmp_3102, and_736_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_6_sva <= COMP_LOOP_6_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_tmp_3102, mux_3171_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_7_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_21_itm <= '0';
        COMP_LOOP_nor_1177_itm <= '0';
        COMP_LOOP_nor_1178_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1325_itm <= '0';
        COMP_LOOP_nor_1180_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1327_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1329_itm <= '0';
        COMP_LOOP_nor_1184_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1333_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1335_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1336_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1337_itm <= '0';
        COMP_LOOP_nor_1192_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1341_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1343_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1344_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1345_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1346_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1347_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1348_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1349_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1350_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1351_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1352_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1353_itm <= '0';
        COMP_LOOP_nor_1207_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1357_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1359_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1360_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1361_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1363_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1364_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1365_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1366_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1367_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1368_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1369_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1371_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1372_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1373_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1374_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1375_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1376_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1377_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1378_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1379_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1380_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1381_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1382_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1383_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1384_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1385_itm <= '0';
      ELSIF ( mux_3175_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_21_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
        COMP_LOOP_nor_1177_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_nor_1178_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1325_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000011"));
        COMP_LOOP_nor_1180_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1327_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000101"));
        COMP_LOOP_COMP_LOOP_and_1329_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000111"));
        COMP_LOOP_nor_1184_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1333_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001011"));
        COMP_LOOP_COMP_LOOP_and_1335_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001101"));
        COMP_LOOP_COMP_LOOP_and_1336_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001110"));
        COMP_LOOP_COMP_LOOP_and_1337_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001111"));
        COMP_LOOP_nor_1192_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1341_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
        COMP_LOOP_COMP_LOOP_and_1343_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
        COMP_LOOP_COMP_LOOP_and_1344_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010110"));
        COMP_LOOP_COMP_LOOP_and_1345_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010111"));
        COMP_LOOP_COMP_LOOP_and_1346_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011000"));
        COMP_LOOP_COMP_LOOP_and_1347_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011001"));
        COMP_LOOP_COMP_LOOP_and_1348_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011010"));
        COMP_LOOP_COMP_LOOP_and_1349_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011011"));
        COMP_LOOP_COMP_LOOP_and_1350_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011100"));
        COMP_LOOP_COMP_LOOP_and_1351_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011101"));
        COMP_LOOP_COMP_LOOP_and_1352_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011110"));
        COMP_LOOP_COMP_LOOP_and_1353_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011111"));
        COMP_LOOP_nor_1207_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_COMP_LOOP_and_1357_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100011"));
        COMP_LOOP_COMP_LOOP_and_1359_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100101"));
        COMP_LOOP_COMP_LOOP_and_1360_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100110"));
        COMP_LOOP_COMP_LOOP_and_1361_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100111"));
        COMP_LOOP_COMP_LOOP_and_1363_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101001"));
        COMP_LOOP_COMP_LOOP_and_1364_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101010"));
        COMP_LOOP_COMP_LOOP_and_1365_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101011"));
        COMP_LOOP_COMP_LOOP_and_1366_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101100"));
        COMP_LOOP_COMP_LOOP_and_1367_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101101"));
        COMP_LOOP_COMP_LOOP_and_1368_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101110"));
        COMP_LOOP_COMP_LOOP_and_1369_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101111"));
        COMP_LOOP_COMP_LOOP_and_1371_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110001"));
        COMP_LOOP_COMP_LOOP_and_1372_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110010"));
        COMP_LOOP_COMP_LOOP_and_1373_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110011"));
        COMP_LOOP_COMP_LOOP_and_1374_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110100"));
        COMP_LOOP_COMP_LOOP_and_1375_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110101"));
        COMP_LOOP_COMP_LOOP_and_1376_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110110"));
        COMP_LOOP_COMP_LOOP_and_1377_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110111"));
        COMP_LOOP_COMP_LOOP_and_1378_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111000"));
        COMP_LOOP_COMP_LOOP_and_1379_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111001"));
        COMP_LOOP_COMP_LOOP_and_1380_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111010"));
        COMP_LOOP_COMP_LOOP_and_1381_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111011"));
        COMP_LOOP_COMP_LOOP_and_1382_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111100"));
        COMP_LOOP_COMP_LOOP_and_1383_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
        COMP_LOOP_COMP_LOOP_and_1384_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111110"));
        COMP_LOOP_COMP_LOOP_and_1385_itm <= CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1185_itm <= '0';
      ELSIF ( and_dcpl_410 = '0' ) THEN
        COMP_LOOP_nor_1185_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1211_itm <= '0';
      ELSIF ( and_dcpl_392 = '0' ) THEN
        COMP_LOOP_nor_1211_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1209_itm <= '0';
      ELSIF ( and_dcpl_404 = '0' ) THEN
        COMP_LOOP_nor_1209_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1196_itm <= '0';
      ELSIF ( and_dcpl_407 = '0' ) THEN
        COMP_LOOP_nor_1196_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1208_itm <= '0';
      ELSIF ( and_dcpl_411 = '0' ) THEN
        COMP_LOOP_nor_1208_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1186_itm <= '0';
      ELSIF ( and_dcpl_411 = '0' ) THEN
        COMP_LOOP_nor_1186_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1182_itm <= '0';
      ELSIF ( and_dcpl_411 = '0' ) THEN
        COMP_LOOP_nor_1182_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1222_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_1222_itm <= NOT(CONV_SL_1_1(COMP_LOOP_6_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1188_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_1188_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1215_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_1215_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1194_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_1194_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1193_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_1193_itm <= NOT((COMP_LOOP_6_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_6_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_6_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_7_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_3182_nl, and_705_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_7_sva <= COMP_LOOP_7_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_3185_itm = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm <= COMP_LOOP_acc_15_nl(7);
        reg_COMP_LOOP_k_10_3_ftd <= z_out_2(6 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_25_itm <= '0';
        COMP_LOOP_nor_1401_itm <= '0';
        COMP_LOOP_nor_1402_itm <= '0';
        COMP_LOOP_nor_1404_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1579_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1580_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1581_itm <= '0';
        COMP_LOOP_nor_1408_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1583_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1585_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1586_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1587_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1588_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1589_itm <= '0';
        COMP_LOOP_nor_1416_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1591_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1592_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1593_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1595_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1596_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1597_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1599_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1600_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1601_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1602_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1603_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1604_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1605_itm <= '0';
        COMP_LOOP_nor_1431_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1608_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1609_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1611_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1612_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1613_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1615_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1616_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1617_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1618_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1619_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1620_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1621_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1623_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1624_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1625_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1626_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1627_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1628_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1629_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1630_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1631_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1632_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1633_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1634_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1635_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1636_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1637_itm <= '0';
      ELSIF ( mux_3187_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_25_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
        COMP_LOOP_nor_1401_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_nor_1402_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
        COMP_LOOP_nor_1404_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1579_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000101"));
        COMP_LOOP_COMP_LOOP_and_1580_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000110"));
        COMP_LOOP_COMP_LOOP_and_1581_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000111"));
        COMP_LOOP_nor_1408_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1583_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001001"));
        COMP_LOOP_COMP_LOOP_and_1585_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001011"));
        COMP_LOOP_COMP_LOOP_and_1586_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001100"));
        COMP_LOOP_COMP_LOOP_and_1587_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001101"));
        COMP_LOOP_COMP_LOOP_and_1588_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001110"));
        COMP_LOOP_COMP_LOOP_and_1589_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001111"));
        COMP_LOOP_nor_1416_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1591_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010001"));
        COMP_LOOP_COMP_LOOP_and_1592_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010010"));
        COMP_LOOP_COMP_LOOP_and_1593_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
        COMP_LOOP_COMP_LOOP_and_1595_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
        COMP_LOOP_COMP_LOOP_and_1596_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010110"));
        COMP_LOOP_COMP_LOOP_and_1597_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010111"));
        COMP_LOOP_COMP_LOOP_and_1599_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011001"));
        COMP_LOOP_COMP_LOOP_and_1600_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011010"));
        COMP_LOOP_COMP_LOOP_and_1601_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011011"));
        COMP_LOOP_COMP_LOOP_and_1602_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011100"));
        COMP_LOOP_COMP_LOOP_and_1603_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011101"));
        COMP_LOOP_COMP_LOOP_and_1604_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011110"));
        COMP_LOOP_COMP_LOOP_and_1605_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011111"));
        COMP_LOOP_nor_1431_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_COMP_LOOP_and_1608_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100010"));
        COMP_LOOP_COMP_LOOP_and_1609_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100011"));
        COMP_LOOP_COMP_LOOP_and_1611_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100101"));
        COMP_LOOP_COMP_LOOP_and_1612_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100110"));
        COMP_LOOP_COMP_LOOP_and_1613_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100111"));
        COMP_LOOP_COMP_LOOP_and_1615_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101001"));
        COMP_LOOP_COMP_LOOP_and_1616_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101010"));
        COMP_LOOP_COMP_LOOP_and_1617_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101011"));
        COMP_LOOP_COMP_LOOP_and_1618_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101100"));
        COMP_LOOP_COMP_LOOP_and_1619_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101101"));
        COMP_LOOP_COMP_LOOP_and_1620_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101110"));
        COMP_LOOP_COMP_LOOP_and_1621_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101111"));
        COMP_LOOP_COMP_LOOP_and_1623_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110001"));
        COMP_LOOP_COMP_LOOP_and_1624_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110010"));
        COMP_LOOP_COMP_LOOP_and_1625_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110011"));
        COMP_LOOP_COMP_LOOP_and_1626_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110100"));
        COMP_LOOP_COMP_LOOP_and_1627_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110101"));
        COMP_LOOP_COMP_LOOP_and_1628_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110110"));
        COMP_LOOP_COMP_LOOP_and_1629_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110111"));
        COMP_LOOP_COMP_LOOP_and_1630_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111000"));
        COMP_LOOP_COMP_LOOP_and_1631_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111001"));
        COMP_LOOP_COMP_LOOP_and_1632_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111010"));
        COMP_LOOP_COMP_LOOP_and_1633_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111011"));
        COMP_LOOP_COMP_LOOP_and_1634_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111100"));
        COMP_LOOP_COMP_LOOP_and_1635_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
        COMP_LOOP_COMP_LOOP_and_1636_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111110"));
        COMP_LOOP_COMP_LOOP_and_1637_itm <= CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1435_itm <= '0';
      ELSIF ( and_dcpl_390 = '0' ) THEN
        COMP_LOOP_nor_1435_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1446_itm <= '0';
      ELSIF ( (NOT(mux_3188_nl AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_nor_1446_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1439_itm <= '0';
      ELSIF ( and_dcpl_410 = '0' ) THEN
        COMP_LOOP_nor_1439_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1420_itm <= '0';
      ELSIF ( and_dcpl_410 = '0' ) THEN
        COMP_LOOP_nor_1420_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1432_itm <= '0';
      ELSIF ( (NOT(mux_3192_nl AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_nor_1432_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(4
            DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1424_itm <= '0';
      ELSIF ( and_dcpl_407 = '0' ) THEN
        COMP_LOOP_nor_1424_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1410_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_1410_itm <= NOT((COMP_LOOP_7_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_7_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_7_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1403_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_1403_itm <= NOT(CONV_SL_1_1(COMP_LOOP_7_acc_10_itm_10_1_1(5
            DOWNTO 2)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_811, mux_3193_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_10_0_sva_9_0)
            + UNSIGNED(COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'( "111")), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(not_tmp_811, and_705_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_sva <= COMP_LOOP_8_acc_10_itm_10_1_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(not_tmp_811, mux_3197_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm <= COMP_LOOP_1_acc_nl(10);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_29_itm <= '0';
        COMP_LOOP_nor_1625_itm <= '0';
        COMP_LOOP_nor_1626_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1829_itm <= '0';
        COMP_LOOP_nor_1628_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1833_itm <= '0';
        COMP_LOOP_nor_1632_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1836_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1837_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1838_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1839_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1840_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1841_itm <= '0';
        COMP_LOOP_nor_1640_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1843_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1845_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1846_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1847_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1848_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1849_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1851_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1852_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1853_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1854_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1855_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1856_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1857_itm <= '0';
        COMP_LOOP_nor_1655_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1859_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1860_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1861_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1863_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1864_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1865_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1867_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1868_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1869_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1870_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1871_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1872_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1873_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1875_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1876_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1877_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1878_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1879_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1880_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1881_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1882_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1883_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1884_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1885_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1886_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1887_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1888_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1889_itm <= '0';
      ELSIF ( mux_3201_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_29_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
        COMP_LOOP_nor_1625_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_nor_1626_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1829_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000011"));
        COMP_LOOP_nor_1628_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1833_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("000111"));
        COMP_LOOP_nor_1632_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1836_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001010"));
        COMP_LOOP_COMP_LOOP_and_1837_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001011"));
        COMP_LOOP_COMP_LOOP_and_1838_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001100"));
        COMP_LOOP_COMP_LOOP_and_1839_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001101"));
        COMP_LOOP_COMP_LOOP_and_1840_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001110"));
        COMP_LOOP_COMP_LOOP_and_1841_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("001111"));
        COMP_LOOP_nor_1640_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(1))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
        COMP_LOOP_COMP_LOOP_and_1843_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010001"));
        COMP_LOOP_COMP_LOOP_and_1845_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010011"));
        COMP_LOOP_COMP_LOOP_and_1846_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010100"));
        COMP_LOOP_COMP_LOOP_and_1847_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010101"));
        COMP_LOOP_COMP_LOOP_and_1848_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010110"));
        COMP_LOOP_COMP_LOOP_and_1849_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("010111"));
        COMP_LOOP_COMP_LOOP_and_1851_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011001"));
        COMP_LOOP_COMP_LOOP_and_1852_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011010"));
        COMP_LOOP_COMP_LOOP_and_1853_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011011"));
        COMP_LOOP_COMP_LOOP_and_1854_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011100"));
        COMP_LOOP_COMP_LOOP_and_1855_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011101"));
        COMP_LOOP_COMP_LOOP_and_1856_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011110"));
        COMP_LOOP_COMP_LOOP_and_1857_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("011111"));
        COMP_LOOP_nor_1655_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(4
            DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
        COMP_LOOP_COMP_LOOP_and_1859_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100001"));
        COMP_LOOP_COMP_LOOP_and_1860_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100010"));
        COMP_LOOP_COMP_LOOP_and_1861_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100011"));
        COMP_LOOP_COMP_LOOP_and_1863_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100101"));
        COMP_LOOP_COMP_LOOP_and_1864_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100110"));
        COMP_LOOP_COMP_LOOP_and_1865_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("100111"));
        COMP_LOOP_COMP_LOOP_and_1867_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101001"));
        COMP_LOOP_COMP_LOOP_and_1868_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101010"));
        COMP_LOOP_COMP_LOOP_and_1869_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101011"));
        COMP_LOOP_COMP_LOOP_and_1870_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101100"));
        COMP_LOOP_COMP_LOOP_and_1871_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101101"));
        COMP_LOOP_COMP_LOOP_and_1872_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101110"));
        COMP_LOOP_COMP_LOOP_and_1873_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("101111"));
        COMP_LOOP_COMP_LOOP_and_1875_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110001"));
        COMP_LOOP_COMP_LOOP_and_1876_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110010"));
        COMP_LOOP_COMP_LOOP_and_1877_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110011"));
        COMP_LOOP_COMP_LOOP_and_1878_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110100"));
        COMP_LOOP_COMP_LOOP_and_1879_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110101"));
        COMP_LOOP_COMP_LOOP_and_1880_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110110"));
        COMP_LOOP_COMP_LOOP_and_1881_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("110111"));
        COMP_LOOP_COMP_LOOP_and_1882_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111000"));
        COMP_LOOP_COMP_LOOP_and_1883_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111001"));
        COMP_LOOP_COMP_LOOP_and_1884_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111010"));
        COMP_LOOP_COMP_LOOP_and_1885_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111011"));
        COMP_LOOP_COMP_LOOP_and_1886_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111100"));
        COMP_LOOP_COMP_LOOP_and_1887_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
        COMP_LOOP_COMP_LOOP_and_1888_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111110"));
        COMP_LOOP_COMP_LOOP_and_1889_itm <= CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(5
            DOWNTO 0)=STD_LOGIC_VECTOR'("111111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1663_itm <= '0';
      ELSIF ( (mux_3205_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_nor_1663_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1659_itm <= '0';
      ELSIF ( (mux_3210_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_nor_1659_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(4)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1633_itm <= '0';
      ELSIF ( (mux_3216_nl OR (fsm_output(7))) = '1' ) THEN
        COMP_LOOP_nor_1633_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1642_itm <= '0';
      ELSIF ( and_dcpl_410 = '0' ) THEN
        COMP_LOOP_nor_1642_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(3))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1648_itm <= '0';
      ELSIF ( and_dcpl_404 = '0' ) THEN
        COMP_LOOP_nor_1648_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(2))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(1)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1630_itm <= '0';
      ELSIF ( (NOT(mux_3219_nl AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_nor_1630_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(0)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1670_itm <= '0';
      ELSIF ( and_dcpl_411 = '0' ) THEN
        COMP_LOOP_nor_1670_itm <= NOT(CONV_SL_1_1(COMP_LOOP_8_acc_10_itm_10_1_1(3
            DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_nor_1629_itm <= '0';
      ELSIF ( or_dcpl_125 = '0' ) THEN
        COMP_LOOP_nor_1629_itm <= NOT((COMP_LOOP_8_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(4))
            OR (COMP_LOOP_8_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_8_acc_10_itm_10_1_1(1)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1104_itm <= '0';
      ELSIF ( (NOT(mux_3223_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1104_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_111_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_24_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_23_cse, COMP_LOOP_COMP_LOOP_and_1104_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_387));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1106_itm <= '0';
      ELSIF ( (NOT(mux_3226_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1106_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_112_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_25_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_24_cse, COMP_LOOP_COMP_LOOP_and_1106_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_388));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1110_itm <= '0';
      ELSIF ( (NOT(mux_3227_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1110_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_113_nl,
            COMP_LOOP_COMP_LOOP_and_1110_nl, and_dcpl_261);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1118_itm <= '0';
      ELSIF ( (NOT(mux_3229_nl AND (NOT (fsm_output(7))))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1118_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_114_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_87_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_25_cse, COMP_LOOP_COMP_LOOP_and_1118_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_421));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1370_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3231_nl, (fsm_output(7)), fsm_output(5))) = '1' )
          THEN
        COMP_LOOP_COMP_LOOP_and_1370_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_65_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_98_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse, COMP_LOOP_COMP_LOOP_and_1370_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_421));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1577_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1584_itm <= '0';
      ELSIF ( COMP_LOOP_or_151_cse = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1577_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_67_nl,
            COMP_LOOP_COMP_LOOP_and_1577_nl, and_dcpl_258);
        COMP_LOOP_COMP_LOOP_and_1584_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_68_nl,
            COMP_LOOP_COMP_LOOP_and_1584_nl, and_dcpl_258);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1594_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_1614_itm <= '0';
      ELSIF ( COMP_LOOP_or_153_cse = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1594_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_317_nl,
            COMP_LOOP_COMP_LOOP_and_1594_nl, and_dcpl_90);
        COMP_LOOP_COMP_LOOP_and_1614_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_324_nl,
            COMP_LOOP_COMP_LOOP_and_1614_nl, and_dcpl_90);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1598_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3243_nl, (fsm_output(7)), fsm_output(6))) = '1' )
          THEN
        COMP_LOOP_COMP_LOOP_and_1598_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_319_nl,
            COMP_LOOP_COMP_LOOP_and_1598_nl, and_dcpl_370);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1607_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_tmp_3102, mux_3246_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1607_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_320_nl,
            COMP_LOOP_COMP_LOOP_and_1607_nl, and_458_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1610_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3253_nl, mux_3249_nl, fsm_output(6))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1610_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_321_nl,
            COMP_LOOP_COMP_LOOP_and_1610_nl, and_dcpl_118);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1622_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_tmp_3102, mux_3256_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1622_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_325_nl,
            COMP_LOOP_COMP_LOOP_and_1622_nl, and_459_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1831_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3264_nl, and_705_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1831_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_69_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_99_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_cse, COMP_LOOP_COMP_LOOP_and_1831_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_112));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1832_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3274_nl, mux_3267_nl, fsm_output(3))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1832_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_326_nl,
            COMP_LOOP_COMP_LOOP_and_1832_nl, and_461_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1835_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3283_nl, mux_297_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1835_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_327_nl,
            COMP_LOOP_COMP_LOOP_and_1835_nl, and_463_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1844_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_tmp_3133, mux_3286_nl, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1844_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_328_nl,
            COMP_LOOP_COMP_LOOP_and_1844_nl, and_dcpl_90);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1850_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_tmp_3133, mux_tmp_3218, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1850_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_329_nl,
            COMP_LOOP_COMP_LOOP_and_1850_nl, and_dcpl_382);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1862_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3292_nl, mux_297_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1862_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_331_nl,
            COMP_LOOP_COMP_LOOP_and_1862_nl, and_465_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1866_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3298_nl, mux_297_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1866_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_332_nl,
            COMP_LOOP_COMP_LOOP_and_1866_nl, and_468_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_1874_itm <= '0';
      ELSIF ( (MUX_s_1_2_2(mux_3302_nl, and_705_cse, fsm_output(5))) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_1874_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_71_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse, COMP_LOOP_COMP_LOOP_and_1874_nl,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt
            & and_dcpl_86));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_583_itm <= '0';
      ELSIF ( (NOT(mux_3306_nl AND nor_399_cse)) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_583_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_72_nl,
            COMP_LOOP_COMP_LOOP_and_583_nl, and_dcpl_258);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse, STD_LOGIC_VECTOR'( and_dcpl_74
            & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_244_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, STD_LOGIC_VECTOR'( and_dcpl_74
            & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_74_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse, STD_LOGIC_VECTOR'( and_dcpl_74
            & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_75_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse, STD_LOGIC_VECTOR'( and_dcpl_74
            & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_nor_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_76_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse, STD_LOGIC_VECTOR'( and_dcpl_74
            & and_dcpl_77 & and_dcpl_258 & COMP_LOOP_or_120_rgt));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm <= '0';
        COMP_LOOP_tmp_nor_10_itm <= '0';
        COMP_LOOP_tmp_nor_151_itm <= '0';
        COMP_LOOP_tmp_nor_153_itm <= '0';
        COMP_LOOP_tmp_nor_157_itm <= '0';
        COMP_LOOP_tmp_nor_165_itm <= '0';
        COMP_LOOP_tmp_nor_180_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_5_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_76_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_77_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_79_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_80_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_81_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_82_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_83_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_84_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_85_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_49_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_86_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_50_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_49_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_87_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_50_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_88_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_52_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_89_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_52_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_90_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_91_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_92_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_56_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_93_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_57_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_56_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_95_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_58_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_57_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_96_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_59_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_58_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_97_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_60_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_59_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_98_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_61_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_60_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_99_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_62_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_61_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_nor_1_nl,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_63_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_62_cse,
            STD_LOGIC_VECTOR'( and_dcpl_74 & and_dcpl_77 & COMP_LOOP_or_120_rgt));
        COMP_LOOP_tmp_nor_10_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_57_nl, COMP_LOOP_tmp_nor_10_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse, COMP_LOOP_tmp_nor_150_cse, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_77 & and_dcpl_259 & COMP_LOOP_or_74_cse));
        COMP_LOOP_tmp_nor_151_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_58_nl, COMP_LOOP_tmp_nor_18_cse,
            COMP_LOOP_tmp_nor_150_cse, COMP_LOOP_tmp_nor_151_cse, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_77 & and_dcpl_259 & COMP_LOOP_or_74_cse));
        COMP_LOOP_tmp_nor_153_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_60_nl, COMP_LOOP_tmp_nor_150_cse,
            COMP_LOOP_tmp_nor_151_cse, COMP_LOOP_tmp_nor_153_cse, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_77 & and_dcpl_259 & COMP_LOOP_or_74_cse));
        COMP_LOOP_tmp_nor_157_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_64_nl, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse,
            COMP_LOOP_tmp_nor_153_cse, COMP_LOOP_tmp_nor_10_cse, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_77 & and_dcpl_259 & COMP_LOOP_or_74_cse));
        COMP_LOOP_tmp_nor_165_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_72_nl, COMP_LOOP_tmp_nor_151_cse,
            COMP_LOOP_tmp_nor_10_cse, COMP_LOOP_tmp_nor_18_cse, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_77 & and_dcpl_259 & COMP_LOOP_or_74_cse));
        COMP_LOOP_tmp_nor_180_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_87_nl, COMP_LOOP_tmp_nor_153_cse,
            COMP_LOOP_tmp_nor_18_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse, STD_LOGIC_VECTOR'(
            and_dcpl_74 & and_dcpl_77 & and_dcpl_259 & COMP_LOOP_or_74_cse));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_2_tmp_mul_idiv_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (and_dcpl_77 OR and_dcpl_259 OR and_dcpl_260) = '1' ) THEN
        COMP_LOOP_2_tmp_mul_idiv_sva <= z_out_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(or_dcpl_134 OR or_dcpl_122)) = '1' ) THEN
        COMP_LOOP_tmp_mux1h_itm <= MUX1HOT_v_64_8_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_8_i_q_d,
            twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_32_i_q_d,
            twiddle_rsc_0_40_i_q_d, twiddle_rsc_0_48_i_q_d, twiddle_rsc_0_56_i_q_d,
            STD_LOGIC_VECTOR'( COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_2_tmp_lshift_ncse_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (and_dcpl_77 OR and_dcpl_263) = '1' ) THEN
        COMP_LOOP_2_tmp_lshift_ncse_sva <= MUX_v_10_2_2(z_out_1, z_out_7, and_dcpl_263);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_77 OR and_dcpl_258 OR and_dcpl_432 OR and_dcpl_263 OR COMP_LOOP_1_acc_8_itm_mx0c4
          OR and_dcpl_86 OR and_dcpl_343 OR and_dcpl_90 OR and_dcpl_346 OR and_dcpl_95
          OR and_dcpl_349 OR and_dcpl_99 OR and_dcpl_351 OR and_dcpl_104 OR and_dcpl_354
          OR and_dcpl_106 OR and_dcpl_357 OR and_dcpl_109 OR and_dcpl_359) = '1'
          ) THEN
        COMP_LOOP_1_acc_8_itm <= MUX1HOT_v_64_68_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
            vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
            vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
            vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
            vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, vec_rsc_0_16_i_q_d, vec_rsc_0_17_i_q_d,
            vec_rsc_0_18_i_q_d, vec_rsc_0_19_i_q_d, vec_rsc_0_20_i_q_d, vec_rsc_0_21_i_q_d,
            vec_rsc_0_22_i_q_d, vec_rsc_0_23_i_q_d, vec_rsc_0_24_i_q_d, vec_rsc_0_25_i_q_d,
            vec_rsc_0_26_i_q_d, vec_rsc_0_27_i_q_d, vec_rsc_0_28_i_q_d, vec_rsc_0_29_i_q_d,
            vec_rsc_0_30_i_q_d, vec_rsc_0_31_i_q_d, vec_rsc_0_32_i_q_d, vec_rsc_0_33_i_q_d,
            vec_rsc_0_34_i_q_d, vec_rsc_0_35_i_q_d, vec_rsc_0_36_i_q_d, vec_rsc_0_37_i_q_d,
            vec_rsc_0_38_i_q_d, vec_rsc_0_39_i_q_d, vec_rsc_0_40_i_q_d, vec_rsc_0_41_i_q_d,
            vec_rsc_0_42_i_q_d, vec_rsc_0_43_i_q_d, vec_rsc_0_44_i_q_d, vec_rsc_0_45_i_q_d,
            vec_rsc_0_46_i_q_d, vec_rsc_0_47_i_q_d, vec_rsc_0_48_i_q_d, vec_rsc_0_49_i_q_d,
            vec_rsc_0_50_i_q_d, vec_rsc_0_51_i_q_d, vec_rsc_0_52_i_q_d, vec_rsc_0_53_i_q_d,
            vec_rsc_0_54_i_q_d, vec_rsc_0_55_i_q_d, vec_rsc_0_56_i_q_d, vec_rsc_0_57_i_q_d,
            vec_rsc_0_58_i_q_d, vec_rsc_0_59_i_q_d, vec_rsc_0_60_i_q_d, vec_rsc_0_61_i_q_d,
            vec_rsc_0_62_i_q_d, vec_rsc_0_63_i_q_d, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_acc_17_nl),
            64)), twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_26_i_q_d, COMP_LOOP_1_modulo_dev_cmp_return_rsc_z,
            STD_LOGIC_VECTOR'( COMP_LOOP_or_nl & COMP_LOOP_or_1_nl & COMP_LOOP_or_2_nl
            & COMP_LOOP_or_3_nl & COMP_LOOP_or_4_nl & COMP_LOOP_or_5_nl & COMP_LOOP_or_6_nl
            & COMP_LOOP_or_7_nl & COMP_LOOP_or_8_nl & COMP_LOOP_or_9_nl & COMP_LOOP_or_10_nl
            & COMP_LOOP_or_11_nl & COMP_LOOP_or_12_nl & COMP_LOOP_or_13_nl & COMP_LOOP_or_14_nl
            & COMP_LOOP_or_15_nl & COMP_LOOP_or_16_nl & COMP_LOOP_or_17_nl & COMP_LOOP_or_18_nl
            & COMP_LOOP_or_19_nl & COMP_LOOP_or_20_nl & COMP_LOOP_or_21_nl & COMP_LOOP_or_22_nl
            & COMP_LOOP_or_23_nl & COMP_LOOP_or_24_nl & COMP_LOOP_or_25_nl & COMP_LOOP_or_26_nl
            & COMP_LOOP_or_27_nl & COMP_LOOP_or_28_nl & COMP_LOOP_or_29_nl & COMP_LOOP_or_30_nl
            & COMP_LOOP_or_31_nl & COMP_LOOP_or_32_nl & COMP_LOOP_or_33_nl & COMP_LOOP_or_34_nl
            & COMP_LOOP_or_35_nl & COMP_LOOP_or_36_nl & COMP_LOOP_or_37_nl & COMP_LOOP_or_38_nl
            & COMP_LOOP_or_39_nl & COMP_LOOP_or_40_nl & COMP_LOOP_or_41_nl & COMP_LOOP_or_42_nl
            & COMP_LOOP_or_43_nl & COMP_LOOP_or_44_nl & COMP_LOOP_or_45_nl & COMP_LOOP_or_46_nl
            & COMP_LOOP_or_47_nl & COMP_LOOP_or_48_nl & COMP_LOOP_or_49_nl & COMP_LOOP_or_50_nl
            & COMP_LOOP_or_51_nl & COMP_LOOP_or_52_nl & COMP_LOOP_or_53_nl & COMP_LOOP_or_54_nl
            & COMP_LOOP_or_55_nl & COMP_LOOP_or_56_nl & COMP_LOOP_or_57_nl & COMP_LOOP_or_58_nl
            & COMP_LOOP_or_59_nl & COMP_LOOP_or_60_nl & COMP_LOOP_or_61_nl & COMP_LOOP_or_62_nl
            & COMP_LOOP_or_63_nl & COMP_LOOP_or_68_itm & and_dcpl_432 & and_dcpl_263
            & COMP_LOOP_1_acc_8_itm_mx0c4));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm <= '0';
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_36_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_64_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_63_cse, COMP_LOOP_or_120_rgt);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_65_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_64_cse, COMP_LOOP_or_120_rgt);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_66_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_65_cse, COMP_LOOP_or_120_rgt);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_67_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_66_cse, COMP_LOOP_or_120_rgt);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_68_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_67_cse, COMP_LOOP_or_120_rgt);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_69_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_68_cse, COMP_LOOP_or_120_rgt);
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse,
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_69_cse, COMP_LOOP_or_120_rgt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_3_tmp_lshift_ncse_sva <= STD_LOGIC_VECTOR'( "000000000");
        COMP_LOOP_tmp_nor_206_itm <= '0';
        COMP_LOOP_tmp_nor_207_itm <= '0';
        COMP_LOOP_tmp_nor_209_itm <= '0';
        COMP_LOOP_tmp_nor_213_itm <= '0';
        COMP_LOOP_tmp_nor_220_itm <= '0';
      ELSIF ( COMP_LOOP_tmp_or_43_cse = '1' ) THEN
        COMP_LOOP_3_tmp_lshift_ncse_sva <= MUX_v_9_2_2((z_out_1(8 DOWNTO 0)), (z_out_7(8
            DOWNTO 0)), and_dcpl_261);
        COMP_LOOP_tmp_nor_206_itm <= COMP_LOOP_tmp_nor_34_cse;
        COMP_LOOP_tmp_nor_207_itm <= COMP_LOOP_tmp_nor_35_cse;
        COMP_LOOP_tmp_nor_209_itm <= COMP_LOOP_tmp_nor_37_cse;
        COMP_LOOP_tmp_nor_213_itm <= COMP_LOOP_tmp_nor_41_cse;
        COMP_LOOP_tmp_nor_220_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_474_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_1_itm <= MUX1HOT_v_64_64_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
            twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d,
            twiddle_rsc_0_5_i_q_d, twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d,
            twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_9_i_q_d, twiddle_rsc_0_10_i_q_d,
            twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_13_i_q_d,
            twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_16_i_q_d,
            twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_19_i_q_d,
            twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_21_i_q_d, twiddle_rsc_0_22_i_q_d,
            twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_25_i_q_d,
            twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_27_i_q_d, twiddle_rsc_0_28_i_q_d,
            twiddle_rsc_0_29_i_q_d, twiddle_rsc_0_30_i_q_d, twiddle_rsc_0_31_i_q_d,
            twiddle_rsc_0_32_i_q_d, twiddle_rsc_0_33_i_q_d, twiddle_rsc_0_34_i_q_d,
            twiddle_rsc_0_35_i_q_d, twiddle_rsc_0_36_i_q_d, twiddle_rsc_0_37_i_q_d,
            twiddle_rsc_0_38_i_q_d, twiddle_rsc_0_39_i_q_d, twiddle_rsc_0_40_i_q_d,
            twiddle_rsc_0_41_i_q_d, twiddle_rsc_0_42_i_q_d, twiddle_rsc_0_43_i_q_d,
            twiddle_rsc_0_44_i_q_d, twiddle_rsc_0_45_i_q_d, twiddle_rsc_0_46_i_q_d,
            twiddle_rsc_0_47_i_q_d, twiddle_rsc_0_48_i_q_d, twiddle_rsc_0_49_i_q_d,
            twiddle_rsc_0_50_i_q_d, twiddle_rsc_0_51_i_q_d, twiddle_rsc_0_52_i_q_d,
            twiddle_rsc_0_53_i_q_d, twiddle_rsc_0_54_i_q_d, twiddle_rsc_0_55_i_q_d,
            twiddle_rsc_0_56_i_q_d, twiddle_rsc_0_57_i_q_d, twiddle_rsc_0_58_i_q_d,
            twiddle_rsc_0_59_i_q_d, twiddle_rsc_0_60_i_q_d, twiddle_rsc_0_61_i_q_d,
            twiddle_rsc_0_62_i_q_d, twiddle_rsc_0_63_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_249_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_nl
            & COMP_LOOP_tmp_and_250_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_nl &
            COMP_LOOP_tmp_and_251_nl & COMP_LOOP_tmp_and_252_nl & COMP_LOOP_tmp_and_253_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_nl & COMP_LOOP_tmp_and_254_nl &
            COMP_LOOP_tmp_and_255_nl & COMP_LOOP_tmp_and_256_nl & COMP_LOOP_tmp_and_257_nl
            & COMP_LOOP_tmp_and_258_nl & COMP_LOOP_tmp_and_259_nl & COMP_LOOP_tmp_and_260_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_22_nl & COMP_LOOP_tmp_and_261_nl &
            COMP_LOOP_tmp_and_262_nl & COMP_LOOP_tmp_and_263_nl & COMP_LOOP_tmp_and_264_nl
            & COMP_LOOP_tmp_and_265_nl & COMP_LOOP_tmp_and_266_nl & COMP_LOOP_tmp_and_267_nl
            & COMP_LOOP_tmp_and_268_nl & COMP_LOOP_tmp_and_269_nl & COMP_LOOP_tmp_and_270_nl
            & COMP_LOOP_tmp_and_271_nl & COMP_LOOP_tmp_and_272_nl & COMP_LOOP_tmp_and_273_nl
            & COMP_LOOP_tmp_and_274_nl & COMP_LOOP_tmp_and_275_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_nl
            & COMP_LOOP_tmp_and_276_nl & COMP_LOOP_tmp_and_277_nl & COMP_LOOP_tmp_and_278_nl
            & COMP_LOOP_tmp_and_279_nl & COMP_LOOP_tmp_and_280_nl & COMP_LOOP_tmp_and_281_nl
            & COMP_LOOP_tmp_and_282_nl & COMP_LOOP_tmp_and_283_nl & COMP_LOOP_tmp_and_284_nl
            & COMP_LOOP_tmp_and_285_nl & COMP_LOOP_tmp_and_286_nl & COMP_LOOP_tmp_and_287_nl
            & COMP_LOOP_tmp_and_288_nl & COMP_LOOP_tmp_and_289_nl & COMP_LOOP_tmp_and_290_nl
            & COMP_LOOP_tmp_and_291_nl & COMP_LOOP_tmp_and_292_nl & COMP_LOOP_tmp_and_293_nl
            & COMP_LOOP_tmp_and_294_nl & COMP_LOOP_tmp_and_295_nl & COMP_LOOP_tmp_and_296_nl
            & COMP_LOOP_tmp_and_297_nl & COMP_LOOP_tmp_and_298_nl & COMP_LOOP_tmp_and_299_nl
            & COMP_LOOP_tmp_and_300_nl & COMP_LOOP_tmp_and_301_nl & COMP_LOOP_tmp_and_302_nl
            & COMP_LOOP_tmp_and_303_nl & COMP_LOOP_tmp_and_304_nl & COMP_LOOP_tmp_and_305_nl
            & COMP_LOOP_tmp_and_306_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( nor_1579_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_2_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_2_i_q_d,
            twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_8_i_q_d,
            twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_14_i_q_d,
            twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_20_i_q_d,
            twiddle_rsc_0_22_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_26_i_q_d,
            twiddle_rsc_0_28_i_q_d, twiddle_rsc_0_30_i_q_d, twiddle_rsc_0_32_i_q_d,
            twiddle_rsc_0_34_i_q_d, twiddle_rsc_0_36_i_q_d, twiddle_rsc_0_38_i_q_d,
            twiddle_rsc_0_40_i_q_d, twiddle_rsc_0_42_i_q_d, twiddle_rsc_0_44_i_q_d,
            twiddle_rsc_0_46_i_q_d, twiddle_rsc_0_48_i_q_d, twiddle_rsc_0_50_i_q_d,
            twiddle_rsc_0_52_i_q_d, twiddle_rsc_0_54_i_q_d, twiddle_rsc_0_56_i_q_d,
            twiddle_rsc_0_58_i_q_d, twiddle_rsc_0_60_i_q_d, twiddle_rsc_0_62_i_q_d,
            STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_222_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_70_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_71_nl & COMP_LOOP_tmp_and_223_nl &
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_73_nl & COMP_LOOP_tmp_and_224_nl & COMP_LOOP_tmp_and_225_nl
            & COMP_LOOP_tmp_and_226_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_77_nl &
            COMP_LOOP_tmp_and_227_nl & COMP_LOOP_tmp_and_228_nl & COMP_LOOP_tmp_and_229_nl
            & COMP_LOOP_tmp_and_230_nl & COMP_LOOP_tmp_and_231_nl & COMP_LOOP_tmp_and_232_nl
            & COMP_LOOP_tmp_and_233_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_nl &
            COMP_LOOP_tmp_and_234_nl & COMP_LOOP_tmp_and_235_nl & COMP_LOOP_tmp_and_236_nl
            & COMP_LOOP_tmp_and_237_nl & COMP_LOOP_tmp_and_238_nl & COMP_LOOP_tmp_and_239_nl
            & COMP_LOOP_tmp_and_240_nl & COMP_LOOP_tmp_and_241_nl & COMP_LOOP_tmp_and_242_nl
            & COMP_LOOP_tmp_and_243_nl & COMP_LOOP_tmp_and_244_nl & COMP_LOOP_tmp_and_245_nl
            & COMP_LOOP_tmp_and_246_nl & COMP_LOOP_tmp_and_247_nl & COMP_LOOP_tmp_and_248_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_476_tmp = '0' ) THEN
        COMP_LOOP_tmp_mux1h_3_itm <= MUX1HOT_v_64_64_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
            twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d,
            twiddle_rsc_0_5_i_q_d, twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d,
            twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_9_i_q_d, twiddle_rsc_0_10_i_q_d,
            twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_13_i_q_d,
            twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_16_i_q_d,
            twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_19_i_q_d,
            twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_21_i_q_d, twiddle_rsc_0_22_i_q_d,
            twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_25_i_q_d,
            twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_27_i_q_d, twiddle_rsc_0_28_i_q_d,
            twiddle_rsc_0_29_i_q_d, twiddle_rsc_0_30_i_q_d, twiddle_rsc_0_31_i_q_d,
            twiddle_rsc_0_32_i_q_d, twiddle_rsc_0_33_i_q_d, twiddle_rsc_0_34_i_q_d,
            twiddle_rsc_0_35_i_q_d, twiddle_rsc_0_36_i_q_d, twiddle_rsc_0_37_i_q_d,
            twiddle_rsc_0_38_i_q_d, twiddle_rsc_0_39_i_q_d, twiddle_rsc_0_40_i_q_d,
            twiddle_rsc_0_41_i_q_d, twiddle_rsc_0_42_i_q_d, twiddle_rsc_0_43_i_q_d,
            twiddle_rsc_0_44_i_q_d, twiddle_rsc_0_45_i_q_d, twiddle_rsc_0_46_i_q_d,
            twiddle_rsc_0_47_i_q_d, twiddle_rsc_0_48_i_q_d, twiddle_rsc_0_49_i_q_d,
            twiddle_rsc_0_50_i_q_d, twiddle_rsc_0_51_i_q_d, twiddle_rsc_0_52_i_q_d,
            twiddle_rsc_0_53_i_q_d, twiddle_rsc_0_54_i_q_d, twiddle_rsc_0_55_i_q_d,
            twiddle_rsc_0_56_i_q_d, twiddle_rsc_0_57_i_q_d, twiddle_rsc_0_58_i_q_d,
            twiddle_rsc_0_59_i_q_d, twiddle_rsc_0_60_i_q_d, twiddle_rsc_0_61_i_q_d,
            twiddle_rsc_0_62_i_q_d, twiddle_rsc_0_63_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_164_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_102_nl
            & COMP_LOOP_tmp_and_165_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_nl &
            COMP_LOOP_tmp_and_166_nl & COMP_LOOP_tmp_and_167_nl & COMP_LOOP_tmp_and_168_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_nl & COMP_LOOP_tmp_and_169_nl &
            COMP_LOOP_tmp_and_170_nl & COMP_LOOP_tmp_and_171_nl & COMP_LOOP_tmp_and_172_nl
            & COMP_LOOP_tmp_and_173_nl & COMP_LOOP_tmp_and_174_nl & COMP_LOOP_tmp_and_175_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_nl & COMP_LOOP_tmp_and_176_nl &
            COMP_LOOP_tmp_and_177_nl & COMP_LOOP_tmp_and_178_nl & COMP_LOOP_tmp_and_179_nl
            & COMP_LOOP_tmp_and_180_nl & COMP_LOOP_tmp_and_181_nl & COMP_LOOP_tmp_and_182_nl
            & COMP_LOOP_tmp_and_183_nl & COMP_LOOP_tmp_and_184_nl & COMP_LOOP_tmp_and_185_nl
            & COMP_LOOP_tmp_and_186_nl & COMP_LOOP_tmp_and_187_nl & COMP_LOOP_tmp_and_188_nl
            & COMP_LOOP_tmp_and_189_nl & COMP_LOOP_tmp_and_190_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_nl
            & COMP_LOOP_tmp_and_191_nl & COMP_LOOP_tmp_and_192_nl & COMP_LOOP_tmp_and_193_nl
            & COMP_LOOP_tmp_and_194_nl & COMP_LOOP_tmp_and_195_nl & COMP_LOOP_tmp_and_196_nl
            & COMP_LOOP_tmp_and_197_nl & COMP_LOOP_tmp_and_198_nl & COMP_LOOP_tmp_and_199_nl
            & COMP_LOOP_tmp_and_200_nl & COMP_LOOP_tmp_and_201_nl & COMP_LOOP_tmp_and_202_nl
            & COMP_LOOP_tmp_and_203_nl & COMP_LOOP_tmp_and_204_nl & COMP_LOOP_tmp_and_205_nl
            & COMP_LOOP_tmp_and_206_nl & COMP_LOOP_tmp_and_207_nl & COMP_LOOP_tmp_and_208_nl
            & COMP_LOOP_tmp_and_209_nl & COMP_LOOP_tmp_and_210_nl & COMP_LOOP_tmp_and_211_nl
            & COMP_LOOP_tmp_and_212_nl & COMP_LOOP_tmp_and_213_nl & COMP_LOOP_tmp_and_214_nl
            & COMP_LOOP_tmp_and_215_nl & COMP_LOOP_tmp_and_216_nl & COMP_LOOP_tmp_and_217_nl
            & COMP_LOOP_tmp_and_218_nl & COMP_LOOP_tmp_and_219_nl & COMP_LOOP_tmp_and_220_nl
            & COMP_LOOP_tmp_and_221_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm <= '0';
      ELSIF ( COMP_LOOP_or_74_cse = '1' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( nor_tmp_396 = '0' ) THEN
        COMP_LOOP_tmp_mux1h_4_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_4_i_q_d,
            twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_16_i_q_d,
            twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_28_i_q_d,
            twiddle_rsc_0_32_i_q_d, twiddle_rsc_0_36_i_q_d, twiddle_rsc_0_40_i_q_d,
            twiddle_rsc_0_44_i_q_d, twiddle_rsc_0_48_i_q_d, twiddle_rsc_0_52_i_q_d,
            twiddle_rsc_0_56_i_q_d, twiddle_rsc_0_60_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_152_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_164_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_165_nl
            & COMP_LOOP_tmp_and_153_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_167_nl &
            COMP_LOOP_tmp_and_154_nl & COMP_LOOP_tmp_and_155_nl & COMP_LOOP_tmp_and_156_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_171_nl & COMP_LOOP_tmp_and_157_nl &
            COMP_LOOP_tmp_and_158_nl & COMP_LOOP_tmp_and_159_nl & COMP_LOOP_tmp_and_160_nl
            & COMP_LOOP_tmp_and_161_nl & COMP_LOOP_tmp_and_162_nl & COMP_LOOP_tmp_and_163_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (((NOT((COMP_LOOP_2_tmp_lshift_ncse_sva(0)) AND COMP_LOOP_tmp_nor_10_itm))
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_274_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_276_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_280_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm OR COMP_LOOP_COMP_LOOP_and_102_itm
          OR COMP_LOOP_COMP_LOOP_and_106_itm OR COMP_LOOP_COMP_LOOP_and_107_itm OR
          COMP_LOOP_COMP_LOOP_and_108_itm OR COMP_LOOP_COMP_LOOP_and_109_itm OR COMP_LOOP_COMP_LOOP_and_110_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_288_rgt OR COMP_LOOP_COMP_LOOP_and_1104_itm
          OR COMP_LOOP_COMP_LOOP_and_1106_itm OR COMP_LOOP_COMP_LOOP_and_1118_itm
          OR COMP_LOOP_COMP_LOOP_and_115_itm OR COMP_LOOP_COMP_LOOP_and_116_itm OR
          COMP_LOOP_COMP_LOOP_and_117_itm OR COMP_LOOP_COMP_LOOP_and_118_itm OR COMP_LOOP_COMP_LOOP_and_120_itm
          OR COMP_LOOP_COMP_LOOP_and_121_itm OR COMP_LOOP_COMP_LOOP_and_122_itm OR
          COMP_LOOP_COMP_LOOP_and_123_itm OR COMP_LOOP_COMP_LOOP_and_124_itm OR COMP_LOOP_COMP_LOOP_and_125_itm
          OR COMP_LOOP_COMP_LOOP_and_1370_itm OR COMP_LOOP_COMP_LOOP_and_1831_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_304_rgt OR COMP_LOOP_COMP_LOOP_and_1874_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm
          OR and_dcpl_432 OR and_dcpl_263) AND mux_3353_nl) = '1' ) THEN
        tmp_21_sva_1 <= MUX1HOT_v_64_65_2(twiddle_rsc_0_1_i_q_d, twiddle_rsc_0_22_i_q_d,
            twiddle_rsc_0_0_i_q_d, tmp_21_sva_2, tmp_21_sva_3, twiddle_rsc_0_4_i_q_d,
            tmp_21_sva_5, tmp_21_sva_6, tmp_21_sva_7, twiddle_rsc_0_8_i_q_d, tmp_21_sva_9,
            COMP_LOOP_1_acc_8_itm, tmp_21_sva_11, twiddle_rsc_0_12_i_q_d, tmp_21_sva_13,
            tmp_21_sva_14, tmp_21_sva_15, twiddle_rsc_0_16_i_q_d, tmp_21_sva_17,
            tmp_21_sva_18, tmp_21_sva_19, twiddle_rsc_0_20_i_q_d, tmp_21_sva_21,
            tmp_21_sva_22, tmp_21_sva_23, twiddle_rsc_0_24_i_q_d, tmp_21_sva_25,
            tmp_21_sva_26, tmp_21_sva_27, twiddle_rsc_0_28_i_q_d, tmp_21_sva_29,
            tmp_21_sva_30, tmp_21_sva_31, twiddle_rsc_0_32_i_q_d, tmp_21_sva_33,
            tmp_21_sva_34, tmp_21_sva_35, twiddle_rsc_0_36_i_q_d, tmp_21_sva_37,
            tmp_21_sva_38, tmp_21_sva_39, twiddle_rsc_0_40_i_q_d, tmp_21_sva_41,
            tmp_21_sva_42, tmp_21_sva_43, twiddle_rsc_0_44_i_q_d, tmp_21_sva_45,
            tmp_21_sva_46, tmp_21_sva_47, twiddle_rsc_0_48_i_q_d, tmp_21_sva_49,
            tmp_21_sva_50, tmp_21_sva_51, twiddle_rsc_0_52_i_q_d, tmp_21_sva_53,
            tmp_21_sva_54, tmp_21_sva_55, twiddle_rsc_0_56_i_q_d, tmp_21_sva_57,
            tmp_21_sva_58, tmp_21_sva_59, twiddle_rsc_0_60_i_q_d, tmp_21_sva_61,
            tmp_21_sva_62, tmp_21_sva_63, STD_LOGIC_VECTOR'( and_dcpl_432 & and_dcpl_263
            & COMP_LOOP_tmp_and_89_nl & COMP_LOOP_tmp_and_90_nl & COMP_LOOP_tmp_and_91_nl
            & COMP_LOOP_tmp_and_92_nl & COMP_LOOP_tmp_and_93_nl & COMP_LOOP_tmp_and_94_nl
            & COMP_LOOP_tmp_and_95_nl & COMP_LOOP_tmp_and_96_nl & COMP_LOOP_tmp_and_97_nl
            & COMP_LOOP_tmp_and_98_nl & COMP_LOOP_tmp_and_99_nl & COMP_LOOP_tmp_and_100_nl
            & COMP_LOOP_tmp_and_101_nl & COMP_LOOP_tmp_and_102_nl & COMP_LOOP_tmp_and_103_nl
            & COMP_LOOP_tmp_and_104_nl & COMP_LOOP_tmp_and_105_nl & COMP_LOOP_tmp_and_106_nl
            & COMP_LOOP_tmp_and_107_nl & COMP_LOOP_tmp_and_108_nl & COMP_LOOP_tmp_and_109_nl
            & COMP_LOOP_tmp_and_110_nl & COMP_LOOP_tmp_and_111_nl & COMP_LOOP_tmp_and_112_nl
            & COMP_LOOP_tmp_and_113_nl & COMP_LOOP_tmp_and_114_nl & COMP_LOOP_tmp_and_115_nl
            & COMP_LOOP_tmp_and_116_nl & COMP_LOOP_tmp_and_117_nl & COMP_LOOP_tmp_and_118_nl
            & COMP_LOOP_tmp_and_119_nl & COMP_LOOP_tmp_and_120_nl & COMP_LOOP_tmp_and_121_nl
            & COMP_LOOP_tmp_and_122_nl & COMP_LOOP_tmp_and_123_nl & COMP_LOOP_tmp_and_124_nl
            & COMP_LOOP_tmp_and_125_nl & COMP_LOOP_tmp_and_126_nl & COMP_LOOP_tmp_and_127_nl
            & COMP_LOOP_tmp_and_128_nl & COMP_LOOP_tmp_and_129_nl & COMP_LOOP_tmp_and_130_nl
            & COMP_LOOP_tmp_and_131_nl & COMP_LOOP_tmp_and_132_nl & COMP_LOOP_tmp_and_133_nl
            & COMP_LOOP_tmp_and_134_nl & COMP_LOOP_tmp_and_135_nl & COMP_LOOP_tmp_and_136_nl
            & COMP_LOOP_tmp_and_137_nl & COMP_LOOP_tmp_and_138_nl & COMP_LOOP_tmp_and_139_nl
            & COMP_LOOP_tmp_and_140_nl & COMP_LOOP_tmp_and_141_nl & COMP_LOOP_tmp_and_142_nl
            & COMP_LOOP_tmp_and_143_nl & COMP_LOOP_tmp_and_144_nl & COMP_LOOP_tmp_and_145_nl
            & COMP_LOOP_tmp_and_146_nl & COMP_LOOP_tmp_and_147_nl & COMP_LOOP_tmp_and_148_nl
            & COMP_LOOP_tmp_and_149_nl & COMP_LOOP_tmp_and_150_nl & COMP_LOOP_tmp_and_151_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm = '1' ) THEN
        tmp_21_sva_3 <= twiddle_rsc_0_3_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm = '1' ) THEN
        tmp_21_sva_5 <= twiddle_rsc_0_5_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm = '1' ) THEN
        tmp_21_sva_7 <= twiddle_rsc_0_7_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm = '1' ) THEN
        tmp_21_sva_9 <= twiddle_rsc_0_9_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_COMP_LOOP_and_123_itm = '1' ) THEN
        tmp_21_sva_27 <= twiddle_rsc_0_27_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_COMP_LOOP_and_125_itm = '1' ) THEN
        tmp_21_sva_29 <= twiddle_rsc_0_29_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_COMP_LOOP_and_1831_itm = '1' ) THEN
        tmp_21_sva_31 <= twiddle_rsc_0_31_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_COMP_LOOP_and_1874_itm = '1' ) THEN
        tmp_21_sva_33 <= twiddle_rsc_0_33_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm = '1' ) THEN
        tmp_21_sva_35 <= twiddle_rsc_0_35_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm = '1' ) THEN
        tmp_21_sva_37 <= twiddle_rsc_0_37_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm = '1' ) THEN
        tmp_21_sva_39 <= twiddle_rsc_0_39_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm = '1' ) THEN
        tmp_21_sva_41 <= twiddle_rsc_0_41_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm = '1' ) THEN
        tmp_21_sva_43 <= twiddle_rsc_0_43_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm = '1' ) THEN
        tmp_21_sva_45 <= twiddle_rsc_0_45_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm = '1' ) THEN
        tmp_21_sva_47 <= twiddle_rsc_0_47_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm = '1' ) THEN
        tmp_21_sva_49 <= twiddle_rsc_0_49_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm = '1' ) THEN
        tmp_21_sva_51 <= twiddle_rsc_0_51_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm = '1' ) THEN
        tmp_21_sva_53 <= twiddle_rsc_0_53_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm = '1' ) THEN
        tmp_21_sva_55 <= twiddle_rsc_0_55_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm = '1' ) THEN
        tmp_21_sva_57 <= twiddle_rsc_0_57_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm = '1' ) THEN
        tmp_21_sva_59 <= twiddle_rsc_0_59_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm = '1' ) THEN
        tmp_21_sva_61 <= twiddle_rsc_0_61_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm = '1' ) THEN
        tmp_21_sva_63 <= twiddle_rsc_0_63_i_q_d;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_74_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_75_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_76_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_78_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_79_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_87_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_88_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_89_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_90_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_91_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_92_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_93_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_94_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_95_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_96_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_97_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_98_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_99_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm <= '0';
      ELSIF ( or_dcpl_150 = '0' ) THEN
        COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_3360_tmp = '1' ) THEN
        COMP_LOOP_tmp_mux1h_5_itm <= MUX1HOT_v_64_64_2(twiddle_rsc_0_0_i_q_d, tmp_21_sva_1,
            tmp_21_sva_2, tmp_21_sva_3, twiddle_rsc_0_4_i_q_d, tmp_21_sva_5, tmp_21_sva_6,
            tmp_21_sva_7, twiddle_rsc_0_8_i_q_d, tmp_21_sva_9, COMP_LOOP_1_acc_8_itm,
            tmp_21_sva_11, twiddle_rsc_0_12_i_q_d, tmp_21_sva_13, tmp_21_sva_14,
            tmp_21_sva_15, twiddle_rsc_0_16_i_q_d, tmp_21_sva_17, tmp_21_sva_18,
            tmp_21_sva_19, twiddle_rsc_0_20_i_q_d, tmp_21_sva_21, tmp_21_sva_22,
            tmp_21_sva_23, twiddle_rsc_0_24_i_q_d, tmp_21_sva_25, tmp_21_sva_26,
            tmp_21_sva_27, twiddle_rsc_0_28_i_q_d, tmp_21_sva_29, tmp_21_sva_30,
            tmp_21_sva_31, twiddle_rsc_0_32_i_q_d, tmp_21_sva_33, tmp_21_sva_34,
            tmp_21_sva_35, twiddle_rsc_0_36_i_q_d, tmp_21_sva_37, tmp_21_sva_38,
            tmp_21_sva_39, twiddle_rsc_0_40_i_q_d, tmp_21_sva_41, tmp_21_sva_42,
            tmp_21_sva_43, twiddle_rsc_0_44_i_q_d, tmp_21_sva_45, tmp_21_sva_46,
            tmp_21_sva_47, twiddle_rsc_0_48_i_q_d, tmp_21_sva_49, tmp_21_sva_50,
            tmp_21_sva_51, twiddle_rsc_0_52_i_q_d, tmp_21_sva_53, tmp_21_sva_54,
            tmp_21_sva_55, twiddle_rsc_0_56_i_q_d, tmp_21_sva_57, tmp_21_sva_58,
            tmp_21_sva_59, twiddle_rsc_0_60_i_q_d, tmp_21_sva_61, tmp_21_sva_62,
            tmp_21_sva_63, STD_LOGIC_VECTOR'( COMP_LOOP_tmp_and_31_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_179_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_180_nl & COMP_LOOP_tmp_and_32_nl &
            COMP_LOOP_tmp_COMP_LOOP_tmp_and_182_nl & COMP_LOOP_tmp_and_33_nl & COMP_LOOP_tmp_and_34_nl
            & COMP_LOOP_tmp_and_35_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_186_nl &
            COMP_LOOP_tmp_and_36_nl & COMP_LOOP_tmp_and_37_nl & COMP_LOOP_tmp_and_38_nl
            & COMP_LOOP_tmp_and_39_nl & COMP_LOOP_tmp_and_40_nl & COMP_LOOP_tmp_and_41_nl
            & COMP_LOOP_tmp_and_42_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_and_194_nl &
            COMP_LOOP_tmp_and_43_nl & COMP_LOOP_tmp_and_44_nl & COMP_LOOP_tmp_and_45_nl
            & COMP_LOOP_tmp_and_46_nl & COMP_LOOP_tmp_and_47_nl & COMP_LOOP_tmp_and_48_nl
            & COMP_LOOP_tmp_and_49_nl & COMP_LOOP_tmp_and_50_nl & COMP_LOOP_tmp_and_51_nl
            & COMP_LOOP_tmp_and_52_nl & COMP_LOOP_tmp_and_53_nl & COMP_LOOP_tmp_and_54_nl
            & COMP_LOOP_tmp_and_55_nl & COMP_LOOP_tmp_and_56_nl & COMP_LOOP_tmp_and_57_nl
            & COMP_LOOP_tmp_COMP_LOOP_tmp_and_210_nl & COMP_LOOP_tmp_and_58_nl &
            COMP_LOOP_tmp_and_59_nl & COMP_LOOP_tmp_and_60_nl & COMP_LOOP_tmp_and_61_nl
            & COMP_LOOP_tmp_and_62_nl & COMP_LOOP_tmp_and_63_nl & COMP_LOOP_tmp_and_64_nl
            & COMP_LOOP_tmp_and_65_nl & COMP_LOOP_tmp_and_66_nl & COMP_LOOP_tmp_and_67_nl
            & COMP_LOOP_tmp_and_68_nl & COMP_LOOP_tmp_and_69_nl & COMP_LOOP_tmp_and_70_nl
            & COMP_LOOP_tmp_and_71_nl & COMP_LOOP_tmp_and_72_nl & COMP_LOOP_tmp_and_73_nl
            & COMP_LOOP_tmp_and_74_nl & COMP_LOOP_tmp_and_75_nl & COMP_LOOP_tmp_and_76_nl
            & COMP_LOOP_tmp_and_77_nl & COMP_LOOP_tmp_and_78_nl & COMP_LOOP_tmp_and_79_nl
            & COMP_LOOP_tmp_and_80_nl & COMP_LOOP_tmp_and_81_nl & COMP_LOOP_tmp_and_82_nl
            & COMP_LOOP_tmp_and_83_nl & COMP_LOOP_tmp_and_84_nl & COMP_LOOP_tmp_and_85_nl
            & COMP_LOOP_tmp_and_86_nl & COMP_LOOP_tmp_and_87_nl & COMP_LOOP_tmp_and_88_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (((NOT(COMP_LOOP_tmp_nor_206_itm AND (COMP_LOOP_3_tmp_lshift_ncse_sva(0))))
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_243_rgt
          OR COMP_LOOP_COMP_LOOP_and_119_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_245_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_249_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_257_rgt
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm
          OR COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm OR and_dcpl_263) AND mux_3364_nl)
          = '1' ) THEN
        COMP_LOOP_tmp_mux1h_6_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_0_i_q_d,
            twiddle_rsc_0_4_i_q_d, tmp_21_sva_21, twiddle_rsc_0_8_i_q_d, tmp_21_sva_23,
            twiddle_rsc_0_12_i_q_d, tmp_21_sva_25, twiddle_rsc_0_16_i_q_d, tmp_21_sva_26,
            twiddle_rsc_0_20_i_q_d, tmp_21_sva_1, twiddle_rsc_0_24_i_q_d, COMP_LOOP_1_acc_8_itm,
            twiddle_rsc_0_28_i_q_d, tmp_21_sva_11, twiddle_rsc_0_32_i_q_d, tmp_21_sva_13,
            twiddle_rsc_0_36_i_q_d, tmp_21_sva_14, twiddle_rsc_0_40_i_q_d, tmp_21_sva_15,
            twiddle_rsc_0_44_i_q_d, tmp_21_sva_17, twiddle_rsc_0_48_i_q_d, tmp_21_sva_18,
            twiddle_rsc_0_52_i_q_d, tmp_21_sva_19, twiddle_rsc_0_56_i_q_d, tmp_21_sva_2,
            twiddle_rsc_0_60_i_q_d, tmp_21_sva_22, STD_LOGIC_VECTOR'( and_dcpl_263
            & COMP_LOOP_tmp_and_nl & COMP_LOOP_tmp_and_1_nl & COMP_LOOP_tmp_and_2_nl
            & COMP_LOOP_tmp_and_3_nl & COMP_LOOP_tmp_and_4_nl & COMP_LOOP_tmp_and_5_nl
            & COMP_LOOP_tmp_and_6_nl & COMP_LOOP_tmp_and_7_nl & COMP_LOOP_tmp_and_8_nl
            & COMP_LOOP_tmp_and_9_nl & COMP_LOOP_tmp_and_10_nl & COMP_LOOP_tmp_and_11_nl
            & COMP_LOOP_tmp_and_12_nl & COMP_LOOP_tmp_and_13_nl & COMP_LOOP_tmp_and_14_nl
            & COMP_LOOP_tmp_and_15_nl & COMP_LOOP_tmp_and_16_nl & COMP_LOOP_tmp_and_17_nl
            & COMP_LOOP_tmp_and_18_nl & COMP_LOOP_tmp_and_19_nl & COMP_LOOP_tmp_and_20_nl
            & COMP_LOOP_tmp_and_21_nl & COMP_LOOP_tmp_and_22_nl & COMP_LOOP_tmp_and_23_nl
            & COMP_LOOP_tmp_and_24_nl & COMP_LOOP_tmp_and_25_nl & COMP_LOOP_tmp_and_26_nl
            & COMP_LOOP_tmp_and_27_nl & COMP_LOOP_tmp_and_28_nl & COMP_LOOP_tmp_and_29_nl
            & COMP_LOOP_tmp_and_30_nl));
      END IF;
    END IF;
  END PROCESS;
  nor_1423_nl <= NOT((fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(4))
      OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_788_nl <= MUX_s_1_2_2(and_tmp_29, and_78_cse, fsm_output(2));
  mux_789_nl <= MUX_s_1_2_2(mux_788_nl, mux_tmp_720, fsm_output(1));
  VEC_LOOP_j_not_1_nl <= NOT VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  nor_422_nl <= NOT((fsm_output(1)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(4))
      OR (fsm_output(3)) OR (fsm_output(7)));
  nor_1426_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(7)));
  and_637_nl <= (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(7));
  mux_781_nl <= MUX_s_1_2_2(nor_1426_nl, and_637_nl, fsm_output(5));
  nand_480_nl <= NOT(mux_781_nl AND and_dcpl_365 AND (NOT (fsm_output(4))) AND (NOT
      (fsm_output(2))));
  or_4159_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 4)/=STD_LOGIC_VECTOR'("000")) OR
      nor_1744_cse OR (fsm_output(3));
  nor_1745_nl <= NOT((CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111")))
      OR (fsm_output(3)));
  or_4154_nl <= (fsm_output(2)) OR and_1046_cse OR (fsm_output(3));
  mux_nl <= MUX_s_1_2_2(nor_1745_nl, or_4154_nl, fsm_output(5));
  mux_3365_nl <= MUX_s_1_2_2(mux_nl, (fsm_output(5)), fsm_output(4));
  nand_493_nl <= NOT((fsm_output(6)) AND (NOT mux_3365_nl));
  COMP_LOOP_COMP_LOOP_and_73_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001011"));
  COMP_LOOP_COMP_LOOP_and_824_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_4_sva(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_734_itm;
  COMP_LOOP_COMP_LOOP_and_74_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001100"));
  COMP_LOOP_COMP_LOOP_and_851_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_4_sva(0))
      AND COMP_LOOP_nor_760_itm;
  COMP_LOOP_COMP_LOOP_and_75_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001101"));
  COMP_LOOP_COMP_LOOP_and_858_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_4_sva(3))
      AND COMP_LOOP_nor_767_itm;
  COMP_LOOP_COMP_LOOP_and_100_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("100110"));
  COMP_LOOP_COMP_LOOP_and_323_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_2_sva(0))
      AND COMP_LOOP_nor_289_itm;
  COMP_LOOP_COMP_LOOP_and_1073_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_955_itm;
  mux_3036_nl <= MUX_s_1_2_2(mux_tmp_2968, mux_tmp_2966, fsm_output(1));
  mux_3037_nl <= MUX_s_1_2_2(or_4057_cse, (NOT mux_3036_nl), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_101_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("100111"));
  COMP_LOOP_COMP_LOOP_and_348_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_2_sva(1))
      AND COMP_LOOP_nor_313_itm;
  COMP_LOOP_COMP_LOOP_and_1075_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(2)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(0))
      AND COMP_LOOP_nor_957_itm;
  and_403_nl <= and_dcpl_76 AND and_dcpl_88;
  nor_420_nl <= NOT(and_507_cse OR (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(3)));
  mux_3039_nl <= MUX_s_1_2_2(nor_420_nl, mux_tmp_2971, fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_102_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("101000"));
  COMP_LOOP_COMP_LOOP_and_1076_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_958_itm;
  COMP_LOOP_COMP_LOOP_and_109_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("101111"));
  COMP_LOOP_COMP_LOOP_and_1094_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(4
      DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_976_itm;
  COMP_LOOP_COMP_LOOP_and_103_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("101001"));
  COMP_LOOP_COMP_LOOP_and_350_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_2_sva(2))
      AND COMP_LOOP_nor_315_itm;
  COMP_LOOP_COMP_LOOP_and_1079_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(0))
      AND COMP_LOOP_nor_961_itm;
  mux_3046_nl <= MUX_s_1_2_2(or_4057_cse, (NOT mux_tmp_2968), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_104_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("101010"));
  COMP_LOOP_COMP_LOOP_and_354_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_2_sva(3))
      AND COMP_LOOP_nor_319_itm;
  COMP_LOOP_COMP_LOOP_and_1080_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(1))
      AND COMP_LOOP_nor_962_itm;
  and_409_nl <= and_dcpl_76 AND and_dcpl_377;
  mux_3047_nl <= MUX_s_1_2_2(or_tmp_3747, (NOT mux_tmp_2966), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_105_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("101011"));
  COMP_LOOP_COMP_LOOP_and_362_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_2_sva(5
      DOWNTO 4)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_326_itm;
  COMP_LOOP_COMP_LOOP_and_1082_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(3
      DOWNTO 2)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_964_itm;
  mux_3048_nl <= MUX_s_1_2_2(or_tmp_3747, (NOT mux_tmp_2968), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_106_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("101100"));
  COMP_LOOP_COMP_LOOP_and_1087_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(0))
      AND COMP_LOOP_nor_969_itm;
  and_411_nl <= and_dcpl_94 AND and_dcpl_113;
  or_3878_nl <= and_507_cse OR (fsm_output(6));
  or_3877_nl <= nor_1744_cse OR (fsm_output(6));
  mux_3051_nl <= MUX_s_1_2_2(or_3878_nl, or_3877_nl, fsm_output(3));
  mux_3052_nl <= MUX_s_1_2_2((fsm_output(6)), mux_3051_nl, nor_358_cse);
  nor_418_nl <= NOT((fsm_output(1)) OR (fsm_output(6)));
  or_3874_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  mux_3049_nl <= MUX_s_1_2_2(nor_418_nl, (fsm_output(6)), or_3874_nl);
  mux_3050_nl <= MUX_s_1_2_2((fsm_output(6)), (NOT mux_3049_nl), fsm_output(5));
  mux_3053_nl <= MUX_s_1_2_2(mux_3052_nl, mux_3050_nl, fsm_output(4));
  COMP_LOOP_COMP_LOOP_and_107_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("101101"));
  COMP_LOOP_COMP_LOOP_and_1088_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(1))
      AND COMP_LOOP_nor_970_itm;
  mux_3055_nl <= MUX_s_1_2_2((NOT and_640_cse), and_640_cse, fsm_output(6));
  mux_3054_nl <= MUX_s_1_2_2((NOT and_640_cse), (fsm_output(4)), fsm_output(6));
  mux_3056_nl <= MUX_s_1_2_2(mux_3055_nl, mux_3054_nl, fsm_output(2));
  mux_3059_nl <= MUX_s_1_2_2((NOT mux_3058_itm), mux_3056_nl, fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_108_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("101110"));
  COMP_LOOP_COMP_LOOP_and_1090_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      AND COMP_LOOP_nor_972_itm;
  mux_3062_nl <= MUX_s_1_2_2(mux_tmp_2994, mux_tmp_2993, fsm_output(1));
  mux_3063_nl <= MUX_s_1_2_2(mux_3062_nl, (NOT mux_180_cse), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_110_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("110000"));
  COMP_LOOP_COMP_LOOP_and_1103_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(0))
      AND COMP_LOOP_nor_984_itm;
  mux_3064_nl <= MUX_s_1_2_2((NOT mux_3058_itm), mux_tmp_2968, fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_115_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("110101"));
  COMP_LOOP_COMP_LOOP_and_1328_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1182_itm;
  COMP_LOOP_COMP_LOOP_and_117_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("110111"));
  COMP_LOOP_COMP_LOOP_and_1332_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(1))
      AND COMP_LOOP_nor_1186_itm;
  COMP_LOOP_COMP_LOOP_and_122_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("111100"));
  COMP_LOOP_COMP_LOOP_and_1355_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(0))
      AND COMP_LOOP_nor_1208_itm;
  COMP_LOOP_COMP_LOOP_and_116_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("110110"));
  COMP_LOOP_COMP_LOOP_and_1331_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(0))
      AND COMP_LOOP_nor_1185_itm;
  or_3889_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_3073_nl <= MUX_s_1_2_2(or_3889_nl, mux_742_cse, fsm_output(2));
  COMP_LOOP_COMP_LOOP_and_118_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("111000"));
  COMP_LOOP_COMP_LOOP_and_1334_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(3
      DOWNTO 2)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1188_itm;
  mux_3081_nl <= MUX_s_1_2_2(mux_tmp_3013, mux_tmp_3012, fsm_output(1));
  COMP_LOOP_COMP_LOOP_and_119_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("111001"));
  COMP_LOOP_COMP_LOOP_and_1339_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(0))
      AND COMP_LOOP_nor_1193_itm;
  nor_414_nl <= NOT((NOT((fsm_output(0)) OR (NOT (fsm_output(3))))) OR (fsm_output(7)));
  mux_3084_nl <= MUX_s_1_2_2(nor_414_nl, (fsm_output(7)), or_341_cse);
  mux_3085_nl <= MUX_s_1_2_2(mux_3084_nl, mux_tmp_3016, or_359_cse);
  COMP_LOOP_COMP_LOOP_and_120_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("111010"));
  COMP_LOOP_COMP_LOOP_and_1340_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(1))
      AND COMP_LOOP_nor_1194_itm;
  mux_3090_nl <= MUX_s_1_2_2((NOT or_tmp_3760), (fsm_output(7)), or_341_cse);
  mux_3091_nl <= MUX_s_1_2_2(mux_3090_nl, mux_tmp_206, fsm_output(2));
  mux_3087_nl <= MUX_s_1_2_2((NOT or_tmp_3757), (fsm_output(7)), or_341_cse);
  mux_3089_nl <= MUX_s_1_2_2(mux_tmp_206, mux_3087_nl, fsm_output(2));
  mux_3092_nl <= MUX_s_1_2_2(mux_3091_nl, mux_3089_nl, fsm_output(1));
  COMP_LOOP_COMP_LOOP_and_121_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("111011"));
  COMP_LOOP_COMP_LOOP_and_1342_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(2))
      AND COMP_LOOP_nor_1196_itm;
  and_503_nl <= (fsm_output(3)) AND (NOT or_tmp_3773);
  mux_3096_nl <= MUX_s_1_2_2(mux_3095_cse, and_503_nl, fsm_output(5));
  mux_3097_nl <= MUX_s_1_2_2(mux_3096_nl, nor_412_cse, fsm_output(4));
  COMP_LOOP_COMP_LOOP_and_123_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("111101"));
  COMP_LOOP_COMP_LOOP_and_1356_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(1))
      AND COMP_LOOP_nor_1209_itm;
  COMP_LOOP_COMP_LOOP_and_124_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("111110"));
  COMP_LOOP_COMP_LOOP_and_1358_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(2))
      AND COMP_LOOP_nor_1211_itm;
  or_3904_nl <= (fsm_output(5)) OR (NOT mux_3095_cse);
  nand_145_nl <= NOT((fsm_output(5)) AND (fsm_output(3)) AND (NOT or_tmp_3773));
  mux_3102_nl <= MUX_s_1_2_2(or_3904_nl, nand_145_nl, fsm_output(4));
  COMP_LOOP_COMP_LOOP_and_125_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("111111"));
  COMP_LOOP_COMP_LOOP_and_1362_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_6_sva(3))
      AND COMP_LOOP_nor_1215_itm;
  mux_3104_nl <= MUX_s_1_2_2((NOT or_tmp_3760), or_tmp_118, fsm_output(4));
  mux_3105_nl <= MUX_s_1_2_2(mux_3104_nl, (fsm_output(7)), fsm_output(6));
  mux_3106_nl <= MUX_s_1_2_2(mux_3105_nl, mux_tmp_444, fsm_output(2));
  mux_3107_nl <= MUX_s_1_2_2(mux_3106_nl, mux_tmp_3012, fsm_output(1));
  mux_3110_nl <= MUX_s_1_2_2(mux_tmp_2955, and_78_cse, fsm_output(2));
  mux_3111_nl <= MUX_s_1_2_2(mux_3110_nl, mux_tmp_3042, fsm_output(1));
  mux_3113_nl <= MUX_s_1_2_2(and_tmp_31, and_673_cse, or_359_cse);
  mux_3115_nl <= MUX_s_1_2_2((NOT mux_3114_itm), mux_3113_nl, fsm_output(5));
  mux_3123_nl <= MUX_s_1_2_2(mux_221_cse, (NOT and_640_cse), fsm_output(5));
  COMP_LOOP_3_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & STD_LOGIC_VECTOR'( "010")), 10), 11) + SIGNED'( "00000000001"), 11));
  nand_149_nl <= NOT(or_359_cse AND CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")));
  mux_3124_nl <= MUX_s_1_2_2(mux_221_cse, nand_149_nl, fsm_output(5));
  mux_3125_nl <= MUX_s_1_2_2(mux_tmp_2971, mux_tmp_3049, fsm_output(1));
  mux_3126_nl <= MUX_s_1_2_2(mux_3125_nl, (fsm_output(6)), fsm_output(5));
  COMP_LOOP_acc_12_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 3)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & '0'), 8), 9) + UNSIGNED'( "000000001"), 9));
  mux_3127_nl <= MUX_s_1_2_2(mux_tmp_2960, mux_tmp_3049, fsm_output(1));
  mux_3128_nl <= MUX_s_1_2_2(mux_3127_nl, (fsm_output(6)), fsm_output(5));
  mux_3130_nl <= MUX_s_1_2_2((NOT mux_3114_itm), and_673_cse, fsm_output(5));
  COMP_LOOP_5_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & STD_LOGIC_VECTOR'( "100")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_3131_nl <= MUX_s_1_2_2(and_677_cse, and_673_cse, or_359_cse);
  mux_3132_nl <= MUX_s_1_2_2((NOT mux_3114_itm), mux_3131_nl, fsm_output(5));
  and_497_nl <= (fsm_output(0)) AND (fsm_output(3)) AND (fsm_output(7));
  mux_3138_nl <= MUX_s_1_2_2(and_497_nl, (fsm_output(7)), or_341_cse);
  mux_3139_nl <= MUX_s_1_2_2(mux_tmp_3016, mux_3138_nl, fsm_output(2));
  mux_3140_nl <= MUX_s_1_2_2(mux_3139_nl, mux_tmp_3070, fsm_output(1));
  mux_3142_nl <= MUX_s_1_2_2(mux_tmp_3016, and_736_cse, fsm_output(2));
  mux_3143_nl <= MUX_s_1_2_2(mux_3142_nl, mux_tmp_3070, fsm_output(1));
  COMP_LOOP_6_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & STD_LOGIC_VECTOR'( "101")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_3146_nl <= MUX_s_1_2_2(mux_tmp_3078, mux_tmp_3070, fsm_output(1));
  mux_212_nl <= MUX_s_1_2_2(and_tmp_10, (fsm_output(4)), or_359_cse);
  mux_3152_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_212_nl), fsm_output(5));
  mux_219_nl <= MUX_s_1_2_2(or_595_cse, or_4007_cse, and_507_cse);
  mux_3160_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_219_nl), fsm_output(5));
  nor_410_nl <= NOT(and_1046_cse OR (fsm_output(5)) OR (fsm_output(7)));
  and_491_nl <= (CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))) AND
      (fsm_output(5)) AND (fsm_output(7));
  mux_3161_nl <= MUX_s_1_2_2(nor_410_nl, and_491_nl, fsm_output(3));
  and_492_nl <= (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(7));
  mux_3162_nl <= MUX_s_1_2_2(mux_3161_nl, and_492_nl, fsm_output(2));
  mux_3163_nl <= MUX_s_1_2_2(mux_3162_nl, and_493_cse, fsm_output(4));
  COMP_LOOP_7_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))) + CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0
      & STD_LOGIC_VECTOR'( "110")), 10), 11) + SIGNED'( "00000000001"), 11));
  mux_3171_nl <= MUX_s_1_2_2(nor_tmp_99, and_736_cse, or_359_cse);
  mux_3181_nl <= MUX_s_1_2_2(mux_tmp_2955, and_705_cse, fsm_output(2));
  mux_3182_nl <= MUX_s_1_2_2(mux_3181_nl, mux_tmp_3042, fsm_output(1));
  COMP_LOOP_acc_15_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 4)))) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_10_3_sva_6_0),
      7), 8) + UNSIGNED'( "00000001"), 8));
  nand_148_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 0)=STD_LOGIC_VECTOR'("11111")));
  mux_3188_nl <= MUX_s_1_2_2(mux_221_cse, nand_148_nl, fsm_output(5));
  mux_359_nl <= MUX_s_1_2_2(and_tmp_10, (fsm_output(4)), fsm_output(2));
  mux_361_nl <= MUX_s_1_2_2(mux_tmp_293, mux_359_nl, fsm_output(1));
  mux_3192_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_361_nl), fsm_output(5));
  mux_3193_nl <= MUX_s_1_2_2(and_78_cse, and_705_cse, or_359_cse);
  COMP_LOOP_1_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(z_out_2 & STD_LOGIC_VECTOR'(
      "000")) + SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10 DOWNTO 1)))) + SIGNED'(
      "00000000001"), 11));
  mux_3197_nl <= MUX_s_1_2_2(and_tmp_29, and_705_cse, or_359_cse);
  and_489_nl <= (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0)) AND (fsm_output(3));
  mux_3203_nl <= MUX_s_1_2_2((NOT or_4057_cse), and_489_nl, fsm_output(2));
  mux_3202_nl <= MUX_s_1_2_2((NOT or_tmp_3801), and_677_cse, fsm_output(2));
  mux_3204_nl <= MUX_s_1_2_2(mux_3203_nl, mux_3202_nl, fsm_output(1));
  mux_3205_nl <= MUX_s_1_2_2(mux_3204_nl, (fsm_output(6)), fsm_output(5));
  and_449_nl <= (fsm_output(6)) AND or_tmp_105;
  mux_3208_nl <= MUX_s_1_2_2(mux_tmp_2965, and_449_nl, fsm_output(2));
  mux_3206_nl <= MUX_s_1_2_2((NOT or_4007_cse), (fsm_output(4)), fsm_output(6));
  mux_3207_nl <= MUX_s_1_2_2(mux_3206_nl, and_tmp_33, fsm_output(2));
  mux_3209_nl <= MUX_s_1_2_2(mux_3208_nl, mux_3207_nl, fsm_output(1));
  mux_3210_nl <= MUX_s_1_2_2(mux_3209_nl, (fsm_output(6)), fsm_output(5));
  mux_3213_nl <= MUX_s_1_2_2((NOT or_595_cse), or_tmp_105, fsm_output(6));
  mux_3214_nl <= MUX_s_1_2_2(mux_3213_nl, and_tmp_33, fsm_output(2));
  mux_3211_nl <= MUX_s_1_2_2((NOT or_4007_cse), or_595_cse, fsm_output(6));
  mux_3212_nl <= MUX_s_1_2_2(mux_3211_nl, and_tmp_33, fsm_output(2));
  mux_3215_nl <= MUX_s_1_2_2(mux_3214_nl, mux_3212_nl, fsm_output(1));
  mux_3216_nl <= MUX_s_1_2_2(mux_3215_nl, (fsm_output(6)), fsm_output(5));
  mux_434_nl <= MUX_s_1_2_2(and_640_cse, and_tmp_10, fsm_output(2));
  mux_435_nl <= MUX_s_1_2_2(mux_434_nl, mux_tmp_293, fsm_output(1));
  mux_3219_nl <= MUX_s_1_2_2(mux_221_cse, (NOT mux_435_nl), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_111_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("110001"));
  COMP_LOOP_COMP_LOOP_and_1104_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(1))
      AND COMP_LOOP_nor_985_itm;
  or_3932_nl <= (fsm_output(6)) OR (fsm_output(4)) OR and_639_cse;
  mux_3221_nl <= MUX_s_1_2_2(or_3932_nl, or_341_cse, fsm_output(2));
  or_3929_nl <= (fsm_output(6)) OR (fsm_output(4)) OR and_dcpl_365;
  mux_3220_nl <= MUX_s_1_2_2(or_341_cse, or_3929_nl, fsm_output(2));
  mux_3222_nl <= MUX_s_1_2_2(mux_3221_nl, mux_3220_nl, fsm_output(1));
  mux_3223_nl <= MUX_s_1_2_2(mux_3222_nl, (NOT mux_180_cse), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_112_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("110010"));
  COMP_LOOP_COMP_LOOP_and_1106_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(2))
      AND COMP_LOOP_nor_987_itm;
  or_3934_nl <= (fsm_output(6)) OR (((fsm_output(4)) OR (fsm_output(0))) AND (fsm_output(3)));
  mux_3224_nl <= MUX_s_1_2_2(or_3934_nl, or_4050_cse, fsm_output(2));
  mux_3225_nl <= MUX_s_1_2_2(mux_3224_nl, mux_tmp_2993, fsm_output(1));
  mux_3226_nl <= MUX_s_1_2_2(mux_3225_nl, (NOT mux_180_cse), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_113_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("110011"));
  COMP_LOOP_COMP_LOOP_and_1110_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_5_sva(3))
      AND COMP_LOOP_nor_991_itm;
  mux_3227_nl <= MUX_s_1_2_2(or_4057_cse, (NOT mux_180_cse), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_114_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("110100"));
  COMP_LOOP_COMP_LOOP_and_1118_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_5_sva(5
      DOWNTO 4)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_998_itm;
  mux_3228_nl <= MUX_s_1_2_2(mux_tmp_2994, mux_tmp_2975, fsm_output(1));
  mux_3229_nl <= MUX_s_1_2_2(mux_3228_nl, (NOT mux_180_cse), fsm_output(5));
  COMP_LOOP_COMP_LOOP_and_65_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("000011"));
  COMP_LOOP_COMP_LOOP_and_1370_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_6_sva(5
      DOWNTO 4)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1222_itm;
  mux_3230_nl <= MUX_s_1_2_2(mux_tmp_656, mux_tmp_3009, fsm_output(2));
  mux_3231_nl <= MUX_s_1_2_2(mux_tmp_3013, mux_3230_nl, fsm_output(1));
  COMP_LOOP_COMP_LOOP_and_67_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("000101"));
  COMP_LOOP_COMP_LOOP_and_1577_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1403_itm;
  COMP_LOOP_COMP_LOOP_and_68_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("000110"));
  COMP_LOOP_COMP_LOOP_and_1584_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(1))
      AND COMP_LOOP_nor_1410_itm;
  COMP_LOOP_COMP_LOOP_and_317_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("000011"));
  COMP_LOOP_COMP_LOOP_and_1594_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      AND COMP_LOOP_nor_1420_itm;
  COMP_LOOP_COMP_LOOP_and_324_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001010"));
  COMP_LOOP_COMP_LOOP_and_1614_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(3))
      AND COMP_LOOP_nor_1439_itm;
  COMP_LOOP_COMP_LOOP_and_319_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("000101"));
  COMP_LOOP_COMP_LOOP_and_1598_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(4
      DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1424_itm;
  nor_403_nl <= NOT((NOT((NOT (fsm_output(3))) OR (fsm_output(5)))) OR (fsm_output(7)));
  nor_405_nl <= NOT((fsm_output(3)) OR nor_358_cse OR (fsm_output(7)));
  mux_3241_nl <= MUX_s_1_2_2(nor_403_nl, nor_405_nl, fsm_output(1));
  mux_3240_nl <= MUX_s_1_2_2(nor_412_cse, and_493_cse, fsm_output(3));
  mux_3242_nl <= MUX_s_1_2_2(mux_3241_nl, mux_3240_nl, fsm_output(2));
  mux_3243_nl <= MUX_s_1_2_2(mux_3242_nl, and_493_cse, fsm_output(4));
  COMP_LOOP_COMP_LOOP_and_320_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("000110"));
  COMP_LOOP_COMP_LOOP_and_1607_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(0))
      AND COMP_LOOP_nor_1432_itm;
  and_458_nl <= and_dcpl_94 AND and_dcpl_88;
  mux_3245_nl <= MUX_s_1_2_2(or_tmp_3717, (fsm_output(7)), or_341_cse);
  mux_3246_nl <= MUX_s_1_2_2(mux_tmp_444, mux_3245_nl, fsm_output(2));
  COMP_LOOP_COMP_LOOP_and_321_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("000111"));
  COMP_LOOP_COMP_LOOP_and_1610_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_7_sva(2))
      AND COMP_LOOP_nor_1435_itm;
  or_3946_nl <= (NOT((NOT (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(5))))
      OR (fsm_output(7));
  mux_3251_nl <= MUX_s_1_2_2(or_3946_nl, or_564_cse, fsm_output(2));
  mux_582_nl <= MUX_s_1_2_2((NOT or_564_cse), (fsm_output(5)), fsm_output(2));
  mux_3252_nl <= MUX_s_1_2_2((NOT mux_3251_nl), mux_582_nl, fsm_output(3));
  mux_3253_nl <= MUX_s_1_2_2(mux_3252_nl, (fsm_output(5)), fsm_output(4));
  or_3943_nl <= (NOT(and_507_cse OR (fsm_output(5)))) OR (fsm_output(7));
  mux_3248_nl <= MUX_s_1_2_2(or_3943_nl, (fsm_output(7)), fsm_output(3));
  mux_3249_nl <= MUX_s_1_2_2(or_564_cse, mux_3248_nl, fsm_output(4));
  COMP_LOOP_COMP_LOOP_and_325_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001011"));
  COMP_LOOP_COMP_LOOP_and_1622_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_7_sva(5
      DOWNTO 4)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1446_itm;
  and_459_nl <= and_dcpl_85 AND and_dcpl_377;
  mux_3255_nl <= MUX_s_1_2_2(or_tmp_404, (fsm_output(7)), fsm_output(6));
  mux_3256_nl <= MUX_s_1_2_2(mux_tmp_656, mux_3255_nl, fsm_output(2));
  COMP_LOOP_COMP_LOOP_and_69_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("000111"));
  COMP_LOOP_COMP_LOOP_and_1831_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(2)) AND (COMP_LOOP_acc_10_cse_10_1_sva(0))
      AND COMP_LOOP_nor_1629_itm;
  mux_3258_nl <= MUX_s_1_2_2(or_tmp_3757, or_tmp_119, fsm_output(4));
  mux_3259_nl <= MUX_s_1_2_2((NOT mux_3258_nl), and_655_cse, fsm_output(6));
  mux_3261_nl <= MUX_s_1_2_2(mux_tmp_3193, mux_3259_nl, fsm_output(2));
  mux_3264_nl <= MUX_s_1_2_2(mux_tmp_3196, mux_3261_nl, fsm_output(1));
  COMP_LOOP_COMP_LOOP_and_326_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001100"));
  COMP_LOOP_COMP_LOOP_and_1832_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1630_itm;
  and_461_nl <= and_dcpl_94 AND and_dcpl_344;
  mux_3271_nl <= MUX_s_1_2_2(nor_399_cse, mux_297_cse, fsm_output(5));
  mux_3272_nl <= MUX_s_1_2_2(mux_3271_nl, and_tmp_35, and_1046_cse);
  mux_3270_nl <= MUX_s_1_2_2(and_705_cse, mux_297_cse, fsm_output(5));
  mux_3273_nl <= MUX_s_1_2_2(mux_3272_nl, mux_3270_nl, fsm_output(4));
  nor_386_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))));
  mux_3268_nl <= MUX_s_1_2_2(and_705_cse, mux_297_cse, nor_386_nl);
  mux_3269_nl <= MUX_s_1_2_2(and_tmp_35, mux_3268_nl, fsm_output(4));
  mux_3274_nl <= MUX_s_1_2_2(mux_3273_nl, mux_3269_nl, fsm_output(2));
  nor_384_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("10")));
  mux_3267_nl <= MUX_s_1_2_2(and_705_cse, mux_297_cse, nor_384_nl);
  COMP_LOOP_COMP_LOOP_and_327_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001101"));
  COMP_LOOP_COMP_LOOP_and_1835_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(3)) AND (COMP_LOOP_acc_10_cse_10_1_sva(0))
      AND COMP_LOOP_nor_1633_itm;
  and_463_nl <= and_dcpl_264 AND and_dcpl_347;
  mux_3282_nl <= MUX_s_1_2_2(mux_tmp_3214, and_tmp_36, fsm_output(2));
  mux_3278_nl <= MUX_s_1_2_2(and_dcpl_60, mux_tmp_3210, fsm_output(6));
  mux_3279_nl <= MUX_s_1_2_2(mux_3278_nl, and_tmp_36, fsm_output(2));
  mux_3283_nl <= MUX_s_1_2_2(mux_3282_nl, mux_3279_nl, fsm_output(1));
  COMP_LOOP_COMP_LOOP_and_328_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001110"));
  COMP_LOOP_COMP_LOOP_and_1844_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_sva(1))
      AND COMP_LOOP_nor_1642_itm;
  mux_3286_nl <= MUX_s_1_2_2(mux_297_cse, mux_tmp_3218, fsm_output(2));
  COMP_LOOP_COMP_LOOP_and_329_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001111"));
  COMP_LOOP_COMP_LOOP_and_1850_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(4
      DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1648_itm;
  COMP_LOOP_COMP_LOOP_and_331_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010001"));
  COMP_LOOP_COMP_LOOP_and_1862_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_sva(2))
      AND COMP_LOOP_nor_1659_itm;
  and_465_nl <= and_dcpl_264 AND and_dcpl_116;
  and_464_nl <= (fsm_output(6)) AND mux_tmp_3213;
  mux_3291_nl <= MUX_s_1_2_2(mux_tmp_3214, and_464_nl, fsm_output(2));
  mux_3289_nl <= MUX_s_1_2_2(and_dcpl_60, mux_tmp_3213, fsm_output(6));
  mux_3290_nl <= MUX_s_1_2_2(mux_3289_nl, and_tmp_36, fsm_output(2));
  mux_3292_nl <= MUX_s_1_2_2(mux_3291_nl, mux_3290_nl, fsm_output(1));
  COMP_LOOP_COMP_LOOP_and_332_nl <= CONV_SL_1_1(COMP_LOOP_2_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010010"));
  COMP_LOOP_COMP_LOOP_and_1866_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(5)) AND (COMP_LOOP_acc_10_cse_10_1_sva(3))
      AND COMP_LOOP_nor_1663_itm;
  and_468_nl <= and_dcpl_85 AND and_dcpl_116;
  mux_3296_nl <= MUX_s_1_2_2((NOT or_477_cse), or_tmp_404, fsm_output(6));
  and_73_nl <= (fsm_output(6)) AND or_tmp_404;
  mux_3297_nl <= MUX_s_1_2_2(mux_3296_nl, and_73_nl, fsm_output(2));
  mux_3294_nl <= MUX_s_1_2_2(and_dcpl_60, or_tmp_404, fsm_output(6));
  and_466_nl <= (fsm_output(6)) AND mux_tmp_3169;
  mux_3295_nl <= MUX_s_1_2_2(mux_3294_nl, and_466_nl, fsm_output(2));
  mux_3298_nl <= MUX_s_1_2_2(mux_3297_nl, mux_3295_nl, fsm_output(1));
  COMP_LOOP_COMP_LOOP_and_71_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001001"));
  COMP_LOOP_COMP_LOOP_and_1874_nl <= CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_sva(5
      DOWNTO 4)=STD_LOGIC_VECTOR'("11")) AND COMP_LOOP_nor_1670_itm;
  nor_397_nl <= NOT(nor_398_cse OR (fsm_output(7)));
  mux_3300_nl <= MUX_s_1_2_2(nor_397_nl, and_655_cse, fsm_output(6));
  mux_3301_nl <= MUX_s_1_2_2(mux_tmp_3193, mux_3300_nl, fsm_output(2));
  mux_3302_nl <= MUX_s_1_2_2(mux_tmp_3196, mux_3301_nl, fsm_output(1));
  COMP_LOOP_COMP_LOOP_and_72_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001010"));
  COMP_LOOP_COMP_LOOP_and_583_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(4)) AND (COMP_LOOP_acc_10_cse_10_1_3_sva(0))
      AND COMP_LOOP_nor_521_itm;
  mux_3306_nl <= MUX_s_1_2_2(mux_3305_itm, (NOT and_779_cse), fsm_output(5));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_nl <= CONV_SL_1_1(z_out_8(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl <= CONV_SL_1_1(z_out_8(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_nl <= CONV_SL_1_1(z_out_8(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_nl <= CONV_SL_1_1(z_out_8(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_nor_nl <= NOT(CONV_SL_1_1(z_out_8(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  COMP_LOOP_COMP_LOOP_and_76_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001110"));
  COMP_LOOP_COMP_LOOP_and_77_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("001111"));
  COMP_LOOP_COMP_LOOP_and_79_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010001"));
  COMP_LOOP_COMP_LOOP_and_80_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010010"));
  COMP_LOOP_COMP_LOOP_and_81_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010011"));
  COMP_LOOP_COMP_LOOP_and_82_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010100"));
  COMP_LOOP_COMP_LOOP_and_83_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010101"));
  COMP_LOOP_COMP_LOOP_and_84_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010110"));
  COMP_LOOP_COMP_LOOP_and_85_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("010111"));
  COMP_LOOP_COMP_LOOP_and_86_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("011000"));
  COMP_LOOP_COMP_LOOP_and_87_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("011001"));
  COMP_LOOP_COMP_LOOP_and_88_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("011010"));
  COMP_LOOP_COMP_LOOP_and_89_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("011011"));
  COMP_LOOP_COMP_LOOP_and_90_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("011100"));
  COMP_LOOP_COMP_LOOP_and_91_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("011101"));
  COMP_LOOP_COMP_LOOP_and_92_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("011110"));
  COMP_LOOP_COMP_LOOP_and_93_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("011111"));
  COMP_LOOP_COMP_LOOP_and_95_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("100001"));
  COMP_LOOP_COMP_LOOP_and_96_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("100010"));
  COMP_LOOP_COMP_LOOP_and_97_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("100011"));
  COMP_LOOP_COMP_LOOP_and_98_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("100100"));
  COMP_LOOP_COMP_LOOP_and_99_nl <= CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO
      0)=STD_LOGIC_VECTOR'("100101"));
  COMP_LOOP_COMP_LOOP_nor_1_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000000")));
  COMP_LOOP_nor_57_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(5 DOWNTO 1)/=STD_LOGIC_VECTOR'("00000")));
  COMP_LOOP_nor_58_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(4))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(2))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_60_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(4))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(3)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(1))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_64_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(4))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(1))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_72_nl <= NOT((COMP_LOOP_1_acc_10_itm_10_1_1(5)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(3))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(2)) OR (COMP_LOOP_1_acc_10_itm_10_1_1(1))
      OR (COMP_LOOP_1_acc_10_itm_10_1_1(0)));
  COMP_LOOP_nor_87_nl <= NOT(CONV_SL_1_1(COMP_LOOP_1_acc_10_itm_10_1_1(4 DOWNTO 0)/=STD_LOGIC_VECTOR'("00000")));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl <= CONV_SL_1_1(COMP_LOOP_1_tmp_mul_idiv_sva_2_0=STD_LOGIC_VECTOR'("001"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl <= CONV_SL_1_1(COMP_LOOP_1_tmp_mul_idiv_sva_2_0=STD_LOGIC_VECTOR'("010"));
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl <= CONV_SL_1_1(COMP_LOOP_1_tmp_mul_idiv_sva_2_0=STD_LOGIC_VECTOR'("100"));
  COMP_LOOP_COMP_LOOP_mux_21_nl <= MUX_v_64_2_2(COMP_LOOP_1_acc_8_itm, z_out_9, COMP_LOOP_or_65_itm);
  COMP_LOOP_acc_17_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_724_cse)
      + UNSIGNED(COMP_LOOP_COMP_LOOP_mux_21_nl), 64));
  COMP_LOOP_or_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm AND and_dcpl_77) OR
      (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_61_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_60_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_59_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_58_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_57_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_56_itm AND and_dcpl_109);
  COMP_LOOP_or_1_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(0)) AND COMP_LOOP_tmp_nor_10_itm
      AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_61_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_60_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_59_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_58_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_57_itm AND and_dcpl_109);
  COMP_LOOP_or_2_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(1)) AND COMP_LOOP_tmp_nor_151_itm
      AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_1518_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_61_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_60_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_59_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_58_itm AND and_dcpl_109);
  COMP_LOOP_or_3_nl <= (COMP_LOOP_COMP_LOOP_and_1370_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_760_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_1518_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_61_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_60_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_59_itm
      AND and_dcpl_109);
  COMP_LOOP_or_4_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(2)) AND COMP_LOOP_tmp_nor_153_itm
      AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_761_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_760_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_1518_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_61_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_60_itm AND and_dcpl_109);
  COMP_LOOP_or_5_nl <= (COMP_LOOP_COMP_LOOP_and_1577_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_509_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_761_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_760_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_1518_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_61_itm
      AND and_dcpl_109);
  COMP_LOOP_or_6_nl <= (COMP_LOOP_COMP_LOOP_and_1584_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_510_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_509_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_761_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_760_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_1518_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_109);
  COMP_LOOP_or_7_nl <= (COMP_LOOP_COMP_LOOP_and_1831_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_258_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_510_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_509_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_761_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_760_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_1518_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_109);
  COMP_LOOP_or_8_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(3)) AND COMP_LOOP_tmp_nor_157_itm
      AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_258_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_510_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_509_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_761_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_760_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_1518_itm AND and_dcpl_109);
  COMP_LOOP_or_9_nl <= (COMP_LOOP_COMP_LOOP_and_1874_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_260_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_258_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_510_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_509_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_761_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_and_760_itm AND and_dcpl_109);
  COMP_LOOP_or_10_nl <= (COMP_LOOP_COMP_LOOP_and_583_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_261_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_260_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_258_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_510_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_509_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_and_761_itm AND and_dcpl_109);
  COMP_LOOP_or_11_nl <= (COMP_LOOP_COMP_LOOP_and_73_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_262_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_261_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_260_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_258_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_510_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_and_509_itm AND and_dcpl_109);
  COMP_LOOP_or_12_nl <= (COMP_LOOP_COMP_LOOP_and_74_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_262_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_261_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_260_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_258_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_and_510_itm AND and_dcpl_109);
  COMP_LOOP_or_13_nl <= (COMP_LOOP_COMP_LOOP_and_75_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_264_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_262_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_261_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_260_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_258_itm
      AND and_dcpl_109);
  COMP_LOOP_or_14_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_264_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_262_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_261_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_260_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_109);
  COMP_LOOP_or_15_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_264_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_262_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_261_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_260_itm AND and_dcpl_109);
  COMP_LOOP_or_16_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(4)) AND COMP_LOOP_tmp_nor_165_itm
      AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_264_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_262_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_261_itm AND and_dcpl_109);
  COMP_LOOP_or_17_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_268_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_264_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_262_itm AND and_dcpl_109);
  COMP_LOOP_or_18_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_522_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_268_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_264_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_109);
  COMP_LOOP_or_19_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_270_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_522_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_268_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_264_itm AND and_dcpl_109);
  COMP_LOOP_or_20_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_18_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_270_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_522_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_268_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_109);
  COMP_LOOP_or_21_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_272_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_18_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_270_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_522_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_268_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_109);
  COMP_LOOP_or_22_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_20_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_272_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_18_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_270_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_522_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_268_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_109);
  COMP_LOOP_or_23_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_21_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_20_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_272_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_18_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_270_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_522_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_268_itm AND and_dcpl_109);
  COMP_LOOP_or_24_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_22_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_21_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_20_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_272_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_18_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_270_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_522_itm AND and_dcpl_109);
  COMP_LOOP_or_25_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_23_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_22_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_21_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_20_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_272_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_18_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_270_itm AND and_dcpl_109);
  COMP_LOOP_or_26_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_24_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_23_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_22_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_21_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_20_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_272_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_18_itm AND and_dcpl_109);
  COMP_LOOP_or_27_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_25_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_24_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_23_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_22_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_21_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_20_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_272_itm AND and_dcpl_109);
  COMP_LOOP_or_28_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_26_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_25_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_24_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_23_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_22_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_21_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_20_itm AND and_dcpl_109);
  COMP_LOOP_or_29_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_27_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_26_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_25_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_24_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_23_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_22_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_21_itm AND and_dcpl_109);
  COMP_LOOP_or_30_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_28_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_27_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_26_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_25_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_24_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_23_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_22_itm AND and_dcpl_109);
  COMP_LOOP_or_31_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_29_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_28_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_27_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_26_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_25_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_24_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_23_itm AND and_dcpl_109);
  COMP_LOOP_or_32_nl <= ((COMP_LOOP_acc_10_cse_10_1_1_sva(5)) AND COMP_LOOP_tmp_nor_180_itm
      AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_29_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_28_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_27_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_26_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_25_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_24_itm AND and_dcpl_109);
  COMP_LOOP_or_33_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_284_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_29_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_28_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_27_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_26_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_25_itm AND and_dcpl_109);
  COMP_LOOP_or_34_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_285_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_284_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_29_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_28_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_27_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_26_itm AND and_dcpl_109);
  COMP_LOOP_or_35_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_286_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_285_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_284_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_29_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_28_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_27_itm AND and_dcpl_109);
  COMP_LOOP_or_36_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_34_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_286_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_285_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_284_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_30_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_29_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_28_itm AND and_dcpl_109);
  COMP_LOOP_or_37_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm AND and_dcpl_77)
      OR (COMP_LOOP_COMP_LOOP_and_288_itm AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_34_itm
      AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_286_itm AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_285_itm
      AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_284_itm AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_30_itm
      AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_29_itm AND and_dcpl_109);
  COMP_LOOP_or_38_nl <= (COMP_LOOP_COMP_LOOP_and_100_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_36_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_288_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_34_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_286_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_285_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_284_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_and_30_itm AND and_dcpl_109);
  COMP_LOOP_or_39_nl <= (COMP_LOOP_COMP_LOOP_and_101_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_37_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_36_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_288_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_34_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_286_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_285_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_and_284_itm AND and_dcpl_109);
  COMP_LOOP_or_40_nl <= (COMP_LOOP_COMP_LOOP_and_102_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_38_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_37_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_36_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_288_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_34_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_286_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_and_285_itm AND and_dcpl_109);
  COMP_LOOP_or_41_nl <= (COMP_LOOP_COMP_LOOP_and_103_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_39_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_38_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_37_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_36_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_288_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_34_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_286_itm
      AND and_dcpl_109);
  COMP_LOOP_or_42_nl <= (COMP_LOOP_COMP_LOOP_and_104_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_40_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_39_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_38_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_37_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_36_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_288_itm AND and_dcpl_106) OR
      (COMP_LOOP_COMP_LOOP_and_34_itm AND and_dcpl_109);
  COMP_LOOP_or_43_nl <= (COMP_LOOP_COMP_LOOP_and_105_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_41_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_40_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_39_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_38_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_37_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_36_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_288_itm
      AND and_dcpl_109);
  COMP_LOOP_or_44_nl <= (COMP_LOOP_COMP_LOOP_and_106_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_42_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_41_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_40_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_39_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_38_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_37_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_36_itm
      AND and_dcpl_109);
  COMP_LOOP_or_45_nl <= (COMP_LOOP_COMP_LOOP_and_107_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_43_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_42_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_41_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_40_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_39_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_38_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_37_itm
      AND and_dcpl_109);
  COMP_LOOP_or_46_nl <= (COMP_LOOP_COMP_LOOP_and_108_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_44_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_43_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_42_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_41_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_40_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_39_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_38_itm
      AND and_dcpl_109);
  COMP_LOOP_or_47_nl <= (COMP_LOOP_COMP_LOOP_and_109_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_45_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_44_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_43_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_42_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_41_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_40_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_39_itm
      AND and_dcpl_109);
  COMP_LOOP_or_48_nl <= (COMP_LOOP_COMP_LOOP_and_110_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_46_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_45_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_44_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_43_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_42_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_41_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_40_itm
      AND and_dcpl_109);
  COMP_LOOP_or_49_nl <= (COMP_LOOP_COMP_LOOP_and_1104_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_47_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_46_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_45_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_44_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_43_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_42_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_41_itm
      AND and_dcpl_109);
  COMP_LOOP_or_50_nl <= (COMP_LOOP_COMP_LOOP_and_1106_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_48_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_47_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_46_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_45_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_44_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_43_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_42_itm
      AND and_dcpl_109);
  COMP_LOOP_or_51_nl <= (COMP_LOOP_COMP_LOOP_and_1110_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_49_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_48_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_47_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_46_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_45_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_44_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_43_itm
      AND and_dcpl_109);
  COMP_LOOP_or_52_nl <= (COMP_LOOP_COMP_LOOP_and_1118_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_50_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_49_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_48_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_47_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_46_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_45_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_44_itm
      AND and_dcpl_109);
  COMP_LOOP_or_53_nl <= (COMP_LOOP_COMP_LOOP_and_115_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_51_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_50_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_49_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_48_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_47_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_46_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_45_itm
      AND and_dcpl_109);
  COMP_LOOP_or_54_nl <= (COMP_LOOP_COMP_LOOP_and_116_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_52_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_51_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_50_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_49_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_48_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_47_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_46_itm
      AND and_dcpl_109);
  COMP_LOOP_or_55_nl <= (COMP_LOOP_COMP_LOOP_and_117_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_53_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_52_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_51_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_50_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_49_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_48_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_47_itm
      AND and_dcpl_109);
  COMP_LOOP_or_56_nl <= (COMP_LOOP_COMP_LOOP_and_118_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_54_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_53_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_52_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_51_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_50_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_49_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_48_itm
      AND and_dcpl_109);
  COMP_LOOP_or_57_nl <= (COMP_LOOP_COMP_LOOP_and_119_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_55_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_54_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_53_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_52_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_51_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_50_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_49_itm
      AND and_dcpl_109);
  COMP_LOOP_or_58_nl <= (COMP_LOOP_COMP_LOOP_and_120_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_56_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_55_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_54_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_53_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_52_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_51_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_50_itm
      AND and_dcpl_109);
  COMP_LOOP_or_59_nl <= (COMP_LOOP_COMP_LOOP_and_121_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_57_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_56_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_55_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_54_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_53_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_52_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_51_itm
      AND and_dcpl_109);
  COMP_LOOP_or_60_nl <= (COMP_LOOP_COMP_LOOP_and_122_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_58_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_57_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_56_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_55_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_54_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_53_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_52_itm
      AND and_dcpl_109);
  COMP_LOOP_or_61_nl <= (COMP_LOOP_COMP_LOOP_and_123_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_59_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_58_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_57_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_56_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_55_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_54_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_53_itm
      AND and_dcpl_109);
  COMP_LOOP_or_62_nl <= (COMP_LOOP_COMP_LOOP_and_124_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_60_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_59_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_58_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_57_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_56_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_55_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_54_itm
      AND and_dcpl_109);
  COMP_LOOP_or_63_nl <= (COMP_LOOP_COMP_LOOP_and_125_itm AND and_dcpl_77) OR (COMP_LOOP_COMP_LOOP_and_61_itm
      AND and_dcpl_86) OR (COMP_LOOP_COMP_LOOP_and_60_itm AND and_dcpl_90) OR (COMP_LOOP_COMP_LOOP_and_59_itm
      AND and_dcpl_95) OR (COMP_LOOP_COMP_LOOP_and_58_itm AND and_dcpl_99) OR (COMP_LOOP_COMP_LOOP_and_57_itm
      AND and_dcpl_104) OR (COMP_LOOP_COMP_LOOP_and_56_itm AND and_dcpl_106) OR (COMP_LOOP_COMP_LOOP_and_55_itm
      AND and_dcpl_109);
  COMP_LOOP_tmp_and_249_nl <= COMP_LOOP_COMP_LOOP_and_119_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(0)) AND COMP_LOOP_tmp_nor_153_itm
      AND (NOT and_474_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(1)) AND COMP_LOOP_tmp_nor_165_itm
      AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_250_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(2)) AND
      COMP_LOOP_tmp_nor_180_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_251_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_252_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_253_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(3)) AND
      COMP_LOOP_tmp_nor_10_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_254_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_255_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_256_nl <= COMP_LOOP_COMP_LOOP_and_102_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_257_nl <= COMP_LOOP_COMP_LOOP_and_106_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_258_nl <= COMP_LOOP_COMP_LOOP_and_107_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_259_nl <= COMP_LOOP_COMP_LOOP_and_108_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_260_nl <= COMP_LOOP_COMP_LOOP_and_109_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_22_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(4)) AND
      COMP_LOOP_tmp_nor_151_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_261_nl <= COMP_LOOP_COMP_LOOP_and_110_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_262_nl <= COMP_LOOP_COMP_LOOP_and_1104_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_263_nl <= COMP_LOOP_COMP_LOOP_and_1106_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_264_nl <= COMP_LOOP_COMP_LOOP_and_1118_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_265_nl <= COMP_LOOP_COMP_LOOP_and_115_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_266_nl <= COMP_LOOP_COMP_LOOP_and_116_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_267_nl <= COMP_LOOP_COMP_LOOP_and_117_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_268_nl <= COMP_LOOP_COMP_LOOP_and_118_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_269_nl <= COMP_LOOP_COMP_LOOP_and_120_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_270_nl <= COMP_LOOP_COMP_LOOP_and_121_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_271_nl <= COMP_LOOP_COMP_LOOP_and_122_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_272_nl <= COMP_LOOP_COMP_LOOP_and_123_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_273_nl <= COMP_LOOP_COMP_LOOP_and_124_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_274_nl <= COMP_LOOP_COMP_LOOP_and_125_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_275_nl <= COMP_LOOP_COMP_LOOP_and_1370_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(5)) AND
      COMP_LOOP_tmp_nor_157_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_276_nl <= COMP_LOOP_COMP_LOOP_and_1831_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_277_nl <= COMP_LOOP_COMP_LOOP_and_1874_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_278_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_279_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_280_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_281_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_282_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_283_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_284_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_285_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_286_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_287_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_288_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_289_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_290_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_291_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_292_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_293_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_294_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_295_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_296_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_297_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_298_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_299_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_300_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_301_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_302_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_303_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_304_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_305_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_306_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm AND (NOT and_474_tmp);
  COMP_LOOP_tmp_and_222_nl <= COMP_LOOP_COMP_LOOP_and_1874_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_70_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_4_0(0))
      AND COMP_LOOP_tmp_nor_206_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_71_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_4_0(1))
      AND COMP_LOOP_tmp_nor_207_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_223_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_73_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_4_0(2))
      AND COMP_LOOP_tmp_nor_209_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_224_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_225_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_226_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_77_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_4_0(3))
      AND COMP_LOOP_tmp_nor_213_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_227_nl <= COMP_LOOP_COMP_LOOP_and_102_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_228_nl <= COMP_LOOP_COMP_LOOP_and_106_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_229_nl <= COMP_LOOP_COMP_LOOP_and_107_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_230_nl <= COMP_LOOP_COMP_LOOP_and_108_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_231_nl <= COMP_LOOP_COMP_LOOP_and_109_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_232_nl <= COMP_LOOP_COMP_LOOP_and_110_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_233_nl <= COMP_LOOP_COMP_LOOP_and_1104_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_nl <= (COMP_LOOP_3_tmp_mul_idiv_sva_4_0(4))
      AND COMP_LOOP_tmp_nor_220_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_234_nl <= COMP_LOOP_COMP_LOOP_and_1106_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_235_nl <= COMP_LOOP_COMP_LOOP_and_1118_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_236_nl <= COMP_LOOP_COMP_LOOP_and_115_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_237_nl <= COMP_LOOP_COMP_LOOP_and_116_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_238_nl <= COMP_LOOP_COMP_LOOP_and_117_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_239_nl <= COMP_LOOP_COMP_LOOP_and_118_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_240_nl <= COMP_LOOP_COMP_LOOP_and_120_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_241_nl <= COMP_LOOP_COMP_LOOP_and_121_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_242_nl <= COMP_LOOP_COMP_LOOP_and_122_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_243_nl <= COMP_LOOP_COMP_LOOP_and_123_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_244_nl <= COMP_LOOP_COMP_LOOP_and_124_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_245_nl <= COMP_LOOP_COMP_LOOP_and_125_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_246_nl <= COMP_LOOP_COMP_LOOP_and_1370_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_247_nl <= COMP_LOOP_COMP_LOOP_and_1831_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_248_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND (NOT nor_1579_tmp);
  COMP_LOOP_tmp_and_164_nl <= COMP_LOOP_COMP_LOOP_and_119_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(0)) AND
      COMP_LOOP_tmp_nor_151_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_102_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(1)) AND
      COMP_LOOP_tmp_nor_153_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_165_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(2)) AND
      COMP_LOOP_tmp_nor_157_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_166_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_167_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_168_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(3)) AND
      COMP_LOOP_tmp_nor_165_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_169_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_170_nl <= COMP_LOOP_COMP_LOOP_and_102_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_171_nl <= COMP_LOOP_COMP_LOOP_and_106_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_172_nl <= COMP_LOOP_COMP_LOOP_and_107_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_173_nl <= COMP_LOOP_COMP_LOOP_and_108_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_174_nl <= COMP_LOOP_COMP_LOOP_and_109_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_175_nl <= COMP_LOOP_COMP_LOOP_and_110_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(4)) AND
      COMP_LOOP_tmp_nor_180_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_176_nl <= COMP_LOOP_COMP_LOOP_and_1104_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_177_nl <= COMP_LOOP_COMP_LOOP_and_1106_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_178_nl <= COMP_LOOP_COMP_LOOP_and_1118_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_179_nl <= COMP_LOOP_COMP_LOOP_and_115_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_180_nl <= COMP_LOOP_COMP_LOOP_and_116_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_181_nl <= COMP_LOOP_COMP_LOOP_and_117_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_182_nl <= COMP_LOOP_COMP_LOOP_and_118_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_183_nl <= COMP_LOOP_COMP_LOOP_and_120_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_184_nl <= COMP_LOOP_COMP_LOOP_and_121_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_185_nl <= COMP_LOOP_COMP_LOOP_and_122_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_186_nl <= COMP_LOOP_COMP_LOOP_and_123_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_187_nl <= COMP_LOOP_COMP_LOOP_and_124_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_188_nl <= COMP_LOOP_COMP_LOOP_and_125_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_189_nl <= COMP_LOOP_COMP_LOOP_and_1370_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_190_nl <= COMP_LOOP_COMP_LOOP_and_1831_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(5)) AND
      COMP_LOOP_tmp_nor_10_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_191_nl <= COMP_LOOP_COMP_LOOP_and_1874_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_192_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_193_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_194_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_195_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_196_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_197_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_198_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_199_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_200_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_201_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_202_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_203_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_204_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_205_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_206_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_207_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_208_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_209_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_210_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_211_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_212_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_213_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_214_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_215_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_216_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_217_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_218_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_219_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_220_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_221_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm AND (NOT and_476_tmp);
  COMP_LOOP_tmp_and_152_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_164_nl <= (COMP_LOOP_5_tmp_mul_idiv_sva(0)) AND
      COMP_LOOP_tmp_nor_140_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_165_nl <= (COMP_LOOP_5_tmp_mul_idiv_sva(1)) AND
      COMP_LOOP_tmp_nor_141_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_153_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_166_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_167_nl <= (COMP_LOOP_5_tmp_mul_idiv_sva(2)) AND
      COMP_LOOP_tmp_nor_143_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_154_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_168_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_155_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_169_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_156_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_170_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_171_nl <= (COMP_LOOP_5_tmp_mul_idiv_sva(3)) AND
      COMP_LOOP_tmp_nor_146_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_157_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_172_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_158_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_173_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_159_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_160_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_175_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_161_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_176_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_162_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_177_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_163_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_178_itm AND (NOT nor_tmp_396);
  COMP_LOOP_tmp_and_89_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_90_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_274_rgt AND and_478_m1c;
  COMP_LOOP_tmp_and_91_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_92_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_276_rgt AND and_478_m1c;
  COMP_LOOP_tmp_and_93_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_94_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_95_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_96_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_280_rgt AND and_478_m1c;
  COMP_LOOP_tmp_and_97_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_98_nl <= COMP_LOOP_COMP_LOOP_and_102_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_99_nl <= COMP_LOOP_COMP_LOOP_and_106_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_100_nl <= COMP_LOOP_COMP_LOOP_and_107_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_101_nl <= COMP_LOOP_COMP_LOOP_and_108_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_102_nl <= COMP_LOOP_COMP_LOOP_and_109_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_103_nl <= COMP_LOOP_COMP_LOOP_and_110_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_104_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_288_rgt AND and_478_m1c;
  COMP_LOOP_tmp_and_105_nl <= COMP_LOOP_COMP_LOOP_and_1104_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_106_nl <= COMP_LOOP_COMP_LOOP_and_1106_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_107_nl <= COMP_LOOP_COMP_LOOP_and_1118_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_108_nl <= COMP_LOOP_COMP_LOOP_and_115_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_109_nl <= COMP_LOOP_COMP_LOOP_and_116_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_110_nl <= COMP_LOOP_COMP_LOOP_and_117_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_111_nl <= COMP_LOOP_COMP_LOOP_and_118_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_112_nl <= COMP_LOOP_COMP_LOOP_and_120_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_113_nl <= COMP_LOOP_COMP_LOOP_and_121_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_114_nl <= COMP_LOOP_COMP_LOOP_and_122_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_115_nl <= COMP_LOOP_COMP_LOOP_and_123_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_116_nl <= COMP_LOOP_COMP_LOOP_and_124_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_117_nl <= COMP_LOOP_COMP_LOOP_and_125_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_118_nl <= COMP_LOOP_COMP_LOOP_and_1370_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_119_nl <= COMP_LOOP_COMP_LOOP_and_1831_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_120_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_304_rgt AND and_478_m1c;
  COMP_LOOP_tmp_and_121_nl <= COMP_LOOP_COMP_LOOP_and_1874_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_122_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_123_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_124_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_125_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_126_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_127_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_128_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_129_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_130_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_131_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_132_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_133_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_134_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_135_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_136_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_137_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_138_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_139_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_140_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_141_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_142_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_143_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_144_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_145_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_146_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_147_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_148_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_149_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_150_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm AND and_478_m1c;
  COMP_LOOP_tmp_and_151_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm AND and_478_m1c;
  mux_3350_nl <= MUX_s_1_2_2(not_tmp_88, nor_tmp_391, fsm_output(6));
  mux_3351_nl <= MUX_s_1_2_2(mux_3350_nl, mux_tmp_3280, fsm_output(2));
  mux_3348_nl <= MUX_s_1_2_2(not_tmp_868, nor_tmp_391, fsm_output(6));
  mux_3349_nl <= MUX_s_1_2_2(mux_3348_nl, mux_tmp_3280, fsm_output(2));
  mux_3352_nl <= MUX_s_1_2_2(mux_3351_nl, mux_3349_nl, fsm_output(1));
  mux_3353_nl <= MUX_s_1_2_2(mux_3352_nl, and_705_cse, fsm_output(5));
  COMP_LOOP_tmp_and_31_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_179_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(0)) AND
      COMP_LOOP_tmp_nor_10_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_180_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(1)) AND
      COMP_LOOP_tmp_nor_151_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_32_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_182_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(2)) AND
      COMP_LOOP_tmp_nor_153_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_33_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_34_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_35_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_186_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(3)) AND
      COMP_LOOP_tmp_nor_157_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_36_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_37_nl <= COMP_LOOP_COMP_LOOP_and_102_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_38_nl <= COMP_LOOP_COMP_LOOP_and_106_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_39_nl <= COMP_LOOP_COMP_LOOP_and_107_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_40_nl <= COMP_LOOP_COMP_LOOP_and_108_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_41_nl <= COMP_LOOP_COMP_LOOP_and_109_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_42_nl <= COMP_LOOP_COMP_LOOP_and_110_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_194_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(4)) AND
      COMP_LOOP_tmp_nor_165_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_43_nl <= COMP_LOOP_COMP_LOOP_and_1104_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_44_nl <= COMP_LOOP_COMP_LOOP_and_1106_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_45_nl <= COMP_LOOP_COMP_LOOP_and_1118_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_46_nl <= COMP_LOOP_COMP_LOOP_and_115_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_47_nl <= COMP_LOOP_COMP_LOOP_and_116_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_48_nl <= COMP_LOOP_COMP_LOOP_and_117_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_49_nl <= COMP_LOOP_COMP_LOOP_and_118_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_50_nl <= COMP_LOOP_COMP_LOOP_and_120_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_51_nl <= COMP_LOOP_COMP_LOOP_and_121_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_52_nl <= COMP_LOOP_COMP_LOOP_and_122_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_53_nl <= COMP_LOOP_COMP_LOOP_and_123_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_54_nl <= COMP_LOOP_COMP_LOOP_and_124_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_55_nl <= COMP_LOOP_COMP_LOOP_and_125_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_56_nl <= COMP_LOOP_COMP_LOOP_and_1370_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_57_nl <= COMP_LOOP_COMP_LOOP_and_1831_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_210_nl <= (COMP_LOOP_2_tmp_mul_idiv_sva(5)) AND
      COMP_LOOP_tmp_nor_180_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_58_nl <= COMP_LOOP_COMP_LOOP_and_1874_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_59_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_60_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_61_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_62_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_63_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_64_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_65_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_66_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_67_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_68_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_69_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_70_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_71_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_72_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_73_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_74_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_75_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_76_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_77_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_78_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_79_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_80_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_81_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_82_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_83_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_84_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_85_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_86_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_87_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_88_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm AND mux_3360_tmp;
  COMP_LOOP_tmp_and_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_1_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_243_rgt AND and_dcpl_265;
  COMP_LOOP_tmp_and_2_nl <= COMP_LOOP_COMP_LOOP_and_119_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_3_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_245_rgt AND and_dcpl_265;
  COMP_LOOP_tmp_and_4_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_5_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_6_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_7_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_249_rgt AND and_dcpl_265;
  COMP_LOOP_tmp_and_8_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_9_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_10_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_11_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_12_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_13_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_14_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_15_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_257_rgt AND and_dcpl_265;
  COMP_LOOP_tmp_and_16_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_17_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_18_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_19_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_20_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_21_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_22_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_23_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_24_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_25_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_26_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_27_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_28_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_29_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm AND and_dcpl_265;
  COMP_LOOP_tmp_and_30_nl <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm AND and_dcpl_265;
  mux_3362_nl <= MUX_s_1_2_2(not_tmp_88, (fsm_output(7)), fsm_output(6));
  mux_3363_nl <= MUX_s_1_2_2(mux_3362_nl, mux_tmp_3100, or_359_cse);
  mux_3361_nl <= MUX_s_1_2_2(nor_tmp_391, (fsm_output(7)), fsm_output(6));
  mux_3364_nl <= MUX_s_1_2_2(mux_3363_nl, mux_3361_nl, fsm_output(5));
  and_1047_nl <= and_dcpl_58 AND (NOT (fsm_output(3))) AND (fsm_output(6)) AND (fsm_output(2))
      AND (NOT (fsm_output(1))) AND (fsm_output(7)) AND (fsm_output(5));
  COMP_LOOP_mux_721_nl <= MUX_v_7_2_2(COMP_LOOP_k_10_3_sva_6_0, (STD_LOGIC_VECTOR'(
      "001") & (NOT z_out_4)), and_1047_nl);
  z_out_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_721_nl),
      8) + UNSIGNED'( "00000001"), 8));
  COMP_LOOP_mux_722_nl <= MUX_v_11_2_2(('1' & (NOT (STAGE_LOOP_lshift_psp_sva(10
      DOWNTO 1)))), STAGE_LOOP_lshift_psp_sva, and_dcpl_488);
  COMP_LOOP_COMP_LOOP_nand_1_nl <= NOT(and_dcpl_488 AND (NOT(and_dcpl_58 AND nor_1715_cse
      AND and_dcpl_477 AND nor_1716_cse)));
  COMP_LOOP_mux_723_nl <= MUX_v_10_2_2((COMP_LOOP_k_10_3_sva_6_0 & STD_LOGIC_VECTOR'(
      "001")), VEC_LOOP_j_10_0_sva_9_0, and_dcpl_488);
  acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_722_nl & COMP_LOOP_COMP_LOOP_nand_1_nl)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_723_nl & '1'), 11), 12),
      12));
  z_out_3 <= acc_1_nl(11 DOWNTO 1);
  STAGE_LOOP_mux_4_nl <= MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, (NOT STAGE_LOOP_i_3_0_sva),
      and_dcpl_501);
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_mux_4_nl) + UNSIGNED('1'
      & (NOT and_dcpl_501) & STD_LOGIC_VECTOR'( "11")), 4));
  COMP_LOOP_mux_724_cse <= MUX_v_64_2_2(z_out_9, COMP_LOOP_1_acc_8_itm, COMP_LOOP_or_65_itm);
  COMP_LOOP_tmp_nor_300_cse <= NOT(and_dcpl_574 OR and_dcpl_589 OR and_dcpl_590);
  COMP_LOOP_tmp_mux_64_nl <= MUX_s_1_2_2((z_out_1(9)), (COMP_LOOP_2_tmp_lshift_ncse_sva(9)),
      COMP_LOOP_tmp_or_54_ssc);
  COMP_LOOP_tmp_COMP_LOOP_tmp_and_337_nl <= COMP_LOOP_tmp_mux_64_nl AND COMP_LOOP_tmp_nor_300_cse;
  COMP_LOOP_tmp_or_88_nl <= and_dcpl_577 OR and_dcpl_589;
  COMP_LOOP_tmp_mux1h_146_nl <= MUX1HOT_v_9_4_2(('0' & (z_out(7 DOWNTO 0))), (z_out_1(8
      DOWNTO 0)), (COMP_LOOP_2_tmp_lshift_ncse_sva(8 DOWNTO 0)), COMP_LOOP_3_tmp_lshift_ncse_sva,
      STD_LOGIC_VECTOR'( and_dcpl_574 & COMP_LOOP_tmp_or_88_nl & COMP_LOOP_tmp_or_54_ssc
      & and_dcpl_590));
  COMP_LOOP_tmp_and_312_nl <= (COMP_LOOP_k_10_3_sva_6_0(6)) AND COMP_LOOP_tmp_nor_300_cse;
  COMP_LOOP_tmp_or_89_nl <= and_dcpl_577 OR and_dcpl_580 OR and_dcpl_583 OR and_dcpl_588;
  COMP_LOOP_tmp_mux1h_147_nl <= MUX1HOT_v_6_3_2(('0' & (COMP_LOOP_k_10_3_sva_6_0(6
      DOWNTO 2))), (COMP_LOOP_k_10_3_sva_6_0(5 DOWNTO 0)), (COMP_LOOP_k_10_3_sva_6_0(6
      DOWNTO 1)), STD_LOGIC_VECTOR'( and_dcpl_574 & COMP_LOOP_tmp_or_89_nl & COMP_LOOP_tmp_or_83_itm));
  COMP_LOOP_tmp_COMP_LOOP_tmp_mux_17_nl <= MUX_s_1_2_2((COMP_LOOP_k_10_3_sva_6_0(1)),
      (COMP_LOOP_k_10_3_sva_6_0(0)), COMP_LOOP_tmp_or_83_itm);
  COMP_LOOP_tmp_or_90_nl <= (COMP_LOOP_tmp_COMP_LOOP_tmp_mux_17_nl AND (NOT(and_dcpl_577
      OR and_dcpl_580))) OR and_dcpl_583 OR and_dcpl_588;
  COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl <= ((COMP_LOOP_k_10_3_sva_6_0(0)) AND (NOT(and_dcpl_577
      OR and_dcpl_583 OR and_dcpl_589))) OR and_dcpl_580 OR and_dcpl_588 OR and_dcpl_590;
  z_out_7 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(COMP_LOOP_tmp_COMP_LOOP_tmp_and_337_nl
      & COMP_LOOP_tmp_mux1h_146_nl) * UNSIGNED(COMP_LOOP_tmp_and_312_nl & COMP_LOOP_tmp_mux1h_147_nl
      & COMP_LOOP_tmp_or_90_nl & COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl & '1')), 10));
  and_1048_nl <= and_dcpl_573 AND CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"))
      AND nor_1716_cse;
  COMP_LOOP_tmp_mux1h_148_nl <= MUX1HOT_v_64_9_2((STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000")
      & (z_out_1(6 DOWNTO 0))), COMP_LOOP_tmp_mux1h_itm, COMP_LOOP_tmp_mux1h_1_itm,
      COMP_LOOP_tmp_mux1h_2_itm, COMP_LOOP_tmp_mux1h_3_itm, COMP_LOOP_tmp_mux1h_4_itm,
      COMP_LOOP_tmp_mux1h_5_itm, COMP_LOOP_tmp_mux1h_6_itm, tmp_21_sva_1, STD_LOGIC_VECTOR'(
      and_1048_nl & and_dcpl_602 & and_dcpl_608 & and_dcpl_611 & and_dcpl_614 & and_dcpl_617
      & and_dcpl_620 & and_dcpl_623 & and_dcpl_625));
  COMP_LOOP_tmp_or_91_nl <= and_dcpl_602 OR and_dcpl_608 OR and_dcpl_611 OR and_dcpl_614
      OR and_dcpl_617 OR and_dcpl_620 OR and_dcpl_623 OR and_dcpl_625;
  COMP_LOOP_tmp_mux_65_nl <= MUX_v_64_2_2((STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000")
      & COMP_LOOP_k_10_3_sva_6_0), COMP_LOOP_1_modulo_dev_cmp_return_rsc_z, COMP_LOOP_tmp_or_91_nl);
  z_out_8 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(COMP_LOOP_tmp_mux1h_148_nl)
      * UNSIGNED(COMP_LOOP_tmp_mux_65_nl)), 64));
  COMP_LOOP_mux1h_1267_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_nor_itm, COMP_LOOP_COMP_LOOP_nor_5_itm,
      COMP_LOOP_COMP_LOOP_nor_9_itm, COMP_LOOP_COMP_LOOP_nor_13_itm, COMP_LOOP_COMP_LOOP_nor_17_itm,
      COMP_LOOP_COMP_LOOP_nor_21_itm, COMP_LOOP_COMP_LOOP_nor_25_itm, COMP_LOOP_COMP_LOOP_nor_29_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_COMP_LOOP_and_1890_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(0)) AND COMP_LOOP_nor_281_itm;
  COMP_LOOP_COMP_LOOP_and_1891_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(0)) AND COMP_LOOP_nor_505_itm;
  COMP_LOOP_COMP_LOOP_and_1892_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(0)) AND COMP_LOOP_nor_729_itm;
  COMP_LOOP_COMP_LOOP_and_1893_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(0)) AND COMP_LOOP_nor_953_itm;
  COMP_LOOP_COMP_LOOP_and_1894_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(0)) AND COMP_LOOP_nor_1177_itm;
  COMP_LOOP_COMP_LOOP_and_1895_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(0)) AND COMP_LOOP_nor_1401_itm;
  COMP_LOOP_COMP_LOOP_and_1896_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(0)) AND COMP_LOOP_nor_1625_itm;
  COMP_LOOP_mux1h_1268_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_1518_itm, COMP_LOOP_COMP_LOOP_and_1890_nl,
      COMP_LOOP_COMP_LOOP_and_1891_nl, COMP_LOOP_COMP_LOOP_and_1892_nl, COMP_LOOP_COMP_LOOP_and_1893_nl,
      COMP_LOOP_COMP_LOOP_and_1894_nl, COMP_LOOP_COMP_LOOP_and_1895_nl, COMP_LOOP_COMP_LOOP_and_1896_nl,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_COMP_LOOP_and_1897_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(1)) AND COMP_LOOP_nor_282_itm;
  COMP_LOOP_COMP_LOOP_and_1898_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(1)) AND COMP_LOOP_nor_506_itm;
  COMP_LOOP_COMP_LOOP_and_1899_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(1)) AND COMP_LOOP_nor_730_itm;
  COMP_LOOP_COMP_LOOP_and_1900_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(1)) AND COMP_LOOP_nor_954_itm;
  COMP_LOOP_COMP_LOOP_and_1901_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(1)) AND COMP_LOOP_nor_1178_itm;
  COMP_LOOP_COMP_LOOP_and_1902_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(1)) AND COMP_LOOP_nor_1402_itm;
  COMP_LOOP_COMP_LOOP_and_1903_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(1)) AND COMP_LOOP_nor_1626_itm;
  COMP_LOOP_mux1h_1269_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_760_itm, COMP_LOOP_COMP_LOOP_and_1897_nl,
      COMP_LOOP_COMP_LOOP_and_1898_nl, COMP_LOOP_COMP_LOOP_and_1899_nl, COMP_LOOP_COMP_LOOP_and_1900_nl,
      COMP_LOOP_COMP_LOOP_and_1901_nl, COMP_LOOP_COMP_LOOP_and_1902_nl, COMP_LOOP_COMP_LOOP_and_1903_nl,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1270_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_761_itm, COMP_LOOP_COMP_LOOP_and_1594_itm,
      COMP_LOOP_COMP_LOOP_and_569_itm, COMP_LOOP_COMP_LOOP_and_821_itm, COMP_LOOP_COMP_LOOP_and_100_itm,
      COMP_LOOP_COMP_LOOP_and_1325_itm, COMP_LOOP_COMP_LOOP_and_1577_itm, COMP_LOOP_COMP_LOOP_and_1829_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_COMP_LOOP_and_1904_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(2)) AND COMP_LOOP_nor_284_itm;
  COMP_LOOP_COMP_LOOP_and_1905_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(2)) AND COMP_LOOP_nor_508_itm;
  COMP_LOOP_COMP_LOOP_and_1906_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(2)) AND COMP_LOOP_nor_732_itm;
  COMP_LOOP_COMP_LOOP_and_1907_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(2)) AND COMP_LOOP_nor_956_itm;
  COMP_LOOP_COMP_LOOP_and_1908_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(2)) AND COMP_LOOP_nor_1180_itm;
  COMP_LOOP_COMP_LOOP_and_1909_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(2)) AND COMP_LOOP_nor_1404_itm;
  COMP_LOOP_COMP_LOOP_and_1910_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(2)) AND COMP_LOOP_nor_1628_itm;
  COMP_LOOP_mux1h_1271_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_509_itm, COMP_LOOP_COMP_LOOP_and_1904_nl,
      COMP_LOOP_COMP_LOOP_and_1905_nl, COMP_LOOP_COMP_LOOP_and_1906_nl, COMP_LOOP_COMP_LOOP_and_1907_nl,
      COMP_LOOP_COMP_LOOP_and_1908_nl, COMP_LOOP_COMP_LOOP_and_1909_nl, COMP_LOOP_COMP_LOOP_and_1910_nl,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1272_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_510_itm, COMP_LOOP_COMP_LOOP_and_1598_itm,
      COMP_LOOP_COMP_LOOP_and_571_itm, COMP_LOOP_COMP_LOOP_and_823_itm, COMP_LOOP_COMP_LOOP_and_101_itm,
      COMP_LOOP_COMP_LOOP_and_1327_itm, COMP_LOOP_COMP_LOOP_and_1579_itm, COMP_LOOP_COMP_LOOP_and_1831_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1273_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_258_itm, COMP_LOOP_COMP_LOOP_and_1607_itm,
      COMP_LOOP_COMP_LOOP_and_572_itm, COMP_LOOP_COMP_LOOP_and_73_itm, COMP_LOOP_COMP_LOOP_and_102_itm,
      COMP_LOOP_COMP_LOOP_and_115_itm, COMP_LOOP_COMP_LOOP_and_1580_itm, COMP_LOOP_COMP_LOOP_and_1832_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1274_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_6_itm, COMP_LOOP_COMP_LOOP_and_1610_itm,
      COMP_LOOP_COMP_LOOP_and_573_itm, COMP_LOOP_COMP_LOOP_and_825_itm, COMP_LOOP_COMP_LOOP_and_1077_itm,
      COMP_LOOP_COMP_LOOP_and_1329_itm, COMP_LOOP_COMP_LOOP_and_1581_itm, COMP_LOOP_COMP_LOOP_and_1833_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_COMP_LOOP_and_1911_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(3)) AND COMP_LOOP_nor_288_itm;
  COMP_LOOP_COMP_LOOP_and_1912_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(3)) AND COMP_LOOP_nor_512_itm;
  COMP_LOOP_COMP_LOOP_and_1913_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(3)) AND COMP_LOOP_nor_736_itm;
  COMP_LOOP_COMP_LOOP_and_1914_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(3)) AND COMP_LOOP_nor_960_itm;
  COMP_LOOP_COMP_LOOP_and_1915_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(3)) AND COMP_LOOP_nor_1184_itm;
  COMP_LOOP_COMP_LOOP_and_1916_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(3)) AND COMP_LOOP_nor_1408_itm;
  COMP_LOOP_COMP_LOOP_and_1917_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(3)) AND COMP_LOOP_nor_1632_itm;
  COMP_LOOP_mux1h_1275_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_260_itm, COMP_LOOP_COMP_LOOP_and_1911_nl,
      COMP_LOOP_COMP_LOOP_and_1912_nl, COMP_LOOP_COMP_LOOP_and_1913_nl, COMP_LOOP_COMP_LOOP_and_1914_nl,
      COMP_LOOP_COMP_LOOP_and_1915_nl, COMP_LOOP_COMP_LOOP_and_1916_nl, COMP_LOOP_COMP_LOOP_and_1917_nl,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1276_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_261_itm, COMP_LOOP_COMP_LOOP_and_100_itm,
      COMP_LOOP_COMP_LOOP_and_575_itm, COMP_LOOP_COMP_LOOP_and_827_itm, COMP_LOOP_COMP_LOOP_and_103_itm,
      COMP_LOOP_COMP_LOOP_and_116_itm, COMP_LOOP_COMP_LOOP_and_1583_itm, COMP_LOOP_COMP_LOOP_and_1835_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1277_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_262_itm, COMP_LOOP_COMP_LOOP_and_1614_itm,
      COMP_LOOP_COMP_LOOP_and_576_itm, COMP_LOOP_COMP_LOOP_and_828_itm, COMP_LOOP_COMP_LOOP_and_104_itm,
      COMP_LOOP_COMP_LOOP_and_117_itm, COMP_LOOP_COMP_LOOP_and_1584_itm, COMP_LOOP_COMP_LOOP_and_1836_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1278_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_10_itm, COMP_LOOP_COMP_LOOP_and_1622_itm,
      COMP_LOOP_COMP_LOOP_and_577_itm, COMP_LOOP_COMP_LOOP_and_829_itm, COMP_LOOP_COMP_LOOP_and_1081_itm,
      COMP_LOOP_COMP_LOOP_and_1333_itm, COMP_LOOP_COMP_LOOP_and_1585_itm, COMP_LOOP_COMP_LOOP_and_1837_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1279_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_264_itm, COMP_LOOP_COMP_LOOP_and_1832_itm,
      COMP_LOOP_COMP_LOOP_and_578_itm, COMP_LOOP_COMP_LOOP_and_830_itm, COMP_LOOP_COMP_LOOP_and_105_itm,
      COMP_LOOP_COMP_LOOP_and_118_itm, COMP_LOOP_COMP_LOOP_and_1586_itm, COMP_LOOP_COMP_LOOP_and_1838_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1280_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_12_itm, COMP_LOOP_COMP_LOOP_and_1835_itm,
      COMP_LOOP_COMP_LOOP_and_579_itm, COMP_LOOP_COMP_LOOP_and_831_itm, COMP_LOOP_COMP_LOOP_and_1083_itm,
      COMP_LOOP_COMP_LOOP_and_1335_itm, COMP_LOOP_COMP_LOOP_and_1587_itm, COMP_LOOP_COMP_LOOP_and_1839_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1281_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_13_itm, COMP_LOOP_COMP_LOOP_and_1844_itm,
      COMP_LOOP_COMP_LOOP_and_580_itm, COMP_LOOP_COMP_LOOP_and_832_itm, COMP_LOOP_COMP_LOOP_and_1084_itm,
      COMP_LOOP_COMP_LOOP_and_1336_itm, COMP_LOOP_COMP_LOOP_and_1588_itm, COMP_LOOP_COMP_LOOP_and_1840_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1282_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_14_itm, COMP_LOOP_COMP_LOOP_and_1850_itm,
      COMP_LOOP_COMP_LOOP_and_581_itm, COMP_LOOP_COMP_LOOP_and_833_itm, COMP_LOOP_COMP_LOOP_and_1085_itm,
      COMP_LOOP_COMP_LOOP_and_1337_itm, COMP_LOOP_COMP_LOOP_and_1589_itm, COMP_LOOP_COMP_LOOP_and_1841_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_COMP_LOOP_and_1918_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(4)) AND COMP_LOOP_nor_296_itm;
  COMP_LOOP_COMP_LOOP_and_1919_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(4)) AND COMP_LOOP_nor_520_itm;
  COMP_LOOP_COMP_LOOP_and_1920_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(4)) AND COMP_LOOP_nor_744_itm;
  COMP_LOOP_COMP_LOOP_and_1921_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(4)) AND COMP_LOOP_nor_968_itm;
  COMP_LOOP_COMP_LOOP_and_1922_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(4)) AND COMP_LOOP_nor_1192_itm;
  COMP_LOOP_COMP_LOOP_and_1923_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(4)) AND COMP_LOOP_nor_1416_itm;
  COMP_LOOP_COMP_LOOP_and_1924_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(4)) AND COMP_LOOP_nor_1640_itm;
  COMP_LOOP_mux1h_1283_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_268_itm, COMP_LOOP_COMP_LOOP_and_1918_nl,
      COMP_LOOP_COMP_LOOP_and_1919_nl, COMP_LOOP_COMP_LOOP_and_1920_nl, COMP_LOOP_COMP_LOOP_and_1921_nl,
      COMP_LOOP_COMP_LOOP_and_1922_nl, COMP_LOOP_COMP_LOOP_and_1923_nl, COMP_LOOP_COMP_LOOP_and_1924_nl,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1284_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_522_itm, COMP_LOOP_COMP_LOOP_and_1862_itm,
      COMP_LOOP_COMP_LOOP_and_583_itm, COMP_LOOP_COMP_LOOP_and_835_itm, COMP_LOOP_COMP_LOOP_and_106_itm,
      COMP_LOOP_COMP_LOOP_and_119_itm, COMP_LOOP_COMP_LOOP_and_1591_itm, COMP_LOOP_COMP_LOOP_and_1843_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1285_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_270_itm, COMP_LOOP_COMP_LOOP_and_1866_itm,
      COMP_LOOP_COMP_LOOP_and_584_itm, COMP_LOOP_COMP_LOOP_and_836_itm, COMP_LOOP_COMP_LOOP_and_107_itm,
      COMP_LOOP_COMP_LOOP_and_120_itm, COMP_LOOP_COMP_LOOP_and_1592_itm, COMP_LOOP_COMP_LOOP_and_1844_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1286_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_18_itm, COMP_LOOP_COMP_LOOP_and_333_itm,
      COMP_LOOP_COMP_LOOP_and_585_itm, COMP_LOOP_COMP_LOOP_and_837_itm, COMP_LOOP_COMP_LOOP_and_1089_itm,
      COMP_LOOP_COMP_LOOP_and_1341_itm, COMP_LOOP_COMP_LOOP_and_1593_itm, COMP_LOOP_COMP_LOOP_and_1845_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1287_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_272_itm, COMP_LOOP_COMP_LOOP_and_334_itm,
      COMP_LOOP_COMP_LOOP_and_586_itm, COMP_LOOP_COMP_LOOP_and_838_itm, COMP_LOOP_COMP_LOOP_and_108_itm,
      COMP_LOOP_COMP_LOOP_and_121_itm, COMP_LOOP_COMP_LOOP_and_1594_itm, COMP_LOOP_COMP_LOOP_and_1846_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1288_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_20_itm, COMP_LOOP_COMP_LOOP_and_335_itm,
      COMP_LOOP_COMP_LOOP_and_587_itm, COMP_LOOP_COMP_LOOP_and_839_itm, COMP_LOOP_COMP_LOOP_and_1091_itm,
      COMP_LOOP_COMP_LOOP_and_1343_itm, COMP_LOOP_COMP_LOOP_and_1595_itm, COMP_LOOP_COMP_LOOP_and_1847_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1289_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_21_itm, COMP_LOOP_COMP_LOOP_and_336_itm,
      COMP_LOOP_COMP_LOOP_and_588_itm, COMP_LOOP_COMP_LOOP_and_840_itm, COMP_LOOP_COMP_LOOP_and_1092_itm,
      COMP_LOOP_COMP_LOOP_and_1344_itm, COMP_LOOP_COMP_LOOP_and_1596_itm, COMP_LOOP_COMP_LOOP_and_1848_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1290_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_22_itm, COMP_LOOP_COMP_LOOP_and_337_itm,
      COMP_LOOP_COMP_LOOP_and_589_itm, COMP_LOOP_COMP_LOOP_and_841_itm, COMP_LOOP_COMP_LOOP_and_1093_itm,
      COMP_LOOP_COMP_LOOP_and_1345_itm, COMP_LOOP_COMP_LOOP_and_1597_itm, COMP_LOOP_COMP_LOOP_and_1849_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1291_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_23_itm, COMP_LOOP_COMP_LOOP_and_338_itm,
      COMP_LOOP_COMP_LOOP_and_590_itm, COMP_LOOP_COMP_LOOP_and_842_itm, COMP_LOOP_COMP_LOOP_and_109_itm,
      COMP_LOOP_COMP_LOOP_and_1346_itm, COMP_LOOP_COMP_LOOP_and_1598_itm, COMP_LOOP_COMP_LOOP_and_1850_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1292_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_24_itm, COMP_LOOP_COMP_LOOP_and_339_itm,
      COMP_LOOP_COMP_LOOP_and_591_itm, COMP_LOOP_COMP_LOOP_and_843_itm, COMP_LOOP_COMP_LOOP_and_1095_itm,
      COMP_LOOP_COMP_LOOP_and_1347_itm, COMP_LOOP_COMP_LOOP_and_1599_itm, COMP_LOOP_COMP_LOOP_and_1851_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1293_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_25_itm, COMP_LOOP_COMP_LOOP_and_340_itm,
      COMP_LOOP_COMP_LOOP_and_592_itm, COMP_LOOP_COMP_LOOP_and_844_itm, COMP_LOOP_COMP_LOOP_and_1096_itm,
      COMP_LOOP_COMP_LOOP_and_1348_itm, COMP_LOOP_COMP_LOOP_and_1600_itm, COMP_LOOP_COMP_LOOP_and_1852_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1294_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_26_itm, COMP_LOOP_COMP_LOOP_and_341_itm,
      COMP_LOOP_COMP_LOOP_and_593_itm, COMP_LOOP_COMP_LOOP_and_845_itm, COMP_LOOP_COMP_LOOP_and_1097_itm,
      COMP_LOOP_COMP_LOOP_and_1349_itm, COMP_LOOP_COMP_LOOP_and_1601_itm, COMP_LOOP_COMP_LOOP_and_1853_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1295_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_27_itm, COMP_LOOP_COMP_LOOP_and_342_itm,
      COMP_LOOP_COMP_LOOP_and_594_itm, COMP_LOOP_COMP_LOOP_and_846_itm, COMP_LOOP_COMP_LOOP_and_1098_itm,
      COMP_LOOP_COMP_LOOP_and_1350_itm, COMP_LOOP_COMP_LOOP_and_1602_itm, COMP_LOOP_COMP_LOOP_and_1854_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1296_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_28_itm, COMP_LOOP_COMP_LOOP_and_343_itm,
      COMP_LOOP_COMP_LOOP_and_595_itm, COMP_LOOP_COMP_LOOP_and_847_itm, COMP_LOOP_COMP_LOOP_and_1099_itm,
      COMP_LOOP_COMP_LOOP_and_1351_itm, COMP_LOOP_COMP_LOOP_and_1603_itm, COMP_LOOP_COMP_LOOP_and_1855_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1297_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_29_itm, COMP_LOOP_COMP_LOOP_and_344_itm,
      COMP_LOOP_COMP_LOOP_and_596_itm, COMP_LOOP_COMP_LOOP_and_848_itm, COMP_LOOP_COMP_LOOP_and_1100_itm,
      COMP_LOOP_COMP_LOOP_and_1352_itm, COMP_LOOP_COMP_LOOP_and_1604_itm, COMP_LOOP_COMP_LOOP_and_1856_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1298_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_30_itm, COMP_LOOP_COMP_LOOP_and_345_itm,
      COMP_LOOP_COMP_LOOP_and_597_itm, COMP_LOOP_COMP_LOOP_and_849_itm, COMP_LOOP_COMP_LOOP_and_1101_itm,
      COMP_LOOP_COMP_LOOP_and_1353_itm, COMP_LOOP_COMP_LOOP_and_1605_itm, COMP_LOOP_COMP_LOOP_and_1857_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_COMP_LOOP_and_1925_nl <= (COMP_LOOP_acc_10_cse_10_1_2_sva(5)) AND COMP_LOOP_nor_311_itm;
  COMP_LOOP_COMP_LOOP_and_1926_nl <= (COMP_LOOP_acc_10_cse_10_1_3_sva(5)) AND COMP_LOOP_nor_535_itm;
  COMP_LOOP_COMP_LOOP_and_1927_nl <= (COMP_LOOP_acc_10_cse_10_1_4_sva(5)) AND COMP_LOOP_nor_759_itm;
  COMP_LOOP_COMP_LOOP_and_1928_nl <= (COMP_LOOP_acc_10_cse_10_1_5_sva(5)) AND COMP_LOOP_nor_983_itm;
  COMP_LOOP_COMP_LOOP_and_1929_nl <= (COMP_LOOP_acc_10_cse_10_1_6_sva(5)) AND COMP_LOOP_nor_1207_itm;
  COMP_LOOP_COMP_LOOP_and_1930_nl <= (COMP_LOOP_acc_10_cse_10_1_7_sva(5)) AND COMP_LOOP_nor_1431_itm;
  COMP_LOOP_COMP_LOOP_and_1931_nl <= (COMP_LOOP_acc_10_cse_10_1_sva(5)) AND COMP_LOOP_nor_1655_itm;
  COMP_LOOP_mux1h_1299_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_284_itm, COMP_LOOP_COMP_LOOP_and_1925_nl,
      COMP_LOOP_COMP_LOOP_and_1926_nl, COMP_LOOP_COMP_LOOP_and_1927_nl, COMP_LOOP_COMP_LOOP_and_1928_nl,
      COMP_LOOP_COMP_LOOP_and_1929_nl, COMP_LOOP_COMP_LOOP_and_1930_nl, COMP_LOOP_COMP_LOOP_and_1931_nl,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1300_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_285_itm, COMP_LOOP_COMP_LOOP_and_347_itm,
      COMP_LOOP_COMP_LOOP_and_599_itm, COMP_LOOP_COMP_LOOP_and_74_itm, COMP_LOOP_COMP_LOOP_and_110_itm,
      COMP_LOOP_COMP_LOOP_and_122_itm, COMP_LOOP_COMP_LOOP_and_1607_itm, COMP_LOOP_COMP_LOOP_and_1859_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1301_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_286_itm, COMP_LOOP_COMP_LOOP_and_101_itm,
      COMP_LOOP_COMP_LOOP_and_600_itm, COMP_LOOP_COMP_LOOP_and_852_itm, COMP_LOOP_COMP_LOOP_and_1104_itm,
      COMP_LOOP_COMP_LOOP_and_123_itm, COMP_LOOP_COMP_LOOP_and_1608_itm, COMP_LOOP_COMP_LOOP_and_1860_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1302_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_34_itm, COMP_LOOP_COMP_LOOP_and_349_itm,
      COMP_LOOP_COMP_LOOP_and_601_itm, COMP_LOOP_COMP_LOOP_and_853_itm, COMP_LOOP_COMP_LOOP_and_1105_itm,
      COMP_LOOP_COMP_LOOP_and_1357_itm, COMP_LOOP_COMP_LOOP_and_1609_itm, COMP_LOOP_COMP_LOOP_and_1861_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1303_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_288_itm, COMP_LOOP_COMP_LOOP_and_103_itm,
      COMP_LOOP_COMP_LOOP_and_602_itm, COMP_LOOP_COMP_LOOP_and_854_itm, COMP_LOOP_COMP_LOOP_and_1106_itm,
      COMP_LOOP_COMP_LOOP_and_124_itm, COMP_LOOP_COMP_LOOP_and_1610_itm, COMP_LOOP_COMP_LOOP_and_1862_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1304_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_36_itm, COMP_LOOP_COMP_LOOP_and_351_itm,
      COMP_LOOP_COMP_LOOP_and_603_itm, COMP_LOOP_COMP_LOOP_and_855_itm, COMP_LOOP_COMP_LOOP_and_1107_itm,
      COMP_LOOP_COMP_LOOP_and_1359_itm, COMP_LOOP_COMP_LOOP_and_1611_itm, COMP_LOOP_COMP_LOOP_and_1863_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1305_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_37_itm, COMP_LOOP_COMP_LOOP_and_352_itm,
      COMP_LOOP_COMP_LOOP_and_604_itm, COMP_LOOP_COMP_LOOP_and_856_itm, COMP_LOOP_COMP_LOOP_and_1108_itm,
      COMP_LOOP_COMP_LOOP_and_1360_itm, COMP_LOOP_COMP_LOOP_and_1612_itm, COMP_LOOP_COMP_LOOP_and_1864_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1306_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_38_itm, COMP_LOOP_COMP_LOOP_and_353_itm,
      COMP_LOOP_COMP_LOOP_and_605_itm, COMP_LOOP_COMP_LOOP_and_857_itm, COMP_LOOP_COMP_LOOP_and_1109_itm,
      COMP_LOOP_COMP_LOOP_and_1361_itm, COMP_LOOP_COMP_LOOP_and_1613_itm, COMP_LOOP_COMP_LOOP_and_1865_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1307_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_39_itm, COMP_LOOP_COMP_LOOP_and_104_itm,
      COMP_LOOP_COMP_LOOP_and_606_itm, COMP_LOOP_COMP_LOOP_and_75_itm, COMP_LOOP_COMP_LOOP_and_1110_itm,
      COMP_LOOP_COMP_LOOP_and_125_itm, COMP_LOOP_COMP_LOOP_and_1614_itm, COMP_LOOP_COMP_LOOP_and_1866_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1308_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_40_itm, COMP_LOOP_COMP_LOOP_and_355_itm,
      COMP_LOOP_COMP_LOOP_and_607_itm, COMP_LOOP_COMP_LOOP_and_859_itm, COMP_LOOP_COMP_LOOP_and_1111_itm,
      COMP_LOOP_COMP_LOOP_and_1363_itm, COMP_LOOP_COMP_LOOP_and_1615_itm, COMP_LOOP_COMP_LOOP_and_1867_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1309_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_41_itm, COMP_LOOP_COMP_LOOP_and_356_itm,
      COMP_LOOP_COMP_LOOP_and_608_itm, COMP_LOOP_COMP_LOOP_and_860_itm, COMP_LOOP_COMP_LOOP_and_1112_itm,
      COMP_LOOP_COMP_LOOP_and_1364_itm, COMP_LOOP_COMP_LOOP_and_1616_itm, COMP_LOOP_COMP_LOOP_and_1868_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1310_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_42_itm, COMP_LOOP_COMP_LOOP_and_357_itm,
      COMP_LOOP_COMP_LOOP_and_609_itm, COMP_LOOP_COMP_LOOP_and_861_itm, COMP_LOOP_COMP_LOOP_and_1113_itm,
      COMP_LOOP_COMP_LOOP_and_1365_itm, COMP_LOOP_COMP_LOOP_and_1617_itm, COMP_LOOP_COMP_LOOP_and_1869_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1311_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_43_itm, COMP_LOOP_COMP_LOOP_and_358_itm,
      COMP_LOOP_COMP_LOOP_and_610_itm, COMP_LOOP_COMP_LOOP_and_862_itm, COMP_LOOP_COMP_LOOP_and_1114_itm,
      COMP_LOOP_COMP_LOOP_and_1366_itm, COMP_LOOP_COMP_LOOP_and_1618_itm, COMP_LOOP_COMP_LOOP_and_1870_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1312_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_44_itm, COMP_LOOP_COMP_LOOP_and_359_itm,
      COMP_LOOP_COMP_LOOP_and_611_itm, COMP_LOOP_COMP_LOOP_and_863_itm, COMP_LOOP_COMP_LOOP_and_1115_itm,
      COMP_LOOP_COMP_LOOP_and_1367_itm, COMP_LOOP_COMP_LOOP_and_1619_itm, COMP_LOOP_COMP_LOOP_and_1871_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1313_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_45_itm, COMP_LOOP_COMP_LOOP_and_360_itm,
      COMP_LOOP_COMP_LOOP_and_612_itm, COMP_LOOP_COMP_LOOP_and_864_itm, COMP_LOOP_COMP_LOOP_and_1116_itm,
      COMP_LOOP_COMP_LOOP_and_1368_itm, COMP_LOOP_COMP_LOOP_and_1620_itm, COMP_LOOP_COMP_LOOP_and_1872_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1314_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_46_itm, COMP_LOOP_COMP_LOOP_and_361_itm,
      COMP_LOOP_COMP_LOOP_and_613_itm, COMP_LOOP_COMP_LOOP_and_865_itm, COMP_LOOP_COMP_LOOP_and_1117_itm,
      COMP_LOOP_COMP_LOOP_and_1369_itm, COMP_LOOP_COMP_LOOP_and_1621_itm, COMP_LOOP_COMP_LOOP_and_1873_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1315_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_47_itm, COMP_LOOP_COMP_LOOP_and_105_itm,
      COMP_LOOP_COMP_LOOP_and_614_itm, COMP_LOOP_COMP_LOOP_and_866_itm, COMP_LOOP_COMP_LOOP_and_1118_itm,
      COMP_LOOP_COMP_LOOP_and_1370_itm, COMP_LOOP_COMP_LOOP_and_1622_itm, COMP_LOOP_COMP_LOOP_and_1874_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1316_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_48_itm, COMP_LOOP_COMP_LOOP_and_363_itm,
      COMP_LOOP_COMP_LOOP_and_615_itm, COMP_LOOP_COMP_LOOP_and_867_itm, COMP_LOOP_COMP_LOOP_and_1119_itm,
      COMP_LOOP_COMP_LOOP_and_1371_itm, COMP_LOOP_COMP_LOOP_and_1623_itm, COMP_LOOP_COMP_LOOP_and_1875_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1317_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_49_itm, COMP_LOOP_COMP_LOOP_and_364_itm,
      COMP_LOOP_COMP_LOOP_and_616_itm, COMP_LOOP_COMP_LOOP_and_868_itm, COMP_LOOP_COMP_LOOP_and_1120_itm,
      COMP_LOOP_COMP_LOOP_and_1372_itm, COMP_LOOP_COMP_LOOP_and_1624_itm, COMP_LOOP_COMP_LOOP_and_1876_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1318_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_50_itm, COMP_LOOP_COMP_LOOP_and_365_itm,
      COMP_LOOP_COMP_LOOP_and_617_itm, COMP_LOOP_COMP_LOOP_and_869_itm, COMP_LOOP_COMP_LOOP_and_1121_itm,
      COMP_LOOP_COMP_LOOP_and_1373_itm, COMP_LOOP_COMP_LOOP_and_1625_itm, COMP_LOOP_COMP_LOOP_and_1877_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1319_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_51_itm, COMP_LOOP_COMP_LOOP_and_366_itm,
      COMP_LOOP_COMP_LOOP_and_618_itm, COMP_LOOP_COMP_LOOP_and_870_itm, COMP_LOOP_COMP_LOOP_and_1122_itm,
      COMP_LOOP_COMP_LOOP_and_1374_itm, COMP_LOOP_COMP_LOOP_and_1626_itm, COMP_LOOP_COMP_LOOP_and_1878_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1320_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_52_itm, COMP_LOOP_COMP_LOOP_and_367_itm,
      COMP_LOOP_COMP_LOOP_and_619_itm, COMP_LOOP_COMP_LOOP_and_871_itm, COMP_LOOP_COMP_LOOP_and_1123_itm,
      COMP_LOOP_COMP_LOOP_and_1375_itm, COMP_LOOP_COMP_LOOP_and_1627_itm, COMP_LOOP_COMP_LOOP_and_1879_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1321_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_53_itm, COMP_LOOP_COMP_LOOP_and_368_itm,
      COMP_LOOP_COMP_LOOP_and_620_itm, COMP_LOOP_COMP_LOOP_and_872_itm, COMP_LOOP_COMP_LOOP_and_1124_itm,
      COMP_LOOP_COMP_LOOP_and_1376_itm, COMP_LOOP_COMP_LOOP_and_1628_itm, COMP_LOOP_COMP_LOOP_and_1880_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1322_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_54_itm, COMP_LOOP_COMP_LOOP_and_369_itm,
      COMP_LOOP_COMP_LOOP_and_621_itm, COMP_LOOP_COMP_LOOP_and_873_itm, COMP_LOOP_COMP_LOOP_and_1125_itm,
      COMP_LOOP_COMP_LOOP_and_1377_itm, COMP_LOOP_COMP_LOOP_and_1629_itm, COMP_LOOP_COMP_LOOP_and_1881_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1323_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_55_itm, COMP_LOOP_COMP_LOOP_and_370_itm,
      COMP_LOOP_COMP_LOOP_and_622_itm, COMP_LOOP_COMP_LOOP_and_874_itm, COMP_LOOP_COMP_LOOP_and_1126_itm,
      COMP_LOOP_COMP_LOOP_and_1378_itm, COMP_LOOP_COMP_LOOP_and_1630_itm, COMP_LOOP_COMP_LOOP_and_1882_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1324_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_56_itm, COMP_LOOP_COMP_LOOP_and_371_itm,
      COMP_LOOP_COMP_LOOP_and_623_itm, COMP_LOOP_COMP_LOOP_and_875_itm, COMP_LOOP_COMP_LOOP_and_1127_itm,
      COMP_LOOP_COMP_LOOP_and_1379_itm, COMP_LOOP_COMP_LOOP_and_1631_itm, COMP_LOOP_COMP_LOOP_and_1883_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1325_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_57_itm, COMP_LOOP_COMP_LOOP_and_372_itm,
      COMP_LOOP_COMP_LOOP_and_624_itm, COMP_LOOP_COMP_LOOP_and_876_itm, COMP_LOOP_COMP_LOOP_and_1128_itm,
      COMP_LOOP_COMP_LOOP_and_1380_itm, COMP_LOOP_COMP_LOOP_and_1632_itm, COMP_LOOP_COMP_LOOP_and_1884_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1326_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_58_itm, COMP_LOOP_COMP_LOOP_and_373_itm,
      COMP_LOOP_COMP_LOOP_and_625_itm, COMP_LOOP_COMP_LOOP_and_877_itm, COMP_LOOP_COMP_LOOP_and_1129_itm,
      COMP_LOOP_COMP_LOOP_and_1381_itm, COMP_LOOP_COMP_LOOP_and_1633_itm, COMP_LOOP_COMP_LOOP_and_1885_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1327_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_59_itm, COMP_LOOP_COMP_LOOP_and_374_itm,
      COMP_LOOP_COMP_LOOP_and_626_itm, COMP_LOOP_COMP_LOOP_and_878_itm, COMP_LOOP_COMP_LOOP_and_1130_itm,
      COMP_LOOP_COMP_LOOP_and_1382_itm, COMP_LOOP_COMP_LOOP_and_1634_itm, COMP_LOOP_COMP_LOOP_and_1886_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1328_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_60_itm, COMP_LOOP_COMP_LOOP_and_375_itm,
      COMP_LOOP_COMP_LOOP_and_627_itm, COMP_LOOP_COMP_LOOP_and_879_itm, COMP_LOOP_COMP_LOOP_and_1131_itm,
      COMP_LOOP_COMP_LOOP_and_1383_itm, COMP_LOOP_COMP_LOOP_and_1635_itm, COMP_LOOP_COMP_LOOP_and_1887_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1329_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_61_itm, COMP_LOOP_COMP_LOOP_and_376_itm,
      COMP_LOOP_COMP_LOOP_and_628_itm, COMP_LOOP_COMP_LOOP_and_880_itm, COMP_LOOP_COMP_LOOP_and_1132_itm,
      COMP_LOOP_COMP_LOOP_and_1384_itm, COMP_LOOP_COMP_LOOP_and_1636_itm, COMP_LOOP_COMP_LOOP_and_1888_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  COMP_LOOP_mux1h_1330_nl <= MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_62_itm, COMP_LOOP_COMP_LOOP_and_377_itm,
      COMP_LOOP_COMP_LOOP_and_629_itm, COMP_LOOP_COMP_LOOP_and_881_itm, COMP_LOOP_COMP_LOOP_and_1133_itm,
      COMP_LOOP_COMP_LOOP_and_1385_itm, COMP_LOOP_COMP_LOOP_and_1637_itm, COMP_LOOP_COMP_LOOP_and_1889_itm,
      STD_LOGIC_VECTOR'( and_dcpl_632 & and_dcpl_636 & and_903_cse & and_907_cse
      & and_910_cse & and_914_cse & and_918_cse & and_920_cse));
  z_out_9 <= MUX1HOT_v_64_64_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d, vec_rsc_0_2_i_q_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d, vec_rsc_0_6_i_q_d,
      vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d, vec_rsc_0_14_i_q_d,
      vec_rsc_0_15_i_q_d, vec_rsc_0_16_i_q_d, vec_rsc_0_17_i_q_d, vec_rsc_0_18_i_q_d,
      vec_rsc_0_19_i_q_d, vec_rsc_0_20_i_q_d, vec_rsc_0_21_i_q_d, vec_rsc_0_22_i_q_d,
      vec_rsc_0_23_i_q_d, vec_rsc_0_24_i_q_d, vec_rsc_0_25_i_q_d, vec_rsc_0_26_i_q_d,
      vec_rsc_0_27_i_q_d, vec_rsc_0_28_i_q_d, vec_rsc_0_29_i_q_d, vec_rsc_0_30_i_q_d,
      vec_rsc_0_31_i_q_d, vec_rsc_0_32_i_q_d, vec_rsc_0_33_i_q_d, vec_rsc_0_34_i_q_d,
      vec_rsc_0_35_i_q_d, vec_rsc_0_36_i_q_d, vec_rsc_0_37_i_q_d, vec_rsc_0_38_i_q_d,
      vec_rsc_0_39_i_q_d, vec_rsc_0_40_i_q_d, vec_rsc_0_41_i_q_d, vec_rsc_0_42_i_q_d,
      vec_rsc_0_43_i_q_d, vec_rsc_0_44_i_q_d, vec_rsc_0_45_i_q_d, vec_rsc_0_46_i_q_d,
      vec_rsc_0_47_i_q_d, vec_rsc_0_48_i_q_d, vec_rsc_0_49_i_q_d, vec_rsc_0_50_i_q_d,
      vec_rsc_0_51_i_q_d, vec_rsc_0_52_i_q_d, vec_rsc_0_53_i_q_d, vec_rsc_0_54_i_q_d,
      vec_rsc_0_55_i_q_d, vec_rsc_0_56_i_q_d, vec_rsc_0_57_i_q_d, vec_rsc_0_58_i_q_d,
      vec_rsc_0_59_i_q_d, vec_rsc_0_60_i_q_d, vec_rsc_0_61_i_q_d, vec_rsc_0_62_i_q_d,
      vec_rsc_0_63_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_mux1h_1267_nl & COMP_LOOP_mux1h_1268_nl
      & COMP_LOOP_mux1h_1269_nl & COMP_LOOP_mux1h_1270_nl & COMP_LOOP_mux1h_1271_nl
      & COMP_LOOP_mux1h_1272_nl & COMP_LOOP_mux1h_1273_nl & COMP_LOOP_mux1h_1274_nl
      & COMP_LOOP_mux1h_1275_nl & COMP_LOOP_mux1h_1276_nl & COMP_LOOP_mux1h_1277_nl
      & COMP_LOOP_mux1h_1278_nl & COMP_LOOP_mux1h_1279_nl & COMP_LOOP_mux1h_1280_nl
      & COMP_LOOP_mux1h_1281_nl & COMP_LOOP_mux1h_1282_nl & COMP_LOOP_mux1h_1283_nl
      & COMP_LOOP_mux1h_1284_nl & COMP_LOOP_mux1h_1285_nl & COMP_LOOP_mux1h_1286_nl
      & COMP_LOOP_mux1h_1287_nl & COMP_LOOP_mux1h_1288_nl & COMP_LOOP_mux1h_1289_nl
      & COMP_LOOP_mux1h_1290_nl & COMP_LOOP_mux1h_1291_nl & COMP_LOOP_mux1h_1292_nl
      & COMP_LOOP_mux1h_1293_nl & COMP_LOOP_mux1h_1294_nl & COMP_LOOP_mux1h_1295_nl
      & COMP_LOOP_mux1h_1296_nl & COMP_LOOP_mux1h_1297_nl & COMP_LOOP_mux1h_1298_nl
      & COMP_LOOP_mux1h_1299_nl & COMP_LOOP_mux1h_1300_nl & COMP_LOOP_mux1h_1301_nl
      & COMP_LOOP_mux1h_1302_nl & COMP_LOOP_mux1h_1303_nl & COMP_LOOP_mux1h_1304_nl
      & COMP_LOOP_mux1h_1305_nl & COMP_LOOP_mux1h_1306_nl & COMP_LOOP_mux1h_1307_nl
      & COMP_LOOP_mux1h_1308_nl & COMP_LOOP_mux1h_1309_nl & COMP_LOOP_mux1h_1310_nl
      & COMP_LOOP_mux1h_1311_nl & COMP_LOOP_mux1h_1312_nl & COMP_LOOP_mux1h_1313_nl
      & COMP_LOOP_mux1h_1314_nl & COMP_LOOP_mux1h_1315_nl & COMP_LOOP_mux1h_1316_nl
      & COMP_LOOP_mux1h_1317_nl & COMP_LOOP_mux1h_1318_nl & COMP_LOOP_mux1h_1319_nl
      & COMP_LOOP_mux1h_1320_nl & COMP_LOOP_mux1h_1321_nl & COMP_LOOP_mux1h_1322_nl
      & COMP_LOOP_mux1h_1323_nl & COMP_LOOP_mux1h_1324_nl & COMP_LOOP_mux1h_1325_nl
      & COMP_LOOP_mux1h_1326_nl & COMP_LOOP_mux1h_1327_nl & COMP_LOOP_mux1h_1328_nl
      & COMP_LOOP_mux1h_1329_nl & COMP_LOOP_mux1h_1330_nl));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIF
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIF IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_0_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_we : OUT STD_LOGIC;
    vec_rsc_0_0_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_0_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_1_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_we : OUT STD_LOGIC;
    vec_rsc_0_1_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_1_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_2_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_we : OUT STD_LOGIC;
    vec_rsc_0_2_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_2_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_3_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_we : OUT STD_LOGIC;
    vec_rsc_0_3_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_3_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_4_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_we : OUT STD_LOGIC;
    vec_rsc_0_4_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_4_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_5_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_we : OUT STD_LOGIC;
    vec_rsc_0_5_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_5_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_6_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_we : OUT STD_LOGIC;
    vec_rsc_0_6_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_6_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_7_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_we : OUT STD_LOGIC;
    vec_rsc_0_7_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_7_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_0_8_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_8_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_we : OUT STD_LOGIC;
    vec_rsc_0_8_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_8_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_0_9_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_9_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_we : OUT STD_LOGIC;
    vec_rsc_0_9_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_9_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_0_10_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_10_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_we : OUT STD_LOGIC;
    vec_rsc_0_10_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_10_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_0_11_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_11_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_we : OUT STD_LOGIC;
    vec_rsc_0_11_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_11_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_0_12_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_12_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_we : OUT STD_LOGIC;
    vec_rsc_0_12_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_12_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_0_13_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_13_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_we : OUT STD_LOGIC;
    vec_rsc_0_13_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_13_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_0_14_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_14_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_we : OUT STD_LOGIC;
    vec_rsc_0_14_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_14_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_0_15_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_15_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_we : OUT STD_LOGIC;
    vec_rsc_0_15_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_15_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    vec_rsc_0_16_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_16_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_16_we : OUT STD_LOGIC;
    vec_rsc_0_16_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_16_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    vec_rsc_0_17_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_17_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_17_we : OUT STD_LOGIC;
    vec_rsc_0_17_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_17_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    vec_rsc_0_18_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_18_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_18_we : OUT STD_LOGIC;
    vec_rsc_0_18_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_18_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    vec_rsc_0_19_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_19_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_19_we : OUT STD_LOGIC;
    vec_rsc_0_19_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_19_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    vec_rsc_0_20_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_20_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_20_we : OUT STD_LOGIC;
    vec_rsc_0_20_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_20_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    vec_rsc_0_21_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_21_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_21_we : OUT STD_LOGIC;
    vec_rsc_0_21_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_21_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    vec_rsc_0_22_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_22_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_22_we : OUT STD_LOGIC;
    vec_rsc_0_22_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_22_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    vec_rsc_0_23_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_23_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_23_we : OUT STD_LOGIC;
    vec_rsc_0_23_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_23_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    vec_rsc_0_24_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_24_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_24_we : OUT STD_LOGIC;
    vec_rsc_0_24_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_24_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    vec_rsc_0_25_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_25_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_25_we : OUT STD_LOGIC;
    vec_rsc_0_25_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_25_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    vec_rsc_0_26_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_26_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_26_we : OUT STD_LOGIC;
    vec_rsc_0_26_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_26_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    vec_rsc_0_27_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_27_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_27_we : OUT STD_LOGIC;
    vec_rsc_0_27_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_27_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    vec_rsc_0_28_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_28_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_28_we : OUT STD_LOGIC;
    vec_rsc_0_28_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_28_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    vec_rsc_0_29_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_29_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_29_we : OUT STD_LOGIC;
    vec_rsc_0_29_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_29_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    vec_rsc_0_30_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_30_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_30_we : OUT STD_LOGIC;
    vec_rsc_0_30_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_30_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    vec_rsc_0_31_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_31_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_31_we : OUT STD_LOGIC;
    vec_rsc_0_31_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_31_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    vec_rsc_0_32_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_32_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_32_we : OUT STD_LOGIC;
    vec_rsc_0_32_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_32_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_32_lz : OUT STD_LOGIC;
    vec_rsc_0_33_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_33_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_33_we : OUT STD_LOGIC;
    vec_rsc_0_33_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_33_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_33_lz : OUT STD_LOGIC;
    vec_rsc_0_34_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_34_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_34_we : OUT STD_LOGIC;
    vec_rsc_0_34_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_34_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_34_lz : OUT STD_LOGIC;
    vec_rsc_0_35_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_35_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_35_we : OUT STD_LOGIC;
    vec_rsc_0_35_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_35_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_35_lz : OUT STD_LOGIC;
    vec_rsc_0_36_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_36_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_36_we : OUT STD_LOGIC;
    vec_rsc_0_36_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_36_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_36_lz : OUT STD_LOGIC;
    vec_rsc_0_37_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_37_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_37_we : OUT STD_LOGIC;
    vec_rsc_0_37_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_37_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_37_lz : OUT STD_LOGIC;
    vec_rsc_0_38_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_38_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_38_we : OUT STD_LOGIC;
    vec_rsc_0_38_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_38_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_38_lz : OUT STD_LOGIC;
    vec_rsc_0_39_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_39_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_39_we : OUT STD_LOGIC;
    vec_rsc_0_39_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_39_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_39_lz : OUT STD_LOGIC;
    vec_rsc_0_40_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_40_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_40_we : OUT STD_LOGIC;
    vec_rsc_0_40_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_40_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_40_lz : OUT STD_LOGIC;
    vec_rsc_0_41_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_41_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_41_we : OUT STD_LOGIC;
    vec_rsc_0_41_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_41_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_41_lz : OUT STD_LOGIC;
    vec_rsc_0_42_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_42_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_42_we : OUT STD_LOGIC;
    vec_rsc_0_42_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_42_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_42_lz : OUT STD_LOGIC;
    vec_rsc_0_43_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_43_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_43_we : OUT STD_LOGIC;
    vec_rsc_0_43_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_43_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_43_lz : OUT STD_LOGIC;
    vec_rsc_0_44_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_44_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_44_we : OUT STD_LOGIC;
    vec_rsc_0_44_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_44_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_44_lz : OUT STD_LOGIC;
    vec_rsc_0_45_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_45_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_45_we : OUT STD_LOGIC;
    vec_rsc_0_45_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_45_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_45_lz : OUT STD_LOGIC;
    vec_rsc_0_46_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_46_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_46_we : OUT STD_LOGIC;
    vec_rsc_0_46_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_46_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_46_lz : OUT STD_LOGIC;
    vec_rsc_0_47_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_47_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_47_we : OUT STD_LOGIC;
    vec_rsc_0_47_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_47_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_47_lz : OUT STD_LOGIC;
    vec_rsc_0_48_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_48_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_48_we : OUT STD_LOGIC;
    vec_rsc_0_48_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_48_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_48_lz : OUT STD_LOGIC;
    vec_rsc_0_49_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_49_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_49_we : OUT STD_LOGIC;
    vec_rsc_0_49_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_49_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_49_lz : OUT STD_LOGIC;
    vec_rsc_0_50_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_50_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_50_we : OUT STD_LOGIC;
    vec_rsc_0_50_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_50_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_50_lz : OUT STD_LOGIC;
    vec_rsc_0_51_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_51_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_51_we : OUT STD_LOGIC;
    vec_rsc_0_51_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_51_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_51_lz : OUT STD_LOGIC;
    vec_rsc_0_52_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_52_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_52_we : OUT STD_LOGIC;
    vec_rsc_0_52_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_52_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_52_lz : OUT STD_LOGIC;
    vec_rsc_0_53_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_53_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_53_we : OUT STD_LOGIC;
    vec_rsc_0_53_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_53_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_53_lz : OUT STD_LOGIC;
    vec_rsc_0_54_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_54_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_54_we : OUT STD_LOGIC;
    vec_rsc_0_54_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_54_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_54_lz : OUT STD_LOGIC;
    vec_rsc_0_55_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_55_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_55_we : OUT STD_LOGIC;
    vec_rsc_0_55_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_55_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_55_lz : OUT STD_LOGIC;
    vec_rsc_0_56_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_56_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_56_we : OUT STD_LOGIC;
    vec_rsc_0_56_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_56_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_56_lz : OUT STD_LOGIC;
    vec_rsc_0_57_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_57_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_57_we : OUT STD_LOGIC;
    vec_rsc_0_57_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_57_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_57_lz : OUT STD_LOGIC;
    vec_rsc_0_58_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_58_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_58_we : OUT STD_LOGIC;
    vec_rsc_0_58_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_58_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_58_lz : OUT STD_LOGIC;
    vec_rsc_0_59_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_59_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_59_we : OUT STD_LOGIC;
    vec_rsc_0_59_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_59_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_59_lz : OUT STD_LOGIC;
    vec_rsc_0_60_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_60_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_60_we : OUT STD_LOGIC;
    vec_rsc_0_60_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_60_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_60_lz : OUT STD_LOGIC;
    vec_rsc_0_61_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_61_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_61_we : OUT STD_LOGIC;
    vec_rsc_0_61_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_61_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_61_lz : OUT STD_LOGIC;
    vec_rsc_0_62_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_62_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_62_we : OUT STD_LOGIC;
    vec_rsc_0_62_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_62_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_62_lz : OUT STD_LOGIC;
    vec_rsc_0_63_wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_63_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_63_we : OUT STD_LOGIC;
    vec_rsc_0_63_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    vec_rsc_0_63_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_63_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_0_0_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_0_1_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_0_2_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_0_3_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_0_4_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_0_5_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_0_6_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_0_7_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_0_8_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_0_9_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_0_10_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_0_11_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_0_12_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_0_13_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_0_14_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_0_15_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_rsc_0_16_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_16_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    twiddle_rsc_0_17_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_17_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    twiddle_rsc_0_18_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_18_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    twiddle_rsc_0_19_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_19_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    twiddle_rsc_0_20_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_20_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    twiddle_rsc_0_21_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_21_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    twiddle_rsc_0_22_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_22_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    twiddle_rsc_0_23_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_23_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    twiddle_rsc_0_24_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_24_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    twiddle_rsc_0_25_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_25_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    twiddle_rsc_0_26_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_26_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    twiddle_rsc_0_27_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_27_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    twiddle_rsc_0_28_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_28_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    twiddle_rsc_0_29_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_29_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    twiddle_rsc_0_30_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_30_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    twiddle_rsc_0_31_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_31_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    twiddle_rsc_0_32_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_32_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_32_lz : OUT STD_LOGIC;
    twiddle_rsc_0_33_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_33_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_33_lz : OUT STD_LOGIC;
    twiddle_rsc_0_34_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_34_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_34_lz : OUT STD_LOGIC;
    twiddle_rsc_0_35_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_35_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_35_lz : OUT STD_LOGIC;
    twiddle_rsc_0_36_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_36_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_36_lz : OUT STD_LOGIC;
    twiddle_rsc_0_37_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_37_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_37_lz : OUT STD_LOGIC;
    twiddle_rsc_0_38_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_38_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_38_lz : OUT STD_LOGIC;
    twiddle_rsc_0_39_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_39_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_39_lz : OUT STD_LOGIC;
    twiddle_rsc_0_40_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_40_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_40_lz : OUT STD_LOGIC;
    twiddle_rsc_0_41_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_41_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_41_lz : OUT STD_LOGIC;
    twiddle_rsc_0_42_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_42_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_42_lz : OUT STD_LOGIC;
    twiddle_rsc_0_43_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_43_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_43_lz : OUT STD_LOGIC;
    twiddle_rsc_0_44_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_44_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_44_lz : OUT STD_LOGIC;
    twiddle_rsc_0_45_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_45_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_45_lz : OUT STD_LOGIC;
    twiddle_rsc_0_46_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_46_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_46_lz : OUT STD_LOGIC;
    twiddle_rsc_0_47_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_47_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_47_lz : OUT STD_LOGIC;
    twiddle_rsc_0_48_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_48_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_48_lz : OUT STD_LOGIC;
    twiddle_rsc_0_49_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_49_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_49_lz : OUT STD_LOGIC;
    twiddle_rsc_0_50_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_50_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_50_lz : OUT STD_LOGIC;
    twiddle_rsc_0_51_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_51_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_51_lz : OUT STD_LOGIC;
    twiddle_rsc_0_52_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_52_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_52_lz : OUT STD_LOGIC;
    twiddle_rsc_0_53_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_53_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_53_lz : OUT STD_LOGIC;
    twiddle_rsc_0_54_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_54_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_54_lz : OUT STD_LOGIC;
    twiddle_rsc_0_55_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_55_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_55_lz : OUT STD_LOGIC;
    twiddle_rsc_0_56_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_56_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_56_lz : OUT STD_LOGIC;
    twiddle_rsc_0_57_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_57_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_57_lz : OUT STD_LOGIC;
    twiddle_rsc_0_58_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_58_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_58_lz : OUT STD_LOGIC;
    twiddle_rsc_0_59_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_59_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_59_lz : OUT STD_LOGIC;
    twiddle_rsc_0_60_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_60_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_60_lz : OUT STD_LOGIC;
    twiddle_rsc_0_61_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_61_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_61_lz : OUT STD_LOGIC;
    twiddle_rsc_0_62_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_62_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_62_lz : OUT STD_LOGIC;
    twiddle_rsc_0_63_radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_63_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    twiddle_rsc_triosy_0_63_lz : OUT STD_LOGIC
  );
END inPlaceNTT_DIF;

ARCHITECTURE v14 OF inPlaceNTT_DIF IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_32_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_33_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_34_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_35_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_36_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_37_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_38_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_39_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_40_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_41_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_42_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_43_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_44_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_45_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_46_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_47_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_48_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_49_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_50_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_51_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_52_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_53_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_54_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_55_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_56_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_57_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_58_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_59_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_60_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_61_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_62_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_63_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_32_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_33_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_34_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_35_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_36_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_37_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_38_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_39_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_40_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_41_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_42_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_43_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_44_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_45_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_46_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_47_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_48_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_49_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_50_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_51_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_52_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_53_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_54_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_55_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_56_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_57_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_58_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_59_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_60_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_61_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_62_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_rsc_0_63_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_d_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_16_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_17_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_18_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_19_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_20_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_21_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_22_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_23_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_24_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_25_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_26_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_27_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_28_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_29_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_30_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_31_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_32_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_33_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_34_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_35_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_36_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_37_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_38_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_39_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_40_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_41_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_42_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_43_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_44_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_45_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_46_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_47_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_48_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_49_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_50_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_51_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_52_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_53_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_54_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_55_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_56_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_57_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_58_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_59_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_60_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_61_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_62_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_63_i_we_d_iff : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_radr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_radr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_8_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_9_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_10_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_11_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_12_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_13_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_14_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_15_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_16_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_16_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_17_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_17_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_18_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_18_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_19_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_19_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_20_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_20_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_21_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_21_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_22_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_22_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_23_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_23_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_24_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_24_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_25_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_25_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_26_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_26_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_27_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_27_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_28_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_28_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_29_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_29_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_30_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_30_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_31_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_31_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_32_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_32_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_32_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_32_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_32_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_32_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_32_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_32_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_33_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_33_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_33_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_33_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_33_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_33_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_33_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_33_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_34_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_34_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_34_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_34_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_34_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_34_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_34_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_34_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_35_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_35_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_35_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_35_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_35_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_35_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_35_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_35_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_36_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_36_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_36_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_36_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_36_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_36_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_36_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_36_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_37_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_37_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_37_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_37_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_37_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_37_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_37_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_37_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_38_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_38_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_38_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_38_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_38_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_38_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_38_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_38_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_39_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_39_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_39_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_39_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_39_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_39_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_39_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_39_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_40_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_40_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_40_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_40_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_40_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_40_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_40_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_40_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_41_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_41_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_41_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_41_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_41_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_41_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_41_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_41_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_42_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_42_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_42_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_42_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_42_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_42_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_42_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_42_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_43_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_43_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_43_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_43_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_43_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_43_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_43_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_43_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_44_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_44_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_44_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_44_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_44_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_44_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_44_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_44_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_45_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_45_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_45_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_45_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_45_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_45_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_45_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_45_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_46_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_46_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_46_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_46_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_46_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_46_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_46_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_46_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_47_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_47_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_47_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_47_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_47_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_47_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_47_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_47_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_48_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_48_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_48_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_48_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_48_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_48_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_48_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_48_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_49_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_49_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_49_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_49_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_49_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_49_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_49_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_49_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_50_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_50_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_50_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_50_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_50_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_50_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_50_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_50_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_51_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_51_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_51_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_51_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_51_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_51_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_51_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_51_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_52_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_52_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_52_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_52_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_52_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_52_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_52_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_52_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_53_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_53_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_53_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_53_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_53_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_53_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_53_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_53_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_54_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_54_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_54_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_54_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_54_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_54_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_54_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_54_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_55_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_55_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_55_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_55_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_55_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_55_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_55_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_55_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_56_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_56_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_56_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_56_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_56_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_56_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_56_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_56_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_57_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_57_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_57_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_57_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_57_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_57_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_57_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_57_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_58_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_58_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_58_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_58_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_58_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_58_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_58_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_58_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_59_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_59_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_59_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_59_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_59_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_59_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_59_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_59_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_60_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_60_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_60_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_60_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_60_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_60_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_60_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_60_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_61_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_61_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_61_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_61_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_61_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_61_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_61_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_61_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_62_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_62_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_62_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_62_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_62_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_62_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_62_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_62_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_63_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_63_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_63_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_63_i_wadr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_63_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_63_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_63_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL vec_rsc_0_63_i_wadr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_0_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_1_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_2_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_3_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_4_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_5_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_6_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_7_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_8_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_9_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_10_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_11_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_12_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_13_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_14_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_15_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_16_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_16_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_16_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_16_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_17_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_17_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_17_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_17_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_18_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_18_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_18_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_18_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_19_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_19_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_19_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_19_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_20_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_20_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_20_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_20_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_21_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_21_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_21_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_21_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_22_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_22_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_22_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_22_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_23_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_23_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_23_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_23_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_24_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_24_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_24_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_24_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_25_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_25_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_25_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_25_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_26_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_26_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_26_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_26_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_27_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_27_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_27_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_27_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_28_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_28_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_28_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_28_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_29_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_29_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_29_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_29_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_30_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_30_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_30_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_30_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_31_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_31_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_31_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_31_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_32_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_32_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_32_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_32_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_33_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_33_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_33_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_33_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_34_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_34_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_34_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_34_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_35_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_35_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_35_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_35_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_36_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_36_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_36_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_36_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_37_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_37_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_37_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_37_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_38_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_38_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_38_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_38_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_39_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_39_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_39_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_39_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_40_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_40_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_40_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_40_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_41_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_41_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_41_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_41_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_42_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_42_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_42_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_42_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_43_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_43_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_43_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_43_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_44_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_44_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_44_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_44_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_45_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_45_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_45_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_45_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_46_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_46_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_46_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_46_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_47_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_47_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_47_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_47_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_48_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_48_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_48_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_48_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_49_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_49_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_49_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_49_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_50_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_50_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_50_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_50_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_51_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_51_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_51_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_51_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_52_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_52_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_52_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_52_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_53_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_53_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_53_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_53_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_54_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_54_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_54_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_54_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_55_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_55_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_55_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_55_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_56_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_56_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_56_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_56_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_57_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_57_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_57_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_57_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_58_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_58_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_58_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_58_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_59_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_59_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_59_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_59_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_60_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_60_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_60_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_60_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_61_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_61_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_61_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_61_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_62_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_62_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_62_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_62_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsc_0_63_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_63_i_radr : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_63_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL twiddle_rsc_0_63_i_radr_d : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT inPlaceNTT_DIF_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_16_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_17_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_18_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_19_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_20_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_21_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_22_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_23_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_24_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_25_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_26_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_27_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_28_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_29_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_30_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_31_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_32_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_33_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_34_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_35_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_36_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_37_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_38_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_39_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_40_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_41_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_42_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_43_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_44_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_45_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_46_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_47_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_48_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_49_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_50_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_51_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_52_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_53_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_54_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_55_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_56_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_57_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_58_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_59_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_60_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_61_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_62_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_63_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_16_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_17_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_18_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_19_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_20_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_21_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_22_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_23_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_24_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_25_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_26_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_27_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_28_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_29_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_30_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_31_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_32_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_33_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_34_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_35_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_36_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_37_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_38_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_39_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_40_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_41_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_42_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_43_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_44_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_45_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_46_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_47_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_48_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_49_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_50_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_51_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_52_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_53_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_54_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_55_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_56_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_57_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_58_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_59_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_60_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_61_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_62_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_0_63_lz : OUT STD_LOGIC;
      vec_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_32_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_33_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_34_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_35_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_36_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_37_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_38_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_39_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_40_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_41_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_42_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_43_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_44_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_45_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_46_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_47_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_48_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_49_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_50_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_51_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_52_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_53_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_54_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_55_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_56_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_57_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_58_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_59_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_60_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_61_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_62_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_63_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_16_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_17_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_18_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_19_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_20_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_21_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_22_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_23_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_24_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_25_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_26_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_27_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_28_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_29_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_30_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_31_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_32_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_33_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_34_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_35_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_36_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_37_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_38_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_39_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_40_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_41_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_42_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_43_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_44_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_45_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_46_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_47_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_48_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_49_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_50_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_51_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_52_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_53_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_54_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_55_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_56_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_57_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_58_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_59_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_60_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_61_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_62_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_rsc_0_63_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      vec_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      vec_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_1_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_2_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_3_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_4_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_5_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_6_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_7_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_8_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_9_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_10_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_11_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_12_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_13_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_14_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_15_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_16_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_17_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_18_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_19_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_20_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_21_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_22_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_23_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_24_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_25_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_26_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_27_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_28_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_29_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_30_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_31_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_32_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_33_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_34_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_35_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_36_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_37_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_38_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_39_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_40_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_41_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_42_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_43_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_44_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_45_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_46_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_47_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_48_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_49_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_50_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_51_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_52_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_53_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_54_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_55_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_56_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_57_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_58_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_59_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_60_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_61_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_62_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_63_i_we_d_pff : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_i_radr_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIF_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_32_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_33_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_34_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_35_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_36_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_37_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_38_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_39_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_40_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_41_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_42_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_43_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_44_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_45_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_46_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_47_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_48_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_49_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_50_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_51_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_52_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_53_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_54_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_55_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_56_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_57_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_58_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_59_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_60_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_61_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_62_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_63_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_16_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_17_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_18_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_19_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_20_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_21_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_22_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_23_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_24_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_25_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_26_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_27_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_28_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_29_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_30_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_31_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_32_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_33_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_34_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_35_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_36_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_37_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_38_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_39_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_40_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_41_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_42_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_43_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_44_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_45_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_46_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_47_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_48_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_49_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_50_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_51_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_52_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_53_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_54_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_55_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_56_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_57_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_58_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_59_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_60_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_61_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_62_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_63_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d_pff : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff : STD_LOGIC_VECTOR
      (3 DOWNTO 0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_0_i_q,
      radr => vec_rsc_0_0_i_radr,
      we => vec_rsc_0_0_we,
      d => vec_rsc_0_0_i_d,
      wadr => vec_rsc_0_0_i_wadr,
      d_d => vec_rsc_0_0_i_d_d,
      q_d => vec_rsc_0_0_i_q_d_1,
      radr_d => vec_rsc_0_0_i_radr_d,
      wadr_d => vec_rsc_0_0_i_wadr_d,
      we_d => vec_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_0_i_q <= vec_rsc_0_0_q;
  vec_rsc_0_0_radr <= vec_rsc_0_0_i_radr;
  vec_rsc_0_0_d <= vec_rsc_0_0_i_d;
  vec_rsc_0_0_wadr <= vec_rsc_0_0_i_wadr;
  vec_rsc_0_0_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_0_i_q_d <= vec_rsc_0_0_i_q_d_1;
  vec_rsc_0_0_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_0_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_1_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_1_i_q,
      radr => vec_rsc_0_1_i_radr,
      we => vec_rsc_0_1_we,
      d => vec_rsc_0_1_i_d,
      wadr => vec_rsc_0_1_i_wadr,
      d_d => vec_rsc_0_1_i_d_d,
      q_d => vec_rsc_0_1_i_q_d_1,
      radr_d => vec_rsc_0_1_i_radr_d,
      wadr_d => vec_rsc_0_1_i_wadr_d,
      we_d => vec_rsc_0_1_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_1_i_q <= vec_rsc_0_1_q;
  vec_rsc_0_1_radr <= vec_rsc_0_1_i_radr;
  vec_rsc_0_1_d <= vec_rsc_0_1_i_d;
  vec_rsc_0_1_wadr <= vec_rsc_0_1_i_wadr;
  vec_rsc_0_1_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_1_i_q_d <= vec_rsc_0_1_i_q_d_1;
  vec_rsc_0_1_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_1_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_2_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_2_i_q,
      radr => vec_rsc_0_2_i_radr,
      we => vec_rsc_0_2_we,
      d => vec_rsc_0_2_i_d,
      wadr => vec_rsc_0_2_i_wadr,
      d_d => vec_rsc_0_2_i_d_d,
      q_d => vec_rsc_0_2_i_q_d_1,
      radr_d => vec_rsc_0_2_i_radr_d,
      wadr_d => vec_rsc_0_2_i_wadr_d,
      we_d => vec_rsc_0_2_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_2_i_q <= vec_rsc_0_2_q;
  vec_rsc_0_2_radr <= vec_rsc_0_2_i_radr;
  vec_rsc_0_2_d <= vec_rsc_0_2_i_d;
  vec_rsc_0_2_wadr <= vec_rsc_0_2_i_wadr;
  vec_rsc_0_2_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_2_i_q_d <= vec_rsc_0_2_i_q_d_1;
  vec_rsc_0_2_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_2_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_3_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_3_i_q,
      radr => vec_rsc_0_3_i_radr,
      we => vec_rsc_0_3_we,
      d => vec_rsc_0_3_i_d,
      wadr => vec_rsc_0_3_i_wadr,
      d_d => vec_rsc_0_3_i_d_d,
      q_d => vec_rsc_0_3_i_q_d_1,
      radr_d => vec_rsc_0_3_i_radr_d,
      wadr_d => vec_rsc_0_3_i_wadr_d,
      we_d => vec_rsc_0_3_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_3_i_q <= vec_rsc_0_3_q;
  vec_rsc_0_3_radr <= vec_rsc_0_3_i_radr;
  vec_rsc_0_3_d <= vec_rsc_0_3_i_d;
  vec_rsc_0_3_wadr <= vec_rsc_0_3_i_wadr;
  vec_rsc_0_3_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_3_i_q_d <= vec_rsc_0_3_i_q_d_1;
  vec_rsc_0_3_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_3_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_4_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_4_i_q,
      radr => vec_rsc_0_4_i_radr,
      we => vec_rsc_0_4_we,
      d => vec_rsc_0_4_i_d,
      wadr => vec_rsc_0_4_i_wadr,
      d_d => vec_rsc_0_4_i_d_d,
      q_d => vec_rsc_0_4_i_q_d_1,
      radr_d => vec_rsc_0_4_i_radr_d,
      wadr_d => vec_rsc_0_4_i_wadr_d,
      we_d => vec_rsc_0_4_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_4_i_q <= vec_rsc_0_4_q;
  vec_rsc_0_4_radr <= vec_rsc_0_4_i_radr;
  vec_rsc_0_4_d <= vec_rsc_0_4_i_d;
  vec_rsc_0_4_wadr <= vec_rsc_0_4_i_wadr;
  vec_rsc_0_4_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_4_i_q_d <= vec_rsc_0_4_i_q_d_1;
  vec_rsc_0_4_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_4_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_5_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_5_i_q,
      radr => vec_rsc_0_5_i_radr,
      we => vec_rsc_0_5_we,
      d => vec_rsc_0_5_i_d,
      wadr => vec_rsc_0_5_i_wadr,
      d_d => vec_rsc_0_5_i_d_d,
      q_d => vec_rsc_0_5_i_q_d_1,
      radr_d => vec_rsc_0_5_i_radr_d,
      wadr_d => vec_rsc_0_5_i_wadr_d,
      we_d => vec_rsc_0_5_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_5_i_q <= vec_rsc_0_5_q;
  vec_rsc_0_5_radr <= vec_rsc_0_5_i_radr;
  vec_rsc_0_5_d <= vec_rsc_0_5_i_d;
  vec_rsc_0_5_wadr <= vec_rsc_0_5_i_wadr;
  vec_rsc_0_5_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_5_i_q_d <= vec_rsc_0_5_i_q_d_1;
  vec_rsc_0_5_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_5_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_6_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_6_i_q,
      radr => vec_rsc_0_6_i_radr,
      we => vec_rsc_0_6_we,
      d => vec_rsc_0_6_i_d,
      wadr => vec_rsc_0_6_i_wadr,
      d_d => vec_rsc_0_6_i_d_d,
      q_d => vec_rsc_0_6_i_q_d_1,
      radr_d => vec_rsc_0_6_i_radr_d,
      wadr_d => vec_rsc_0_6_i_wadr_d,
      we_d => vec_rsc_0_6_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_6_i_q <= vec_rsc_0_6_q;
  vec_rsc_0_6_radr <= vec_rsc_0_6_i_radr;
  vec_rsc_0_6_d <= vec_rsc_0_6_i_d;
  vec_rsc_0_6_wadr <= vec_rsc_0_6_i_wadr;
  vec_rsc_0_6_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_6_i_q_d <= vec_rsc_0_6_i_q_d_1;
  vec_rsc_0_6_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_6_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_7_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_7_i_q,
      radr => vec_rsc_0_7_i_radr,
      we => vec_rsc_0_7_we,
      d => vec_rsc_0_7_i_d,
      wadr => vec_rsc_0_7_i_wadr,
      d_d => vec_rsc_0_7_i_d_d,
      q_d => vec_rsc_0_7_i_q_d_1,
      radr_d => vec_rsc_0_7_i_radr_d,
      wadr_d => vec_rsc_0_7_i_wadr_d,
      we_d => vec_rsc_0_7_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_7_i_q <= vec_rsc_0_7_q;
  vec_rsc_0_7_radr <= vec_rsc_0_7_i_radr;
  vec_rsc_0_7_d <= vec_rsc_0_7_i_d;
  vec_rsc_0_7_wadr <= vec_rsc_0_7_i_wadr;
  vec_rsc_0_7_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_7_i_q_d <= vec_rsc_0_7_i_q_d_1;
  vec_rsc_0_7_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_7_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_8_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_8_i_q,
      radr => vec_rsc_0_8_i_radr,
      we => vec_rsc_0_8_we,
      d => vec_rsc_0_8_i_d,
      wadr => vec_rsc_0_8_i_wadr,
      d_d => vec_rsc_0_8_i_d_d,
      q_d => vec_rsc_0_8_i_q_d_1,
      radr_d => vec_rsc_0_8_i_radr_d,
      wadr_d => vec_rsc_0_8_i_wadr_d,
      we_d => vec_rsc_0_8_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_8_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_8_i_q <= vec_rsc_0_8_q;
  vec_rsc_0_8_radr <= vec_rsc_0_8_i_radr;
  vec_rsc_0_8_d <= vec_rsc_0_8_i_d;
  vec_rsc_0_8_wadr <= vec_rsc_0_8_i_wadr;
  vec_rsc_0_8_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_8_i_q_d <= vec_rsc_0_8_i_q_d_1;
  vec_rsc_0_8_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_8_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_9_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_9_i_q,
      radr => vec_rsc_0_9_i_radr,
      we => vec_rsc_0_9_we,
      d => vec_rsc_0_9_i_d,
      wadr => vec_rsc_0_9_i_wadr,
      d_d => vec_rsc_0_9_i_d_d,
      q_d => vec_rsc_0_9_i_q_d_1,
      radr_d => vec_rsc_0_9_i_radr_d,
      wadr_d => vec_rsc_0_9_i_wadr_d,
      we_d => vec_rsc_0_9_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_9_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_9_i_q <= vec_rsc_0_9_q;
  vec_rsc_0_9_radr <= vec_rsc_0_9_i_radr;
  vec_rsc_0_9_d <= vec_rsc_0_9_i_d;
  vec_rsc_0_9_wadr <= vec_rsc_0_9_i_wadr;
  vec_rsc_0_9_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_9_i_q_d <= vec_rsc_0_9_i_q_d_1;
  vec_rsc_0_9_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_9_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_10_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_10_i_q,
      radr => vec_rsc_0_10_i_radr,
      we => vec_rsc_0_10_we,
      d => vec_rsc_0_10_i_d,
      wadr => vec_rsc_0_10_i_wadr,
      d_d => vec_rsc_0_10_i_d_d,
      q_d => vec_rsc_0_10_i_q_d_1,
      radr_d => vec_rsc_0_10_i_radr_d,
      wadr_d => vec_rsc_0_10_i_wadr_d,
      we_d => vec_rsc_0_10_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_10_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_10_i_q <= vec_rsc_0_10_q;
  vec_rsc_0_10_radr <= vec_rsc_0_10_i_radr;
  vec_rsc_0_10_d <= vec_rsc_0_10_i_d;
  vec_rsc_0_10_wadr <= vec_rsc_0_10_i_wadr;
  vec_rsc_0_10_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_10_i_q_d <= vec_rsc_0_10_i_q_d_1;
  vec_rsc_0_10_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_10_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_11_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_11_i_q,
      radr => vec_rsc_0_11_i_radr,
      we => vec_rsc_0_11_we,
      d => vec_rsc_0_11_i_d,
      wadr => vec_rsc_0_11_i_wadr,
      d_d => vec_rsc_0_11_i_d_d,
      q_d => vec_rsc_0_11_i_q_d_1,
      radr_d => vec_rsc_0_11_i_radr_d,
      wadr_d => vec_rsc_0_11_i_wadr_d,
      we_d => vec_rsc_0_11_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_11_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_11_i_q <= vec_rsc_0_11_q;
  vec_rsc_0_11_radr <= vec_rsc_0_11_i_radr;
  vec_rsc_0_11_d <= vec_rsc_0_11_i_d;
  vec_rsc_0_11_wadr <= vec_rsc_0_11_i_wadr;
  vec_rsc_0_11_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_11_i_q_d <= vec_rsc_0_11_i_q_d_1;
  vec_rsc_0_11_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_11_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_12_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_12_i_q,
      radr => vec_rsc_0_12_i_radr,
      we => vec_rsc_0_12_we,
      d => vec_rsc_0_12_i_d,
      wadr => vec_rsc_0_12_i_wadr,
      d_d => vec_rsc_0_12_i_d_d,
      q_d => vec_rsc_0_12_i_q_d_1,
      radr_d => vec_rsc_0_12_i_radr_d,
      wadr_d => vec_rsc_0_12_i_wadr_d,
      we_d => vec_rsc_0_12_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_12_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_12_i_q <= vec_rsc_0_12_q;
  vec_rsc_0_12_radr <= vec_rsc_0_12_i_radr;
  vec_rsc_0_12_d <= vec_rsc_0_12_i_d;
  vec_rsc_0_12_wadr <= vec_rsc_0_12_i_wadr;
  vec_rsc_0_12_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_12_i_q_d <= vec_rsc_0_12_i_q_d_1;
  vec_rsc_0_12_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_12_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_13_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_13_i_q,
      radr => vec_rsc_0_13_i_radr,
      we => vec_rsc_0_13_we,
      d => vec_rsc_0_13_i_d,
      wadr => vec_rsc_0_13_i_wadr,
      d_d => vec_rsc_0_13_i_d_d,
      q_d => vec_rsc_0_13_i_q_d_1,
      radr_d => vec_rsc_0_13_i_radr_d,
      wadr_d => vec_rsc_0_13_i_wadr_d,
      we_d => vec_rsc_0_13_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_13_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_13_i_q <= vec_rsc_0_13_q;
  vec_rsc_0_13_radr <= vec_rsc_0_13_i_radr;
  vec_rsc_0_13_d <= vec_rsc_0_13_i_d;
  vec_rsc_0_13_wadr <= vec_rsc_0_13_i_wadr;
  vec_rsc_0_13_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_13_i_q_d <= vec_rsc_0_13_i_q_d_1;
  vec_rsc_0_13_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_13_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_14_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_14_i_q,
      radr => vec_rsc_0_14_i_radr,
      we => vec_rsc_0_14_we,
      d => vec_rsc_0_14_i_d,
      wadr => vec_rsc_0_14_i_wadr,
      d_d => vec_rsc_0_14_i_d_d,
      q_d => vec_rsc_0_14_i_q_d_1,
      radr_d => vec_rsc_0_14_i_radr_d,
      wadr_d => vec_rsc_0_14_i_wadr_d,
      we_d => vec_rsc_0_14_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_14_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_14_i_q <= vec_rsc_0_14_q;
  vec_rsc_0_14_radr <= vec_rsc_0_14_i_radr;
  vec_rsc_0_14_d <= vec_rsc_0_14_i_d;
  vec_rsc_0_14_wadr <= vec_rsc_0_14_i_wadr;
  vec_rsc_0_14_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_14_i_q_d <= vec_rsc_0_14_i_q_d_1;
  vec_rsc_0_14_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_14_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_15_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_15_i_q,
      radr => vec_rsc_0_15_i_radr,
      we => vec_rsc_0_15_we,
      d => vec_rsc_0_15_i_d,
      wadr => vec_rsc_0_15_i_wadr,
      d_d => vec_rsc_0_15_i_d_d,
      q_d => vec_rsc_0_15_i_q_d_1,
      radr_d => vec_rsc_0_15_i_radr_d,
      wadr_d => vec_rsc_0_15_i_wadr_d,
      we_d => vec_rsc_0_15_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_15_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_15_i_q <= vec_rsc_0_15_q;
  vec_rsc_0_15_radr <= vec_rsc_0_15_i_radr;
  vec_rsc_0_15_d <= vec_rsc_0_15_i_d;
  vec_rsc_0_15_wadr <= vec_rsc_0_15_i_wadr;
  vec_rsc_0_15_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_15_i_q_d <= vec_rsc_0_15_i_q_d_1;
  vec_rsc_0_15_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_15_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_16_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_16_i_q,
      radr => vec_rsc_0_16_i_radr,
      we => vec_rsc_0_16_we,
      d => vec_rsc_0_16_i_d,
      wadr => vec_rsc_0_16_i_wadr,
      d_d => vec_rsc_0_16_i_d_d,
      q_d => vec_rsc_0_16_i_q_d_1,
      radr_d => vec_rsc_0_16_i_radr_d,
      wadr_d => vec_rsc_0_16_i_wadr_d,
      we_d => vec_rsc_0_16_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_16_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_16_i_q <= vec_rsc_0_16_q;
  vec_rsc_0_16_radr <= vec_rsc_0_16_i_radr;
  vec_rsc_0_16_d <= vec_rsc_0_16_i_d;
  vec_rsc_0_16_wadr <= vec_rsc_0_16_i_wadr;
  vec_rsc_0_16_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_16_i_q_d <= vec_rsc_0_16_i_q_d_1;
  vec_rsc_0_16_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_16_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_17_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_17_i_q,
      radr => vec_rsc_0_17_i_radr,
      we => vec_rsc_0_17_we,
      d => vec_rsc_0_17_i_d,
      wadr => vec_rsc_0_17_i_wadr,
      d_d => vec_rsc_0_17_i_d_d,
      q_d => vec_rsc_0_17_i_q_d_1,
      radr_d => vec_rsc_0_17_i_radr_d,
      wadr_d => vec_rsc_0_17_i_wadr_d,
      we_d => vec_rsc_0_17_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_17_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_17_i_q <= vec_rsc_0_17_q;
  vec_rsc_0_17_radr <= vec_rsc_0_17_i_radr;
  vec_rsc_0_17_d <= vec_rsc_0_17_i_d;
  vec_rsc_0_17_wadr <= vec_rsc_0_17_i_wadr;
  vec_rsc_0_17_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_17_i_q_d <= vec_rsc_0_17_i_q_d_1;
  vec_rsc_0_17_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_17_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_18_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_18_i_q,
      radr => vec_rsc_0_18_i_radr,
      we => vec_rsc_0_18_we,
      d => vec_rsc_0_18_i_d,
      wadr => vec_rsc_0_18_i_wadr,
      d_d => vec_rsc_0_18_i_d_d,
      q_d => vec_rsc_0_18_i_q_d_1,
      radr_d => vec_rsc_0_18_i_radr_d,
      wadr_d => vec_rsc_0_18_i_wadr_d,
      we_d => vec_rsc_0_18_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_18_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_18_i_q <= vec_rsc_0_18_q;
  vec_rsc_0_18_radr <= vec_rsc_0_18_i_radr;
  vec_rsc_0_18_d <= vec_rsc_0_18_i_d;
  vec_rsc_0_18_wadr <= vec_rsc_0_18_i_wadr;
  vec_rsc_0_18_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_18_i_q_d <= vec_rsc_0_18_i_q_d_1;
  vec_rsc_0_18_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_18_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_19_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_19_i_q,
      radr => vec_rsc_0_19_i_radr,
      we => vec_rsc_0_19_we,
      d => vec_rsc_0_19_i_d,
      wadr => vec_rsc_0_19_i_wadr,
      d_d => vec_rsc_0_19_i_d_d,
      q_d => vec_rsc_0_19_i_q_d_1,
      radr_d => vec_rsc_0_19_i_radr_d,
      wadr_d => vec_rsc_0_19_i_wadr_d,
      we_d => vec_rsc_0_19_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_19_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_19_i_q <= vec_rsc_0_19_q;
  vec_rsc_0_19_radr <= vec_rsc_0_19_i_radr;
  vec_rsc_0_19_d <= vec_rsc_0_19_i_d;
  vec_rsc_0_19_wadr <= vec_rsc_0_19_i_wadr;
  vec_rsc_0_19_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_19_i_q_d <= vec_rsc_0_19_i_q_d_1;
  vec_rsc_0_19_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_19_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_20_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_20_i_q,
      radr => vec_rsc_0_20_i_radr,
      we => vec_rsc_0_20_we,
      d => vec_rsc_0_20_i_d,
      wadr => vec_rsc_0_20_i_wadr,
      d_d => vec_rsc_0_20_i_d_d,
      q_d => vec_rsc_0_20_i_q_d_1,
      radr_d => vec_rsc_0_20_i_radr_d,
      wadr_d => vec_rsc_0_20_i_wadr_d,
      we_d => vec_rsc_0_20_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_20_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_20_i_q <= vec_rsc_0_20_q;
  vec_rsc_0_20_radr <= vec_rsc_0_20_i_radr;
  vec_rsc_0_20_d <= vec_rsc_0_20_i_d;
  vec_rsc_0_20_wadr <= vec_rsc_0_20_i_wadr;
  vec_rsc_0_20_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_20_i_q_d <= vec_rsc_0_20_i_q_d_1;
  vec_rsc_0_20_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_20_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_21_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_21_i_q,
      radr => vec_rsc_0_21_i_radr,
      we => vec_rsc_0_21_we,
      d => vec_rsc_0_21_i_d,
      wadr => vec_rsc_0_21_i_wadr,
      d_d => vec_rsc_0_21_i_d_d,
      q_d => vec_rsc_0_21_i_q_d_1,
      radr_d => vec_rsc_0_21_i_radr_d,
      wadr_d => vec_rsc_0_21_i_wadr_d,
      we_d => vec_rsc_0_21_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_21_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_21_i_q <= vec_rsc_0_21_q;
  vec_rsc_0_21_radr <= vec_rsc_0_21_i_radr;
  vec_rsc_0_21_d <= vec_rsc_0_21_i_d;
  vec_rsc_0_21_wadr <= vec_rsc_0_21_i_wadr;
  vec_rsc_0_21_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_21_i_q_d <= vec_rsc_0_21_i_q_d_1;
  vec_rsc_0_21_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_21_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_22_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_22_i_q,
      radr => vec_rsc_0_22_i_radr,
      we => vec_rsc_0_22_we,
      d => vec_rsc_0_22_i_d,
      wadr => vec_rsc_0_22_i_wadr,
      d_d => vec_rsc_0_22_i_d_d,
      q_d => vec_rsc_0_22_i_q_d_1,
      radr_d => vec_rsc_0_22_i_radr_d,
      wadr_d => vec_rsc_0_22_i_wadr_d,
      we_d => vec_rsc_0_22_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_22_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_22_i_q <= vec_rsc_0_22_q;
  vec_rsc_0_22_radr <= vec_rsc_0_22_i_radr;
  vec_rsc_0_22_d <= vec_rsc_0_22_i_d;
  vec_rsc_0_22_wadr <= vec_rsc_0_22_i_wadr;
  vec_rsc_0_22_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_22_i_q_d <= vec_rsc_0_22_i_q_d_1;
  vec_rsc_0_22_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_22_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_23_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_23_i_q,
      radr => vec_rsc_0_23_i_radr,
      we => vec_rsc_0_23_we,
      d => vec_rsc_0_23_i_d,
      wadr => vec_rsc_0_23_i_wadr,
      d_d => vec_rsc_0_23_i_d_d,
      q_d => vec_rsc_0_23_i_q_d_1,
      radr_d => vec_rsc_0_23_i_radr_d,
      wadr_d => vec_rsc_0_23_i_wadr_d,
      we_d => vec_rsc_0_23_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_23_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_23_i_q <= vec_rsc_0_23_q;
  vec_rsc_0_23_radr <= vec_rsc_0_23_i_radr;
  vec_rsc_0_23_d <= vec_rsc_0_23_i_d;
  vec_rsc_0_23_wadr <= vec_rsc_0_23_i_wadr;
  vec_rsc_0_23_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_23_i_q_d <= vec_rsc_0_23_i_q_d_1;
  vec_rsc_0_23_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_23_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_24_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_24_i_q,
      radr => vec_rsc_0_24_i_radr,
      we => vec_rsc_0_24_we,
      d => vec_rsc_0_24_i_d,
      wadr => vec_rsc_0_24_i_wadr,
      d_d => vec_rsc_0_24_i_d_d,
      q_d => vec_rsc_0_24_i_q_d_1,
      radr_d => vec_rsc_0_24_i_radr_d,
      wadr_d => vec_rsc_0_24_i_wadr_d,
      we_d => vec_rsc_0_24_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_24_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_24_i_q <= vec_rsc_0_24_q;
  vec_rsc_0_24_radr <= vec_rsc_0_24_i_radr;
  vec_rsc_0_24_d <= vec_rsc_0_24_i_d;
  vec_rsc_0_24_wadr <= vec_rsc_0_24_i_wadr;
  vec_rsc_0_24_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_24_i_q_d <= vec_rsc_0_24_i_q_d_1;
  vec_rsc_0_24_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_24_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_25_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_25_i_q,
      radr => vec_rsc_0_25_i_radr,
      we => vec_rsc_0_25_we,
      d => vec_rsc_0_25_i_d,
      wadr => vec_rsc_0_25_i_wadr,
      d_d => vec_rsc_0_25_i_d_d,
      q_d => vec_rsc_0_25_i_q_d_1,
      radr_d => vec_rsc_0_25_i_radr_d,
      wadr_d => vec_rsc_0_25_i_wadr_d,
      we_d => vec_rsc_0_25_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_25_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_25_i_q <= vec_rsc_0_25_q;
  vec_rsc_0_25_radr <= vec_rsc_0_25_i_radr;
  vec_rsc_0_25_d <= vec_rsc_0_25_i_d;
  vec_rsc_0_25_wadr <= vec_rsc_0_25_i_wadr;
  vec_rsc_0_25_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_25_i_q_d <= vec_rsc_0_25_i_q_d_1;
  vec_rsc_0_25_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_25_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_26_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_26_i_q,
      radr => vec_rsc_0_26_i_radr,
      we => vec_rsc_0_26_we,
      d => vec_rsc_0_26_i_d,
      wadr => vec_rsc_0_26_i_wadr,
      d_d => vec_rsc_0_26_i_d_d,
      q_d => vec_rsc_0_26_i_q_d_1,
      radr_d => vec_rsc_0_26_i_radr_d,
      wadr_d => vec_rsc_0_26_i_wadr_d,
      we_d => vec_rsc_0_26_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_26_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_26_i_q <= vec_rsc_0_26_q;
  vec_rsc_0_26_radr <= vec_rsc_0_26_i_radr;
  vec_rsc_0_26_d <= vec_rsc_0_26_i_d;
  vec_rsc_0_26_wadr <= vec_rsc_0_26_i_wadr;
  vec_rsc_0_26_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_26_i_q_d <= vec_rsc_0_26_i_q_d_1;
  vec_rsc_0_26_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_26_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_27_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_27_i_q,
      radr => vec_rsc_0_27_i_radr,
      we => vec_rsc_0_27_we,
      d => vec_rsc_0_27_i_d,
      wadr => vec_rsc_0_27_i_wadr,
      d_d => vec_rsc_0_27_i_d_d,
      q_d => vec_rsc_0_27_i_q_d_1,
      radr_d => vec_rsc_0_27_i_radr_d,
      wadr_d => vec_rsc_0_27_i_wadr_d,
      we_d => vec_rsc_0_27_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_27_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_27_i_q <= vec_rsc_0_27_q;
  vec_rsc_0_27_radr <= vec_rsc_0_27_i_radr;
  vec_rsc_0_27_d <= vec_rsc_0_27_i_d;
  vec_rsc_0_27_wadr <= vec_rsc_0_27_i_wadr;
  vec_rsc_0_27_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_27_i_q_d <= vec_rsc_0_27_i_q_d_1;
  vec_rsc_0_27_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_27_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_28_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_28_i_q,
      radr => vec_rsc_0_28_i_radr,
      we => vec_rsc_0_28_we,
      d => vec_rsc_0_28_i_d,
      wadr => vec_rsc_0_28_i_wadr,
      d_d => vec_rsc_0_28_i_d_d,
      q_d => vec_rsc_0_28_i_q_d_1,
      radr_d => vec_rsc_0_28_i_radr_d,
      wadr_d => vec_rsc_0_28_i_wadr_d,
      we_d => vec_rsc_0_28_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_28_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_28_i_q <= vec_rsc_0_28_q;
  vec_rsc_0_28_radr <= vec_rsc_0_28_i_radr;
  vec_rsc_0_28_d <= vec_rsc_0_28_i_d;
  vec_rsc_0_28_wadr <= vec_rsc_0_28_i_wadr;
  vec_rsc_0_28_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_28_i_q_d <= vec_rsc_0_28_i_q_d_1;
  vec_rsc_0_28_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_28_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_29_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_29_i_q,
      radr => vec_rsc_0_29_i_radr,
      we => vec_rsc_0_29_we,
      d => vec_rsc_0_29_i_d,
      wadr => vec_rsc_0_29_i_wadr,
      d_d => vec_rsc_0_29_i_d_d,
      q_d => vec_rsc_0_29_i_q_d_1,
      radr_d => vec_rsc_0_29_i_radr_d,
      wadr_d => vec_rsc_0_29_i_wadr_d,
      we_d => vec_rsc_0_29_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_29_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_29_i_q <= vec_rsc_0_29_q;
  vec_rsc_0_29_radr <= vec_rsc_0_29_i_radr;
  vec_rsc_0_29_d <= vec_rsc_0_29_i_d;
  vec_rsc_0_29_wadr <= vec_rsc_0_29_i_wadr;
  vec_rsc_0_29_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_29_i_q_d <= vec_rsc_0_29_i_q_d_1;
  vec_rsc_0_29_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_29_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_30_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_30_i_q,
      radr => vec_rsc_0_30_i_radr,
      we => vec_rsc_0_30_we,
      d => vec_rsc_0_30_i_d,
      wadr => vec_rsc_0_30_i_wadr,
      d_d => vec_rsc_0_30_i_d_d,
      q_d => vec_rsc_0_30_i_q_d_1,
      radr_d => vec_rsc_0_30_i_radr_d,
      wadr_d => vec_rsc_0_30_i_wadr_d,
      we_d => vec_rsc_0_30_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_30_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_30_i_q <= vec_rsc_0_30_q;
  vec_rsc_0_30_radr <= vec_rsc_0_30_i_radr;
  vec_rsc_0_30_d <= vec_rsc_0_30_i_d;
  vec_rsc_0_30_wadr <= vec_rsc_0_30_i_wadr;
  vec_rsc_0_30_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_30_i_q_d <= vec_rsc_0_30_i_q_d_1;
  vec_rsc_0_30_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_30_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_31_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_31_i_q,
      radr => vec_rsc_0_31_i_radr,
      we => vec_rsc_0_31_we,
      d => vec_rsc_0_31_i_d,
      wadr => vec_rsc_0_31_i_wadr,
      d_d => vec_rsc_0_31_i_d_d,
      q_d => vec_rsc_0_31_i_q_d_1,
      radr_d => vec_rsc_0_31_i_radr_d,
      wadr_d => vec_rsc_0_31_i_wadr_d,
      we_d => vec_rsc_0_31_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_31_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_31_i_q <= vec_rsc_0_31_q;
  vec_rsc_0_31_radr <= vec_rsc_0_31_i_radr;
  vec_rsc_0_31_d <= vec_rsc_0_31_i_d;
  vec_rsc_0_31_wadr <= vec_rsc_0_31_i_wadr;
  vec_rsc_0_31_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_31_i_q_d <= vec_rsc_0_31_i_q_d_1;
  vec_rsc_0_31_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_31_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_32_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_32_i_q,
      radr => vec_rsc_0_32_i_radr,
      we => vec_rsc_0_32_we,
      d => vec_rsc_0_32_i_d,
      wadr => vec_rsc_0_32_i_wadr,
      d_d => vec_rsc_0_32_i_d_d,
      q_d => vec_rsc_0_32_i_q_d_1,
      radr_d => vec_rsc_0_32_i_radr_d,
      wadr_d => vec_rsc_0_32_i_wadr_d,
      we_d => vec_rsc_0_32_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_32_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_32_i_q <= vec_rsc_0_32_q;
  vec_rsc_0_32_radr <= vec_rsc_0_32_i_radr;
  vec_rsc_0_32_d <= vec_rsc_0_32_i_d;
  vec_rsc_0_32_wadr <= vec_rsc_0_32_i_wadr;
  vec_rsc_0_32_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_32_i_q_d <= vec_rsc_0_32_i_q_d_1;
  vec_rsc_0_32_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_32_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_33_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_33_i_q,
      radr => vec_rsc_0_33_i_radr,
      we => vec_rsc_0_33_we,
      d => vec_rsc_0_33_i_d,
      wadr => vec_rsc_0_33_i_wadr,
      d_d => vec_rsc_0_33_i_d_d,
      q_d => vec_rsc_0_33_i_q_d_1,
      radr_d => vec_rsc_0_33_i_radr_d,
      wadr_d => vec_rsc_0_33_i_wadr_d,
      we_d => vec_rsc_0_33_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_33_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_33_i_q <= vec_rsc_0_33_q;
  vec_rsc_0_33_radr <= vec_rsc_0_33_i_radr;
  vec_rsc_0_33_d <= vec_rsc_0_33_i_d;
  vec_rsc_0_33_wadr <= vec_rsc_0_33_i_wadr;
  vec_rsc_0_33_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_33_i_q_d <= vec_rsc_0_33_i_q_d_1;
  vec_rsc_0_33_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_33_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_34_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_34_i_q,
      radr => vec_rsc_0_34_i_radr,
      we => vec_rsc_0_34_we,
      d => vec_rsc_0_34_i_d,
      wadr => vec_rsc_0_34_i_wadr,
      d_d => vec_rsc_0_34_i_d_d,
      q_d => vec_rsc_0_34_i_q_d_1,
      radr_d => vec_rsc_0_34_i_radr_d,
      wadr_d => vec_rsc_0_34_i_wadr_d,
      we_d => vec_rsc_0_34_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_34_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_34_i_q <= vec_rsc_0_34_q;
  vec_rsc_0_34_radr <= vec_rsc_0_34_i_radr;
  vec_rsc_0_34_d <= vec_rsc_0_34_i_d;
  vec_rsc_0_34_wadr <= vec_rsc_0_34_i_wadr;
  vec_rsc_0_34_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_34_i_q_d <= vec_rsc_0_34_i_q_d_1;
  vec_rsc_0_34_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_34_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_35_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_35_i_q,
      radr => vec_rsc_0_35_i_radr,
      we => vec_rsc_0_35_we,
      d => vec_rsc_0_35_i_d,
      wadr => vec_rsc_0_35_i_wadr,
      d_d => vec_rsc_0_35_i_d_d,
      q_d => vec_rsc_0_35_i_q_d_1,
      radr_d => vec_rsc_0_35_i_radr_d,
      wadr_d => vec_rsc_0_35_i_wadr_d,
      we_d => vec_rsc_0_35_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_35_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_35_i_q <= vec_rsc_0_35_q;
  vec_rsc_0_35_radr <= vec_rsc_0_35_i_radr;
  vec_rsc_0_35_d <= vec_rsc_0_35_i_d;
  vec_rsc_0_35_wadr <= vec_rsc_0_35_i_wadr;
  vec_rsc_0_35_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_35_i_q_d <= vec_rsc_0_35_i_q_d_1;
  vec_rsc_0_35_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_35_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_36_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_36_i_q,
      radr => vec_rsc_0_36_i_radr,
      we => vec_rsc_0_36_we,
      d => vec_rsc_0_36_i_d,
      wadr => vec_rsc_0_36_i_wadr,
      d_d => vec_rsc_0_36_i_d_d,
      q_d => vec_rsc_0_36_i_q_d_1,
      radr_d => vec_rsc_0_36_i_radr_d,
      wadr_d => vec_rsc_0_36_i_wadr_d,
      we_d => vec_rsc_0_36_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_36_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_36_i_q <= vec_rsc_0_36_q;
  vec_rsc_0_36_radr <= vec_rsc_0_36_i_radr;
  vec_rsc_0_36_d <= vec_rsc_0_36_i_d;
  vec_rsc_0_36_wadr <= vec_rsc_0_36_i_wadr;
  vec_rsc_0_36_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_36_i_q_d <= vec_rsc_0_36_i_q_d_1;
  vec_rsc_0_36_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_36_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_37_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_37_i_q,
      radr => vec_rsc_0_37_i_radr,
      we => vec_rsc_0_37_we,
      d => vec_rsc_0_37_i_d,
      wadr => vec_rsc_0_37_i_wadr,
      d_d => vec_rsc_0_37_i_d_d,
      q_d => vec_rsc_0_37_i_q_d_1,
      radr_d => vec_rsc_0_37_i_radr_d,
      wadr_d => vec_rsc_0_37_i_wadr_d,
      we_d => vec_rsc_0_37_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_37_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_37_i_q <= vec_rsc_0_37_q;
  vec_rsc_0_37_radr <= vec_rsc_0_37_i_radr;
  vec_rsc_0_37_d <= vec_rsc_0_37_i_d;
  vec_rsc_0_37_wadr <= vec_rsc_0_37_i_wadr;
  vec_rsc_0_37_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_37_i_q_d <= vec_rsc_0_37_i_q_d_1;
  vec_rsc_0_37_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_37_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_38_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_38_i_q,
      radr => vec_rsc_0_38_i_radr,
      we => vec_rsc_0_38_we,
      d => vec_rsc_0_38_i_d,
      wadr => vec_rsc_0_38_i_wadr,
      d_d => vec_rsc_0_38_i_d_d,
      q_d => vec_rsc_0_38_i_q_d_1,
      radr_d => vec_rsc_0_38_i_radr_d,
      wadr_d => vec_rsc_0_38_i_wadr_d,
      we_d => vec_rsc_0_38_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_38_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_38_i_q <= vec_rsc_0_38_q;
  vec_rsc_0_38_radr <= vec_rsc_0_38_i_radr;
  vec_rsc_0_38_d <= vec_rsc_0_38_i_d;
  vec_rsc_0_38_wadr <= vec_rsc_0_38_i_wadr;
  vec_rsc_0_38_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_38_i_q_d <= vec_rsc_0_38_i_q_d_1;
  vec_rsc_0_38_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_38_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_39_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_39_i_q,
      radr => vec_rsc_0_39_i_radr,
      we => vec_rsc_0_39_we,
      d => vec_rsc_0_39_i_d,
      wadr => vec_rsc_0_39_i_wadr,
      d_d => vec_rsc_0_39_i_d_d,
      q_d => vec_rsc_0_39_i_q_d_1,
      radr_d => vec_rsc_0_39_i_radr_d,
      wadr_d => vec_rsc_0_39_i_wadr_d,
      we_d => vec_rsc_0_39_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_39_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_39_i_q <= vec_rsc_0_39_q;
  vec_rsc_0_39_radr <= vec_rsc_0_39_i_radr;
  vec_rsc_0_39_d <= vec_rsc_0_39_i_d;
  vec_rsc_0_39_wadr <= vec_rsc_0_39_i_wadr;
  vec_rsc_0_39_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_39_i_q_d <= vec_rsc_0_39_i_q_d_1;
  vec_rsc_0_39_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_39_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_40_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_40_i_q,
      radr => vec_rsc_0_40_i_radr,
      we => vec_rsc_0_40_we,
      d => vec_rsc_0_40_i_d,
      wadr => vec_rsc_0_40_i_wadr,
      d_d => vec_rsc_0_40_i_d_d,
      q_d => vec_rsc_0_40_i_q_d_1,
      radr_d => vec_rsc_0_40_i_radr_d,
      wadr_d => vec_rsc_0_40_i_wadr_d,
      we_d => vec_rsc_0_40_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_40_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_40_i_q <= vec_rsc_0_40_q;
  vec_rsc_0_40_radr <= vec_rsc_0_40_i_radr;
  vec_rsc_0_40_d <= vec_rsc_0_40_i_d;
  vec_rsc_0_40_wadr <= vec_rsc_0_40_i_wadr;
  vec_rsc_0_40_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_40_i_q_d <= vec_rsc_0_40_i_q_d_1;
  vec_rsc_0_40_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_40_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_41_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_41_i_q,
      radr => vec_rsc_0_41_i_radr,
      we => vec_rsc_0_41_we,
      d => vec_rsc_0_41_i_d,
      wadr => vec_rsc_0_41_i_wadr,
      d_d => vec_rsc_0_41_i_d_d,
      q_d => vec_rsc_0_41_i_q_d_1,
      radr_d => vec_rsc_0_41_i_radr_d,
      wadr_d => vec_rsc_0_41_i_wadr_d,
      we_d => vec_rsc_0_41_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_41_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_41_i_q <= vec_rsc_0_41_q;
  vec_rsc_0_41_radr <= vec_rsc_0_41_i_radr;
  vec_rsc_0_41_d <= vec_rsc_0_41_i_d;
  vec_rsc_0_41_wadr <= vec_rsc_0_41_i_wadr;
  vec_rsc_0_41_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_41_i_q_d <= vec_rsc_0_41_i_q_d_1;
  vec_rsc_0_41_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_41_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_42_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_42_i_q,
      radr => vec_rsc_0_42_i_radr,
      we => vec_rsc_0_42_we,
      d => vec_rsc_0_42_i_d,
      wadr => vec_rsc_0_42_i_wadr,
      d_d => vec_rsc_0_42_i_d_d,
      q_d => vec_rsc_0_42_i_q_d_1,
      radr_d => vec_rsc_0_42_i_radr_d,
      wadr_d => vec_rsc_0_42_i_wadr_d,
      we_d => vec_rsc_0_42_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_42_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_42_i_q <= vec_rsc_0_42_q;
  vec_rsc_0_42_radr <= vec_rsc_0_42_i_radr;
  vec_rsc_0_42_d <= vec_rsc_0_42_i_d;
  vec_rsc_0_42_wadr <= vec_rsc_0_42_i_wadr;
  vec_rsc_0_42_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_42_i_q_d <= vec_rsc_0_42_i_q_d_1;
  vec_rsc_0_42_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_42_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_43_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_43_i_q,
      radr => vec_rsc_0_43_i_radr,
      we => vec_rsc_0_43_we,
      d => vec_rsc_0_43_i_d,
      wadr => vec_rsc_0_43_i_wadr,
      d_d => vec_rsc_0_43_i_d_d,
      q_d => vec_rsc_0_43_i_q_d_1,
      radr_d => vec_rsc_0_43_i_radr_d,
      wadr_d => vec_rsc_0_43_i_wadr_d,
      we_d => vec_rsc_0_43_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_43_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_43_i_q <= vec_rsc_0_43_q;
  vec_rsc_0_43_radr <= vec_rsc_0_43_i_radr;
  vec_rsc_0_43_d <= vec_rsc_0_43_i_d;
  vec_rsc_0_43_wadr <= vec_rsc_0_43_i_wadr;
  vec_rsc_0_43_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_43_i_q_d <= vec_rsc_0_43_i_q_d_1;
  vec_rsc_0_43_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_43_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_44_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_44_i_q,
      radr => vec_rsc_0_44_i_radr,
      we => vec_rsc_0_44_we,
      d => vec_rsc_0_44_i_d,
      wadr => vec_rsc_0_44_i_wadr,
      d_d => vec_rsc_0_44_i_d_d,
      q_d => vec_rsc_0_44_i_q_d_1,
      radr_d => vec_rsc_0_44_i_radr_d,
      wadr_d => vec_rsc_0_44_i_wadr_d,
      we_d => vec_rsc_0_44_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_44_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_44_i_q <= vec_rsc_0_44_q;
  vec_rsc_0_44_radr <= vec_rsc_0_44_i_radr;
  vec_rsc_0_44_d <= vec_rsc_0_44_i_d;
  vec_rsc_0_44_wadr <= vec_rsc_0_44_i_wadr;
  vec_rsc_0_44_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_44_i_q_d <= vec_rsc_0_44_i_q_d_1;
  vec_rsc_0_44_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_44_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_45_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_45_i_q,
      radr => vec_rsc_0_45_i_radr,
      we => vec_rsc_0_45_we,
      d => vec_rsc_0_45_i_d,
      wadr => vec_rsc_0_45_i_wadr,
      d_d => vec_rsc_0_45_i_d_d,
      q_d => vec_rsc_0_45_i_q_d_1,
      radr_d => vec_rsc_0_45_i_radr_d,
      wadr_d => vec_rsc_0_45_i_wadr_d,
      we_d => vec_rsc_0_45_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_45_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_45_i_q <= vec_rsc_0_45_q;
  vec_rsc_0_45_radr <= vec_rsc_0_45_i_radr;
  vec_rsc_0_45_d <= vec_rsc_0_45_i_d;
  vec_rsc_0_45_wadr <= vec_rsc_0_45_i_wadr;
  vec_rsc_0_45_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_45_i_q_d <= vec_rsc_0_45_i_q_d_1;
  vec_rsc_0_45_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_45_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_46_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_46_i_q,
      radr => vec_rsc_0_46_i_radr,
      we => vec_rsc_0_46_we,
      d => vec_rsc_0_46_i_d,
      wadr => vec_rsc_0_46_i_wadr,
      d_d => vec_rsc_0_46_i_d_d,
      q_d => vec_rsc_0_46_i_q_d_1,
      radr_d => vec_rsc_0_46_i_radr_d,
      wadr_d => vec_rsc_0_46_i_wadr_d,
      we_d => vec_rsc_0_46_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_46_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_46_i_q <= vec_rsc_0_46_q;
  vec_rsc_0_46_radr <= vec_rsc_0_46_i_radr;
  vec_rsc_0_46_d <= vec_rsc_0_46_i_d;
  vec_rsc_0_46_wadr <= vec_rsc_0_46_i_wadr;
  vec_rsc_0_46_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_46_i_q_d <= vec_rsc_0_46_i_q_d_1;
  vec_rsc_0_46_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_46_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_47_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_47_i_q,
      radr => vec_rsc_0_47_i_radr,
      we => vec_rsc_0_47_we,
      d => vec_rsc_0_47_i_d,
      wadr => vec_rsc_0_47_i_wadr,
      d_d => vec_rsc_0_47_i_d_d,
      q_d => vec_rsc_0_47_i_q_d_1,
      radr_d => vec_rsc_0_47_i_radr_d,
      wadr_d => vec_rsc_0_47_i_wadr_d,
      we_d => vec_rsc_0_47_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_47_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_47_i_q <= vec_rsc_0_47_q;
  vec_rsc_0_47_radr <= vec_rsc_0_47_i_radr;
  vec_rsc_0_47_d <= vec_rsc_0_47_i_d;
  vec_rsc_0_47_wadr <= vec_rsc_0_47_i_wadr;
  vec_rsc_0_47_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_47_i_q_d <= vec_rsc_0_47_i_q_d_1;
  vec_rsc_0_47_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_47_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_48_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_48_i_q,
      radr => vec_rsc_0_48_i_radr,
      we => vec_rsc_0_48_we,
      d => vec_rsc_0_48_i_d,
      wadr => vec_rsc_0_48_i_wadr,
      d_d => vec_rsc_0_48_i_d_d,
      q_d => vec_rsc_0_48_i_q_d_1,
      radr_d => vec_rsc_0_48_i_radr_d,
      wadr_d => vec_rsc_0_48_i_wadr_d,
      we_d => vec_rsc_0_48_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_48_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_48_i_q <= vec_rsc_0_48_q;
  vec_rsc_0_48_radr <= vec_rsc_0_48_i_radr;
  vec_rsc_0_48_d <= vec_rsc_0_48_i_d;
  vec_rsc_0_48_wadr <= vec_rsc_0_48_i_wadr;
  vec_rsc_0_48_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_48_i_q_d <= vec_rsc_0_48_i_q_d_1;
  vec_rsc_0_48_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_48_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_49_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_49_i_q,
      radr => vec_rsc_0_49_i_radr,
      we => vec_rsc_0_49_we,
      d => vec_rsc_0_49_i_d,
      wadr => vec_rsc_0_49_i_wadr,
      d_d => vec_rsc_0_49_i_d_d,
      q_d => vec_rsc_0_49_i_q_d_1,
      radr_d => vec_rsc_0_49_i_radr_d,
      wadr_d => vec_rsc_0_49_i_wadr_d,
      we_d => vec_rsc_0_49_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_49_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_49_i_q <= vec_rsc_0_49_q;
  vec_rsc_0_49_radr <= vec_rsc_0_49_i_radr;
  vec_rsc_0_49_d <= vec_rsc_0_49_i_d;
  vec_rsc_0_49_wadr <= vec_rsc_0_49_i_wadr;
  vec_rsc_0_49_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_49_i_q_d <= vec_rsc_0_49_i_q_d_1;
  vec_rsc_0_49_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_49_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_50_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_50_i_q,
      radr => vec_rsc_0_50_i_radr,
      we => vec_rsc_0_50_we,
      d => vec_rsc_0_50_i_d,
      wadr => vec_rsc_0_50_i_wadr,
      d_d => vec_rsc_0_50_i_d_d,
      q_d => vec_rsc_0_50_i_q_d_1,
      radr_d => vec_rsc_0_50_i_radr_d,
      wadr_d => vec_rsc_0_50_i_wadr_d,
      we_d => vec_rsc_0_50_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_50_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_50_i_q <= vec_rsc_0_50_q;
  vec_rsc_0_50_radr <= vec_rsc_0_50_i_radr;
  vec_rsc_0_50_d <= vec_rsc_0_50_i_d;
  vec_rsc_0_50_wadr <= vec_rsc_0_50_i_wadr;
  vec_rsc_0_50_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_50_i_q_d <= vec_rsc_0_50_i_q_d_1;
  vec_rsc_0_50_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_50_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_51_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_51_i_q,
      radr => vec_rsc_0_51_i_radr,
      we => vec_rsc_0_51_we,
      d => vec_rsc_0_51_i_d,
      wadr => vec_rsc_0_51_i_wadr,
      d_d => vec_rsc_0_51_i_d_d,
      q_d => vec_rsc_0_51_i_q_d_1,
      radr_d => vec_rsc_0_51_i_radr_d,
      wadr_d => vec_rsc_0_51_i_wadr_d,
      we_d => vec_rsc_0_51_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_51_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_51_i_q <= vec_rsc_0_51_q;
  vec_rsc_0_51_radr <= vec_rsc_0_51_i_radr;
  vec_rsc_0_51_d <= vec_rsc_0_51_i_d;
  vec_rsc_0_51_wadr <= vec_rsc_0_51_i_wadr;
  vec_rsc_0_51_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_51_i_q_d <= vec_rsc_0_51_i_q_d_1;
  vec_rsc_0_51_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_51_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_52_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_52_i_q,
      radr => vec_rsc_0_52_i_radr,
      we => vec_rsc_0_52_we,
      d => vec_rsc_0_52_i_d,
      wadr => vec_rsc_0_52_i_wadr,
      d_d => vec_rsc_0_52_i_d_d,
      q_d => vec_rsc_0_52_i_q_d_1,
      radr_d => vec_rsc_0_52_i_radr_d,
      wadr_d => vec_rsc_0_52_i_wadr_d,
      we_d => vec_rsc_0_52_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_52_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_52_i_q <= vec_rsc_0_52_q;
  vec_rsc_0_52_radr <= vec_rsc_0_52_i_radr;
  vec_rsc_0_52_d <= vec_rsc_0_52_i_d;
  vec_rsc_0_52_wadr <= vec_rsc_0_52_i_wadr;
  vec_rsc_0_52_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_52_i_q_d <= vec_rsc_0_52_i_q_d_1;
  vec_rsc_0_52_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_52_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_53_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_53_i_q,
      radr => vec_rsc_0_53_i_radr,
      we => vec_rsc_0_53_we,
      d => vec_rsc_0_53_i_d,
      wadr => vec_rsc_0_53_i_wadr,
      d_d => vec_rsc_0_53_i_d_d,
      q_d => vec_rsc_0_53_i_q_d_1,
      radr_d => vec_rsc_0_53_i_radr_d,
      wadr_d => vec_rsc_0_53_i_wadr_d,
      we_d => vec_rsc_0_53_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_53_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_53_i_q <= vec_rsc_0_53_q;
  vec_rsc_0_53_radr <= vec_rsc_0_53_i_radr;
  vec_rsc_0_53_d <= vec_rsc_0_53_i_d;
  vec_rsc_0_53_wadr <= vec_rsc_0_53_i_wadr;
  vec_rsc_0_53_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_53_i_q_d <= vec_rsc_0_53_i_q_d_1;
  vec_rsc_0_53_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_53_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_54_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_54_i_q,
      radr => vec_rsc_0_54_i_radr,
      we => vec_rsc_0_54_we,
      d => vec_rsc_0_54_i_d,
      wadr => vec_rsc_0_54_i_wadr,
      d_d => vec_rsc_0_54_i_d_d,
      q_d => vec_rsc_0_54_i_q_d_1,
      radr_d => vec_rsc_0_54_i_radr_d,
      wadr_d => vec_rsc_0_54_i_wadr_d,
      we_d => vec_rsc_0_54_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_54_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_54_i_q <= vec_rsc_0_54_q;
  vec_rsc_0_54_radr <= vec_rsc_0_54_i_radr;
  vec_rsc_0_54_d <= vec_rsc_0_54_i_d;
  vec_rsc_0_54_wadr <= vec_rsc_0_54_i_wadr;
  vec_rsc_0_54_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_54_i_q_d <= vec_rsc_0_54_i_q_d_1;
  vec_rsc_0_54_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_54_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_55_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_55_i_q,
      radr => vec_rsc_0_55_i_radr,
      we => vec_rsc_0_55_we,
      d => vec_rsc_0_55_i_d,
      wadr => vec_rsc_0_55_i_wadr,
      d_d => vec_rsc_0_55_i_d_d,
      q_d => vec_rsc_0_55_i_q_d_1,
      radr_d => vec_rsc_0_55_i_radr_d,
      wadr_d => vec_rsc_0_55_i_wadr_d,
      we_d => vec_rsc_0_55_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_55_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_55_i_q <= vec_rsc_0_55_q;
  vec_rsc_0_55_radr <= vec_rsc_0_55_i_radr;
  vec_rsc_0_55_d <= vec_rsc_0_55_i_d;
  vec_rsc_0_55_wadr <= vec_rsc_0_55_i_wadr;
  vec_rsc_0_55_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_55_i_q_d <= vec_rsc_0_55_i_q_d_1;
  vec_rsc_0_55_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_55_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_56_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_56_i_q,
      radr => vec_rsc_0_56_i_radr,
      we => vec_rsc_0_56_we,
      d => vec_rsc_0_56_i_d,
      wadr => vec_rsc_0_56_i_wadr,
      d_d => vec_rsc_0_56_i_d_d,
      q_d => vec_rsc_0_56_i_q_d_1,
      radr_d => vec_rsc_0_56_i_radr_d,
      wadr_d => vec_rsc_0_56_i_wadr_d,
      we_d => vec_rsc_0_56_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_56_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_56_i_q <= vec_rsc_0_56_q;
  vec_rsc_0_56_radr <= vec_rsc_0_56_i_radr;
  vec_rsc_0_56_d <= vec_rsc_0_56_i_d;
  vec_rsc_0_56_wadr <= vec_rsc_0_56_i_wadr;
  vec_rsc_0_56_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_56_i_q_d <= vec_rsc_0_56_i_q_d_1;
  vec_rsc_0_56_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_56_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_57_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_57_i_q,
      radr => vec_rsc_0_57_i_radr,
      we => vec_rsc_0_57_we,
      d => vec_rsc_0_57_i_d,
      wadr => vec_rsc_0_57_i_wadr,
      d_d => vec_rsc_0_57_i_d_d,
      q_d => vec_rsc_0_57_i_q_d_1,
      radr_d => vec_rsc_0_57_i_radr_d,
      wadr_d => vec_rsc_0_57_i_wadr_d,
      we_d => vec_rsc_0_57_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_57_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_57_i_q <= vec_rsc_0_57_q;
  vec_rsc_0_57_radr <= vec_rsc_0_57_i_radr;
  vec_rsc_0_57_d <= vec_rsc_0_57_i_d;
  vec_rsc_0_57_wadr <= vec_rsc_0_57_i_wadr;
  vec_rsc_0_57_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_57_i_q_d <= vec_rsc_0_57_i_q_d_1;
  vec_rsc_0_57_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_57_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_58_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_58_i_q,
      radr => vec_rsc_0_58_i_radr,
      we => vec_rsc_0_58_we,
      d => vec_rsc_0_58_i_d,
      wadr => vec_rsc_0_58_i_wadr,
      d_d => vec_rsc_0_58_i_d_d,
      q_d => vec_rsc_0_58_i_q_d_1,
      radr_d => vec_rsc_0_58_i_radr_d,
      wadr_d => vec_rsc_0_58_i_wadr_d,
      we_d => vec_rsc_0_58_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_58_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_58_i_q <= vec_rsc_0_58_q;
  vec_rsc_0_58_radr <= vec_rsc_0_58_i_radr;
  vec_rsc_0_58_d <= vec_rsc_0_58_i_d;
  vec_rsc_0_58_wadr <= vec_rsc_0_58_i_wadr;
  vec_rsc_0_58_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_58_i_q_d <= vec_rsc_0_58_i_q_d_1;
  vec_rsc_0_58_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_58_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_59_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_59_i_q,
      radr => vec_rsc_0_59_i_radr,
      we => vec_rsc_0_59_we,
      d => vec_rsc_0_59_i_d,
      wadr => vec_rsc_0_59_i_wadr,
      d_d => vec_rsc_0_59_i_d_d,
      q_d => vec_rsc_0_59_i_q_d_1,
      radr_d => vec_rsc_0_59_i_radr_d,
      wadr_d => vec_rsc_0_59_i_wadr_d,
      we_d => vec_rsc_0_59_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_59_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_59_i_q <= vec_rsc_0_59_q;
  vec_rsc_0_59_radr <= vec_rsc_0_59_i_radr;
  vec_rsc_0_59_d <= vec_rsc_0_59_i_d;
  vec_rsc_0_59_wadr <= vec_rsc_0_59_i_wadr;
  vec_rsc_0_59_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_59_i_q_d <= vec_rsc_0_59_i_q_d_1;
  vec_rsc_0_59_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_59_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_60_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_60_i_q,
      radr => vec_rsc_0_60_i_radr,
      we => vec_rsc_0_60_we,
      d => vec_rsc_0_60_i_d,
      wadr => vec_rsc_0_60_i_wadr,
      d_d => vec_rsc_0_60_i_d_d,
      q_d => vec_rsc_0_60_i_q_d_1,
      radr_d => vec_rsc_0_60_i_radr_d,
      wadr_d => vec_rsc_0_60_i_wadr_d,
      we_d => vec_rsc_0_60_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_60_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_60_i_q <= vec_rsc_0_60_q;
  vec_rsc_0_60_radr <= vec_rsc_0_60_i_radr;
  vec_rsc_0_60_d <= vec_rsc_0_60_i_d;
  vec_rsc_0_60_wadr <= vec_rsc_0_60_i_wadr;
  vec_rsc_0_60_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_60_i_q_d <= vec_rsc_0_60_i_q_d_1;
  vec_rsc_0_60_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_60_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_61_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_61_i_q,
      radr => vec_rsc_0_61_i_radr,
      we => vec_rsc_0_61_we,
      d => vec_rsc_0_61_i_d,
      wadr => vec_rsc_0_61_i_wadr,
      d_d => vec_rsc_0_61_i_d_d,
      q_d => vec_rsc_0_61_i_q_d_1,
      radr_d => vec_rsc_0_61_i_radr_d,
      wadr_d => vec_rsc_0_61_i_wadr_d,
      we_d => vec_rsc_0_61_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_61_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_61_i_q <= vec_rsc_0_61_q;
  vec_rsc_0_61_radr <= vec_rsc_0_61_i_radr;
  vec_rsc_0_61_d <= vec_rsc_0_61_i_d;
  vec_rsc_0_61_wadr <= vec_rsc_0_61_i_wadr;
  vec_rsc_0_61_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_61_i_q_d <= vec_rsc_0_61_i_q_d_1;
  vec_rsc_0_61_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_61_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_62_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_62_i_q,
      radr => vec_rsc_0_62_i_radr,
      we => vec_rsc_0_62_we,
      d => vec_rsc_0_62_i_d,
      wadr => vec_rsc_0_62_i_wadr,
      d_d => vec_rsc_0_62_i_d_d,
      q_d => vec_rsc_0_62_i_q_d_1,
      radr_d => vec_rsc_0_62_i_radr_d,
      wadr_d => vec_rsc_0_62_i_wadr_d,
      we_d => vec_rsc_0_62_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_62_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_62_i_q <= vec_rsc_0_62_q;
  vec_rsc_0_62_radr <= vec_rsc_0_62_i_radr;
  vec_rsc_0_62_d <= vec_rsc_0_62_i_d;
  vec_rsc_0_62_wadr <= vec_rsc_0_62_i_wadr;
  vec_rsc_0_62_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_62_i_q_d <= vec_rsc_0_62_i_q_d_1;
  vec_rsc_0_62_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_62_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_63_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen
    PORT MAP(
      q => vec_rsc_0_63_i_q,
      radr => vec_rsc_0_63_i_radr,
      we => vec_rsc_0_63_we,
      d => vec_rsc_0_63_i_d,
      wadr => vec_rsc_0_63_i_wadr,
      d_d => vec_rsc_0_63_i_d_d,
      q_d => vec_rsc_0_63_i_q_d_1,
      radr_d => vec_rsc_0_63_i_radr_d,
      wadr_d => vec_rsc_0_63_i_wadr_d,
      we_d => vec_rsc_0_63_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_63_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_63_i_q <= vec_rsc_0_63_q;
  vec_rsc_0_63_radr <= vec_rsc_0_63_i_radr;
  vec_rsc_0_63_d <= vec_rsc_0_63_i_d;
  vec_rsc_0_63_wadr <= vec_rsc_0_63_i_wadr;
  vec_rsc_0_63_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_63_i_q_d <= vec_rsc_0_63_i_q_d_1;
  vec_rsc_0_63_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_63_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  twiddle_rsc_0_0_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_0_i_q,
      radr => twiddle_rsc_0_0_i_radr,
      q_d => twiddle_rsc_0_0_i_q_d_1,
      radr_d => twiddle_rsc_0_0_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_0_i_q <= twiddle_rsc_0_0_q;
  twiddle_rsc_0_0_radr <= twiddle_rsc_0_0_i_radr;
  twiddle_rsc_0_0_i_q_d <= twiddle_rsc_0_0_i_q_d_1;
  twiddle_rsc_0_0_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_1_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_1_i_q,
      radr => twiddle_rsc_0_1_i_radr,
      q_d => twiddle_rsc_0_1_i_q_d_1,
      radr_d => twiddle_rsc_0_1_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_1_i_q <= twiddle_rsc_0_1_q;
  twiddle_rsc_0_1_radr <= twiddle_rsc_0_1_i_radr;
  twiddle_rsc_0_1_i_q_d <= twiddle_rsc_0_1_i_q_d_1;
  twiddle_rsc_0_1_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_2_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_2_i_q,
      radr => twiddle_rsc_0_2_i_radr,
      q_d => twiddle_rsc_0_2_i_q_d_1,
      radr_d => twiddle_rsc_0_2_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_2_i_q <= twiddle_rsc_0_2_q;
  twiddle_rsc_0_2_radr <= twiddle_rsc_0_2_i_radr;
  twiddle_rsc_0_2_i_q_d <= twiddle_rsc_0_2_i_q_d_1;
  twiddle_rsc_0_2_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_3_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_3_i_q,
      radr => twiddle_rsc_0_3_i_radr,
      q_d => twiddle_rsc_0_3_i_q_d_1,
      radr_d => twiddle_rsc_0_3_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_3_i_q <= twiddle_rsc_0_3_q;
  twiddle_rsc_0_3_radr <= twiddle_rsc_0_3_i_radr;
  twiddle_rsc_0_3_i_q_d <= twiddle_rsc_0_3_i_q_d_1;
  twiddle_rsc_0_3_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_4_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_4_i_q,
      radr => twiddle_rsc_0_4_i_radr,
      q_d => twiddle_rsc_0_4_i_q_d_1,
      radr_d => twiddle_rsc_0_4_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_4_i_q <= twiddle_rsc_0_4_q;
  twiddle_rsc_0_4_radr <= twiddle_rsc_0_4_i_radr;
  twiddle_rsc_0_4_i_q_d <= twiddle_rsc_0_4_i_q_d_1;
  twiddle_rsc_0_4_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_5_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_5_i_q,
      radr => twiddle_rsc_0_5_i_radr,
      q_d => twiddle_rsc_0_5_i_q_d_1,
      radr_d => twiddle_rsc_0_5_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_5_i_q <= twiddle_rsc_0_5_q;
  twiddle_rsc_0_5_radr <= twiddle_rsc_0_5_i_radr;
  twiddle_rsc_0_5_i_q_d <= twiddle_rsc_0_5_i_q_d_1;
  twiddle_rsc_0_5_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_6_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_6_i_q,
      radr => twiddle_rsc_0_6_i_radr,
      q_d => twiddle_rsc_0_6_i_q_d_1,
      radr_d => twiddle_rsc_0_6_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_6_i_q <= twiddle_rsc_0_6_q;
  twiddle_rsc_0_6_radr <= twiddle_rsc_0_6_i_radr;
  twiddle_rsc_0_6_i_q_d <= twiddle_rsc_0_6_i_q_d_1;
  twiddle_rsc_0_6_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_7_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_7_i_q,
      radr => twiddle_rsc_0_7_i_radr,
      q_d => twiddle_rsc_0_7_i_q_d_1,
      radr_d => twiddle_rsc_0_7_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_7_i_q <= twiddle_rsc_0_7_q;
  twiddle_rsc_0_7_radr <= twiddle_rsc_0_7_i_radr;
  twiddle_rsc_0_7_i_q_d <= twiddle_rsc_0_7_i_q_d_1;
  twiddle_rsc_0_7_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_8_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_8_i_q,
      radr => twiddle_rsc_0_8_i_radr,
      q_d => twiddle_rsc_0_8_i_q_d_1,
      radr_d => twiddle_rsc_0_8_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_8_i_q <= twiddle_rsc_0_8_q;
  twiddle_rsc_0_8_radr <= twiddle_rsc_0_8_i_radr;
  twiddle_rsc_0_8_i_q_d <= twiddle_rsc_0_8_i_q_d_1;
  twiddle_rsc_0_8_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_9_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_9_i_q,
      radr => twiddle_rsc_0_9_i_radr,
      q_d => twiddle_rsc_0_9_i_q_d_1,
      radr_d => twiddle_rsc_0_9_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_9_i_q <= twiddle_rsc_0_9_q;
  twiddle_rsc_0_9_radr <= twiddle_rsc_0_9_i_radr;
  twiddle_rsc_0_9_i_q_d <= twiddle_rsc_0_9_i_q_d_1;
  twiddle_rsc_0_9_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_10_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_10_i_q,
      radr => twiddle_rsc_0_10_i_radr,
      q_d => twiddle_rsc_0_10_i_q_d_1,
      radr_d => twiddle_rsc_0_10_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_10_i_q <= twiddle_rsc_0_10_q;
  twiddle_rsc_0_10_radr <= twiddle_rsc_0_10_i_radr;
  twiddle_rsc_0_10_i_q_d <= twiddle_rsc_0_10_i_q_d_1;
  twiddle_rsc_0_10_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_11_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_11_i_q,
      radr => twiddle_rsc_0_11_i_radr,
      q_d => twiddle_rsc_0_11_i_q_d_1,
      radr_d => twiddle_rsc_0_11_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_11_i_q <= twiddle_rsc_0_11_q;
  twiddle_rsc_0_11_radr <= twiddle_rsc_0_11_i_radr;
  twiddle_rsc_0_11_i_q_d <= twiddle_rsc_0_11_i_q_d_1;
  twiddle_rsc_0_11_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_12_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_12_i_q,
      radr => twiddle_rsc_0_12_i_radr,
      q_d => twiddle_rsc_0_12_i_q_d_1,
      radr_d => twiddle_rsc_0_12_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_12_i_q <= twiddle_rsc_0_12_q;
  twiddle_rsc_0_12_radr <= twiddle_rsc_0_12_i_radr;
  twiddle_rsc_0_12_i_q_d <= twiddle_rsc_0_12_i_q_d_1;
  twiddle_rsc_0_12_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_13_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_13_i_q,
      radr => twiddle_rsc_0_13_i_radr,
      q_d => twiddle_rsc_0_13_i_q_d_1,
      radr_d => twiddle_rsc_0_13_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_13_i_q <= twiddle_rsc_0_13_q;
  twiddle_rsc_0_13_radr <= twiddle_rsc_0_13_i_radr;
  twiddle_rsc_0_13_i_q_d <= twiddle_rsc_0_13_i_q_d_1;
  twiddle_rsc_0_13_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_14_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_14_i_q,
      radr => twiddle_rsc_0_14_i_radr,
      q_d => twiddle_rsc_0_14_i_q_d_1,
      radr_d => twiddle_rsc_0_14_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_14_i_q <= twiddle_rsc_0_14_q;
  twiddle_rsc_0_14_radr <= twiddle_rsc_0_14_i_radr;
  twiddle_rsc_0_14_i_q_d <= twiddle_rsc_0_14_i_q_d_1;
  twiddle_rsc_0_14_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_15_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_15_i_q,
      radr => twiddle_rsc_0_15_i_radr,
      q_d => twiddle_rsc_0_15_i_q_d_1,
      radr_d => twiddle_rsc_0_15_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_15_i_q <= twiddle_rsc_0_15_q;
  twiddle_rsc_0_15_radr <= twiddle_rsc_0_15_i_radr;
  twiddle_rsc_0_15_i_q_d <= twiddle_rsc_0_15_i_q_d_1;
  twiddle_rsc_0_15_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_16_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_16_i_q,
      radr => twiddle_rsc_0_16_i_radr,
      q_d => twiddle_rsc_0_16_i_q_d_1,
      radr_d => twiddle_rsc_0_16_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_16_i_q <= twiddle_rsc_0_16_q;
  twiddle_rsc_0_16_radr <= twiddle_rsc_0_16_i_radr;
  twiddle_rsc_0_16_i_q_d <= twiddle_rsc_0_16_i_q_d_1;
  twiddle_rsc_0_16_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_17_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_17_i_q,
      radr => twiddle_rsc_0_17_i_radr,
      q_d => twiddle_rsc_0_17_i_q_d_1,
      radr_d => twiddle_rsc_0_17_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_17_i_q <= twiddle_rsc_0_17_q;
  twiddle_rsc_0_17_radr <= twiddle_rsc_0_17_i_radr;
  twiddle_rsc_0_17_i_q_d <= twiddle_rsc_0_17_i_q_d_1;
  twiddle_rsc_0_17_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_18_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_18_i_q,
      radr => twiddle_rsc_0_18_i_radr,
      q_d => twiddle_rsc_0_18_i_q_d_1,
      radr_d => twiddle_rsc_0_18_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_18_i_q <= twiddle_rsc_0_18_q;
  twiddle_rsc_0_18_radr <= twiddle_rsc_0_18_i_radr;
  twiddle_rsc_0_18_i_q_d <= twiddle_rsc_0_18_i_q_d_1;
  twiddle_rsc_0_18_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_19_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_19_i_q,
      radr => twiddle_rsc_0_19_i_radr,
      q_d => twiddle_rsc_0_19_i_q_d_1,
      radr_d => twiddle_rsc_0_19_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_19_i_q <= twiddle_rsc_0_19_q;
  twiddle_rsc_0_19_radr <= twiddle_rsc_0_19_i_radr;
  twiddle_rsc_0_19_i_q_d <= twiddle_rsc_0_19_i_q_d_1;
  twiddle_rsc_0_19_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_20_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_20_i_q,
      radr => twiddle_rsc_0_20_i_radr,
      q_d => twiddle_rsc_0_20_i_q_d_1,
      radr_d => twiddle_rsc_0_20_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_20_i_q <= twiddle_rsc_0_20_q;
  twiddle_rsc_0_20_radr <= twiddle_rsc_0_20_i_radr;
  twiddle_rsc_0_20_i_q_d <= twiddle_rsc_0_20_i_q_d_1;
  twiddle_rsc_0_20_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_21_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_21_i_q,
      radr => twiddle_rsc_0_21_i_radr,
      q_d => twiddle_rsc_0_21_i_q_d_1,
      radr_d => twiddle_rsc_0_21_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_21_i_q <= twiddle_rsc_0_21_q;
  twiddle_rsc_0_21_radr <= twiddle_rsc_0_21_i_radr;
  twiddle_rsc_0_21_i_q_d <= twiddle_rsc_0_21_i_q_d_1;
  twiddle_rsc_0_21_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_22_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_22_i_q,
      radr => twiddle_rsc_0_22_i_radr,
      q_d => twiddle_rsc_0_22_i_q_d_1,
      radr_d => twiddle_rsc_0_22_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_22_i_q <= twiddle_rsc_0_22_q;
  twiddle_rsc_0_22_radr <= twiddle_rsc_0_22_i_radr;
  twiddle_rsc_0_22_i_q_d <= twiddle_rsc_0_22_i_q_d_1;
  twiddle_rsc_0_22_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_23_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_23_i_q,
      radr => twiddle_rsc_0_23_i_radr,
      q_d => twiddle_rsc_0_23_i_q_d_1,
      radr_d => twiddle_rsc_0_23_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_23_i_q <= twiddle_rsc_0_23_q;
  twiddle_rsc_0_23_radr <= twiddle_rsc_0_23_i_radr;
  twiddle_rsc_0_23_i_q_d <= twiddle_rsc_0_23_i_q_d_1;
  twiddle_rsc_0_23_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_24_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_24_i_q,
      radr => twiddle_rsc_0_24_i_radr,
      q_d => twiddle_rsc_0_24_i_q_d_1,
      radr_d => twiddle_rsc_0_24_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_24_i_q <= twiddle_rsc_0_24_q;
  twiddle_rsc_0_24_radr <= twiddle_rsc_0_24_i_radr;
  twiddle_rsc_0_24_i_q_d <= twiddle_rsc_0_24_i_q_d_1;
  twiddle_rsc_0_24_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_25_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_25_i_q,
      radr => twiddle_rsc_0_25_i_radr,
      q_d => twiddle_rsc_0_25_i_q_d_1,
      radr_d => twiddle_rsc_0_25_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_25_i_q <= twiddle_rsc_0_25_q;
  twiddle_rsc_0_25_radr <= twiddle_rsc_0_25_i_radr;
  twiddle_rsc_0_25_i_q_d <= twiddle_rsc_0_25_i_q_d_1;
  twiddle_rsc_0_25_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_26_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_26_i_q,
      radr => twiddle_rsc_0_26_i_radr,
      q_d => twiddle_rsc_0_26_i_q_d_1,
      radr_d => twiddle_rsc_0_26_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_26_i_q <= twiddle_rsc_0_26_q;
  twiddle_rsc_0_26_radr <= twiddle_rsc_0_26_i_radr;
  twiddle_rsc_0_26_i_q_d <= twiddle_rsc_0_26_i_q_d_1;
  twiddle_rsc_0_26_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_27_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_27_i_q,
      radr => twiddle_rsc_0_27_i_radr,
      q_d => twiddle_rsc_0_27_i_q_d_1,
      radr_d => twiddle_rsc_0_27_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_27_i_q <= twiddle_rsc_0_27_q;
  twiddle_rsc_0_27_radr <= twiddle_rsc_0_27_i_radr;
  twiddle_rsc_0_27_i_q_d <= twiddle_rsc_0_27_i_q_d_1;
  twiddle_rsc_0_27_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_28_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_28_i_q,
      radr => twiddle_rsc_0_28_i_radr,
      q_d => twiddle_rsc_0_28_i_q_d_1,
      radr_d => twiddle_rsc_0_28_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_28_i_q <= twiddle_rsc_0_28_q;
  twiddle_rsc_0_28_radr <= twiddle_rsc_0_28_i_radr;
  twiddle_rsc_0_28_i_q_d <= twiddle_rsc_0_28_i_q_d_1;
  twiddle_rsc_0_28_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_29_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_29_i_q,
      radr => twiddle_rsc_0_29_i_radr,
      q_d => twiddle_rsc_0_29_i_q_d_1,
      radr_d => twiddle_rsc_0_29_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_29_i_q <= twiddle_rsc_0_29_q;
  twiddle_rsc_0_29_radr <= twiddle_rsc_0_29_i_radr;
  twiddle_rsc_0_29_i_q_d <= twiddle_rsc_0_29_i_q_d_1;
  twiddle_rsc_0_29_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_30_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_30_i_q,
      radr => twiddle_rsc_0_30_i_radr,
      q_d => twiddle_rsc_0_30_i_q_d_1,
      radr_d => twiddle_rsc_0_30_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_30_i_q <= twiddle_rsc_0_30_q;
  twiddle_rsc_0_30_radr <= twiddle_rsc_0_30_i_radr;
  twiddle_rsc_0_30_i_q_d <= twiddle_rsc_0_30_i_q_d_1;
  twiddle_rsc_0_30_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_31_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_31_i_q,
      radr => twiddle_rsc_0_31_i_radr,
      q_d => twiddle_rsc_0_31_i_q_d_1,
      radr_d => twiddle_rsc_0_31_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_31_i_q <= twiddle_rsc_0_31_q;
  twiddle_rsc_0_31_radr <= twiddle_rsc_0_31_i_radr;
  twiddle_rsc_0_31_i_q_d <= twiddle_rsc_0_31_i_q_d_1;
  twiddle_rsc_0_31_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_32_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_32_i_q,
      radr => twiddle_rsc_0_32_i_radr,
      q_d => twiddle_rsc_0_32_i_q_d_1,
      radr_d => twiddle_rsc_0_32_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_32_i_q <= twiddle_rsc_0_32_q;
  twiddle_rsc_0_32_radr <= twiddle_rsc_0_32_i_radr;
  twiddle_rsc_0_32_i_q_d <= twiddle_rsc_0_32_i_q_d_1;
  twiddle_rsc_0_32_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_33_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_33_i_q,
      radr => twiddle_rsc_0_33_i_radr,
      q_d => twiddle_rsc_0_33_i_q_d_1,
      radr_d => twiddle_rsc_0_33_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_33_i_q <= twiddle_rsc_0_33_q;
  twiddle_rsc_0_33_radr <= twiddle_rsc_0_33_i_radr;
  twiddle_rsc_0_33_i_q_d <= twiddle_rsc_0_33_i_q_d_1;
  twiddle_rsc_0_33_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_34_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_34_i_q,
      radr => twiddle_rsc_0_34_i_radr,
      q_d => twiddle_rsc_0_34_i_q_d_1,
      radr_d => twiddle_rsc_0_34_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_34_i_q <= twiddle_rsc_0_34_q;
  twiddle_rsc_0_34_radr <= twiddle_rsc_0_34_i_radr;
  twiddle_rsc_0_34_i_q_d <= twiddle_rsc_0_34_i_q_d_1;
  twiddle_rsc_0_34_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_35_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_35_i_q,
      radr => twiddle_rsc_0_35_i_radr,
      q_d => twiddle_rsc_0_35_i_q_d_1,
      radr_d => twiddle_rsc_0_35_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_35_i_q <= twiddle_rsc_0_35_q;
  twiddle_rsc_0_35_radr <= twiddle_rsc_0_35_i_radr;
  twiddle_rsc_0_35_i_q_d <= twiddle_rsc_0_35_i_q_d_1;
  twiddle_rsc_0_35_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_36_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_36_i_q,
      radr => twiddle_rsc_0_36_i_radr,
      q_d => twiddle_rsc_0_36_i_q_d_1,
      radr_d => twiddle_rsc_0_36_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_36_i_q <= twiddle_rsc_0_36_q;
  twiddle_rsc_0_36_radr <= twiddle_rsc_0_36_i_radr;
  twiddle_rsc_0_36_i_q_d <= twiddle_rsc_0_36_i_q_d_1;
  twiddle_rsc_0_36_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_37_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_37_i_q,
      radr => twiddle_rsc_0_37_i_radr,
      q_d => twiddle_rsc_0_37_i_q_d_1,
      radr_d => twiddle_rsc_0_37_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_37_i_q <= twiddle_rsc_0_37_q;
  twiddle_rsc_0_37_radr <= twiddle_rsc_0_37_i_radr;
  twiddle_rsc_0_37_i_q_d <= twiddle_rsc_0_37_i_q_d_1;
  twiddle_rsc_0_37_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_38_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_38_i_q,
      radr => twiddle_rsc_0_38_i_radr,
      q_d => twiddle_rsc_0_38_i_q_d_1,
      radr_d => twiddle_rsc_0_38_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_38_i_q <= twiddle_rsc_0_38_q;
  twiddle_rsc_0_38_radr <= twiddle_rsc_0_38_i_radr;
  twiddle_rsc_0_38_i_q_d <= twiddle_rsc_0_38_i_q_d_1;
  twiddle_rsc_0_38_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_39_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_39_i_q,
      radr => twiddle_rsc_0_39_i_radr,
      q_d => twiddle_rsc_0_39_i_q_d_1,
      radr_d => twiddle_rsc_0_39_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_39_i_q <= twiddle_rsc_0_39_q;
  twiddle_rsc_0_39_radr <= twiddle_rsc_0_39_i_radr;
  twiddle_rsc_0_39_i_q_d <= twiddle_rsc_0_39_i_q_d_1;
  twiddle_rsc_0_39_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_40_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_40_i_q,
      radr => twiddle_rsc_0_40_i_radr,
      q_d => twiddle_rsc_0_40_i_q_d_1,
      radr_d => twiddle_rsc_0_40_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_40_i_q <= twiddle_rsc_0_40_q;
  twiddle_rsc_0_40_radr <= twiddle_rsc_0_40_i_radr;
  twiddle_rsc_0_40_i_q_d <= twiddle_rsc_0_40_i_q_d_1;
  twiddle_rsc_0_40_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_41_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_41_i_q,
      radr => twiddle_rsc_0_41_i_radr,
      q_d => twiddle_rsc_0_41_i_q_d_1,
      radr_d => twiddle_rsc_0_41_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_41_i_q <= twiddle_rsc_0_41_q;
  twiddle_rsc_0_41_radr <= twiddle_rsc_0_41_i_radr;
  twiddle_rsc_0_41_i_q_d <= twiddle_rsc_0_41_i_q_d_1;
  twiddle_rsc_0_41_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_42_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_42_i_q,
      radr => twiddle_rsc_0_42_i_radr,
      q_d => twiddle_rsc_0_42_i_q_d_1,
      radr_d => twiddle_rsc_0_42_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_42_i_q <= twiddle_rsc_0_42_q;
  twiddle_rsc_0_42_radr <= twiddle_rsc_0_42_i_radr;
  twiddle_rsc_0_42_i_q_d <= twiddle_rsc_0_42_i_q_d_1;
  twiddle_rsc_0_42_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_43_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_43_i_q,
      radr => twiddle_rsc_0_43_i_radr,
      q_d => twiddle_rsc_0_43_i_q_d_1,
      radr_d => twiddle_rsc_0_43_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_43_i_q <= twiddle_rsc_0_43_q;
  twiddle_rsc_0_43_radr <= twiddle_rsc_0_43_i_radr;
  twiddle_rsc_0_43_i_q_d <= twiddle_rsc_0_43_i_q_d_1;
  twiddle_rsc_0_43_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_44_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_44_i_q,
      radr => twiddle_rsc_0_44_i_radr,
      q_d => twiddle_rsc_0_44_i_q_d_1,
      radr_d => twiddle_rsc_0_44_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_44_i_q <= twiddle_rsc_0_44_q;
  twiddle_rsc_0_44_radr <= twiddle_rsc_0_44_i_radr;
  twiddle_rsc_0_44_i_q_d <= twiddle_rsc_0_44_i_q_d_1;
  twiddle_rsc_0_44_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_45_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_45_i_q,
      radr => twiddle_rsc_0_45_i_radr,
      q_d => twiddle_rsc_0_45_i_q_d_1,
      radr_d => twiddle_rsc_0_45_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_45_i_q <= twiddle_rsc_0_45_q;
  twiddle_rsc_0_45_radr <= twiddle_rsc_0_45_i_radr;
  twiddle_rsc_0_45_i_q_d <= twiddle_rsc_0_45_i_q_d_1;
  twiddle_rsc_0_45_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_46_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_46_i_q,
      radr => twiddle_rsc_0_46_i_radr,
      q_d => twiddle_rsc_0_46_i_q_d_1,
      radr_d => twiddle_rsc_0_46_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_46_i_q <= twiddle_rsc_0_46_q;
  twiddle_rsc_0_46_radr <= twiddle_rsc_0_46_i_radr;
  twiddle_rsc_0_46_i_q_d <= twiddle_rsc_0_46_i_q_d_1;
  twiddle_rsc_0_46_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_47_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_47_i_q,
      radr => twiddle_rsc_0_47_i_radr,
      q_d => twiddle_rsc_0_47_i_q_d_1,
      radr_d => twiddle_rsc_0_47_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_47_i_q <= twiddle_rsc_0_47_q;
  twiddle_rsc_0_47_radr <= twiddle_rsc_0_47_i_radr;
  twiddle_rsc_0_47_i_q_d <= twiddle_rsc_0_47_i_q_d_1;
  twiddle_rsc_0_47_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_48_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_48_i_q,
      radr => twiddle_rsc_0_48_i_radr,
      q_d => twiddle_rsc_0_48_i_q_d_1,
      radr_d => twiddle_rsc_0_48_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_48_i_q <= twiddle_rsc_0_48_q;
  twiddle_rsc_0_48_radr <= twiddle_rsc_0_48_i_radr;
  twiddle_rsc_0_48_i_q_d <= twiddle_rsc_0_48_i_q_d_1;
  twiddle_rsc_0_48_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_49_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_49_i_q,
      radr => twiddle_rsc_0_49_i_radr,
      q_d => twiddle_rsc_0_49_i_q_d_1,
      radr_d => twiddle_rsc_0_49_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_49_i_q <= twiddle_rsc_0_49_q;
  twiddle_rsc_0_49_radr <= twiddle_rsc_0_49_i_radr;
  twiddle_rsc_0_49_i_q_d <= twiddle_rsc_0_49_i_q_d_1;
  twiddle_rsc_0_49_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_50_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_50_i_q,
      radr => twiddle_rsc_0_50_i_radr,
      q_d => twiddle_rsc_0_50_i_q_d_1,
      radr_d => twiddle_rsc_0_50_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_50_i_q <= twiddle_rsc_0_50_q;
  twiddle_rsc_0_50_radr <= twiddle_rsc_0_50_i_radr;
  twiddle_rsc_0_50_i_q_d <= twiddle_rsc_0_50_i_q_d_1;
  twiddle_rsc_0_50_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_51_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_51_i_q,
      radr => twiddle_rsc_0_51_i_radr,
      q_d => twiddle_rsc_0_51_i_q_d_1,
      radr_d => twiddle_rsc_0_51_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_51_i_q <= twiddle_rsc_0_51_q;
  twiddle_rsc_0_51_radr <= twiddle_rsc_0_51_i_radr;
  twiddle_rsc_0_51_i_q_d <= twiddle_rsc_0_51_i_q_d_1;
  twiddle_rsc_0_51_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_52_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_52_i_q,
      radr => twiddle_rsc_0_52_i_radr,
      q_d => twiddle_rsc_0_52_i_q_d_1,
      radr_d => twiddle_rsc_0_52_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_52_i_q <= twiddle_rsc_0_52_q;
  twiddle_rsc_0_52_radr <= twiddle_rsc_0_52_i_radr;
  twiddle_rsc_0_52_i_q_d <= twiddle_rsc_0_52_i_q_d_1;
  twiddle_rsc_0_52_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_53_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_53_i_q,
      radr => twiddle_rsc_0_53_i_radr,
      q_d => twiddle_rsc_0_53_i_q_d_1,
      radr_d => twiddle_rsc_0_53_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_53_i_q <= twiddle_rsc_0_53_q;
  twiddle_rsc_0_53_radr <= twiddle_rsc_0_53_i_radr;
  twiddle_rsc_0_53_i_q_d <= twiddle_rsc_0_53_i_q_d_1;
  twiddle_rsc_0_53_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_54_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_54_i_q,
      radr => twiddle_rsc_0_54_i_radr,
      q_d => twiddle_rsc_0_54_i_q_d_1,
      radr_d => twiddle_rsc_0_54_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_54_i_q <= twiddle_rsc_0_54_q;
  twiddle_rsc_0_54_radr <= twiddle_rsc_0_54_i_radr;
  twiddle_rsc_0_54_i_q_d <= twiddle_rsc_0_54_i_q_d_1;
  twiddle_rsc_0_54_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_55_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_55_i_q,
      radr => twiddle_rsc_0_55_i_radr,
      q_d => twiddle_rsc_0_55_i_q_d_1,
      radr_d => twiddle_rsc_0_55_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_55_i_q <= twiddle_rsc_0_55_q;
  twiddle_rsc_0_55_radr <= twiddle_rsc_0_55_i_radr;
  twiddle_rsc_0_55_i_q_d <= twiddle_rsc_0_55_i_q_d_1;
  twiddle_rsc_0_55_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_56_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_56_i_q,
      radr => twiddle_rsc_0_56_i_radr,
      q_d => twiddle_rsc_0_56_i_q_d_1,
      radr_d => twiddle_rsc_0_56_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_56_i_q <= twiddle_rsc_0_56_q;
  twiddle_rsc_0_56_radr <= twiddle_rsc_0_56_i_radr;
  twiddle_rsc_0_56_i_q_d <= twiddle_rsc_0_56_i_q_d_1;
  twiddle_rsc_0_56_i_radr_d <= twiddle_rsc_0_0_i_radr_d_iff;

  twiddle_rsc_0_57_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_57_i_q,
      radr => twiddle_rsc_0_57_i_radr,
      q_d => twiddle_rsc_0_57_i_q_d_1,
      radr_d => twiddle_rsc_0_57_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_57_i_q <= twiddle_rsc_0_57_q;
  twiddle_rsc_0_57_radr <= twiddle_rsc_0_57_i_radr;
  twiddle_rsc_0_57_i_q_d <= twiddle_rsc_0_57_i_q_d_1;
  twiddle_rsc_0_57_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_58_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_58_i_q,
      radr => twiddle_rsc_0_58_i_radr,
      q_d => twiddle_rsc_0_58_i_q_d_1,
      radr_d => twiddle_rsc_0_58_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_58_i_q <= twiddle_rsc_0_58_q;
  twiddle_rsc_0_58_radr <= twiddle_rsc_0_58_i_radr;
  twiddle_rsc_0_58_i_q_d <= twiddle_rsc_0_58_i_q_d_1;
  twiddle_rsc_0_58_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_59_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_59_i_q,
      radr => twiddle_rsc_0_59_i_radr,
      q_d => twiddle_rsc_0_59_i_q_d_1,
      radr_d => twiddle_rsc_0_59_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_59_i_q <= twiddle_rsc_0_59_q;
  twiddle_rsc_0_59_radr <= twiddle_rsc_0_59_i_radr;
  twiddle_rsc_0_59_i_q_d <= twiddle_rsc_0_59_i_q_d_1;
  twiddle_rsc_0_59_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_60_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_60_i_q,
      radr => twiddle_rsc_0_60_i_radr,
      q_d => twiddle_rsc_0_60_i_q_d_1,
      radr_d => twiddle_rsc_0_60_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_60_i_q <= twiddle_rsc_0_60_q;
  twiddle_rsc_0_60_radr <= twiddle_rsc_0_60_i_radr;
  twiddle_rsc_0_60_i_q_d <= twiddle_rsc_0_60_i_q_d_1;
  twiddle_rsc_0_60_i_radr_d <= twiddle_rsc_0_4_i_radr_d_iff;

  twiddle_rsc_0_61_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_61_i_q,
      radr => twiddle_rsc_0_61_i_radr,
      q_d => twiddle_rsc_0_61_i_q_d_1,
      radr_d => twiddle_rsc_0_61_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_61_i_q <= twiddle_rsc_0_61_q;
  twiddle_rsc_0_61_radr <= twiddle_rsc_0_61_i_radr;
  twiddle_rsc_0_61_i_q_d <= twiddle_rsc_0_61_i_q_d_1;
  twiddle_rsc_0_61_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  twiddle_rsc_0_62_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_62_i_q,
      radr => twiddle_rsc_0_62_i_radr,
      q_d => twiddle_rsc_0_62_i_q_d_1,
      radr_d => twiddle_rsc_0_62_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_62_i_q <= twiddle_rsc_0_62_q;
  twiddle_rsc_0_62_radr <= twiddle_rsc_0_62_i_radr;
  twiddle_rsc_0_62_i_q_d <= twiddle_rsc_0_62_i_q_d_1;
  twiddle_rsc_0_62_i_radr_d <= twiddle_rsc_0_2_i_radr_d_iff;

  twiddle_rsc_0_63_i : inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen
    PORT MAP(
      q => twiddle_rsc_0_63_i_q,
      radr => twiddle_rsc_0_63_i_radr,
      q_d => twiddle_rsc_0_63_i_q_d_1,
      radr_d => twiddle_rsc_0_63_i_radr_d,
      readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsc_0_63_i_q <= twiddle_rsc_0_63_q;
  twiddle_rsc_0_63_radr <= twiddle_rsc_0_63_i_radr;
  twiddle_rsc_0_63_i_q_d <= twiddle_rsc_0_63_i_q_d_1;
  twiddle_rsc_0_63_i_radr_d <= twiddle_rsc_0_1_i_radr_d_iff;

  inPlaceNTT_DIF_core_inst : inPlaceNTT_DIF_core
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      vec_rsc_triosy_0_8_lz => vec_rsc_triosy_0_8_lz,
      vec_rsc_triosy_0_9_lz => vec_rsc_triosy_0_9_lz,
      vec_rsc_triosy_0_10_lz => vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz => vec_rsc_triosy_0_11_lz,
      vec_rsc_triosy_0_12_lz => vec_rsc_triosy_0_12_lz,
      vec_rsc_triosy_0_13_lz => vec_rsc_triosy_0_13_lz,
      vec_rsc_triosy_0_14_lz => vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz => vec_rsc_triosy_0_15_lz,
      vec_rsc_triosy_0_16_lz => vec_rsc_triosy_0_16_lz,
      vec_rsc_triosy_0_17_lz => vec_rsc_triosy_0_17_lz,
      vec_rsc_triosy_0_18_lz => vec_rsc_triosy_0_18_lz,
      vec_rsc_triosy_0_19_lz => vec_rsc_triosy_0_19_lz,
      vec_rsc_triosy_0_20_lz => vec_rsc_triosy_0_20_lz,
      vec_rsc_triosy_0_21_lz => vec_rsc_triosy_0_21_lz,
      vec_rsc_triosy_0_22_lz => vec_rsc_triosy_0_22_lz,
      vec_rsc_triosy_0_23_lz => vec_rsc_triosy_0_23_lz,
      vec_rsc_triosy_0_24_lz => vec_rsc_triosy_0_24_lz,
      vec_rsc_triosy_0_25_lz => vec_rsc_triosy_0_25_lz,
      vec_rsc_triosy_0_26_lz => vec_rsc_triosy_0_26_lz,
      vec_rsc_triosy_0_27_lz => vec_rsc_triosy_0_27_lz,
      vec_rsc_triosy_0_28_lz => vec_rsc_triosy_0_28_lz,
      vec_rsc_triosy_0_29_lz => vec_rsc_triosy_0_29_lz,
      vec_rsc_triosy_0_30_lz => vec_rsc_triosy_0_30_lz,
      vec_rsc_triosy_0_31_lz => vec_rsc_triosy_0_31_lz,
      vec_rsc_triosy_0_32_lz => vec_rsc_triosy_0_32_lz,
      vec_rsc_triosy_0_33_lz => vec_rsc_triosy_0_33_lz,
      vec_rsc_triosy_0_34_lz => vec_rsc_triosy_0_34_lz,
      vec_rsc_triosy_0_35_lz => vec_rsc_triosy_0_35_lz,
      vec_rsc_triosy_0_36_lz => vec_rsc_triosy_0_36_lz,
      vec_rsc_triosy_0_37_lz => vec_rsc_triosy_0_37_lz,
      vec_rsc_triosy_0_38_lz => vec_rsc_triosy_0_38_lz,
      vec_rsc_triosy_0_39_lz => vec_rsc_triosy_0_39_lz,
      vec_rsc_triosy_0_40_lz => vec_rsc_triosy_0_40_lz,
      vec_rsc_triosy_0_41_lz => vec_rsc_triosy_0_41_lz,
      vec_rsc_triosy_0_42_lz => vec_rsc_triosy_0_42_lz,
      vec_rsc_triosy_0_43_lz => vec_rsc_triosy_0_43_lz,
      vec_rsc_triosy_0_44_lz => vec_rsc_triosy_0_44_lz,
      vec_rsc_triosy_0_45_lz => vec_rsc_triosy_0_45_lz,
      vec_rsc_triosy_0_46_lz => vec_rsc_triosy_0_46_lz,
      vec_rsc_triosy_0_47_lz => vec_rsc_triosy_0_47_lz,
      vec_rsc_triosy_0_48_lz => vec_rsc_triosy_0_48_lz,
      vec_rsc_triosy_0_49_lz => vec_rsc_triosy_0_49_lz,
      vec_rsc_triosy_0_50_lz => vec_rsc_triosy_0_50_lz,
      vec_rsc_triosy_0_51_lz => vec_rsc_triosy_0_51_lz,
      vec_rsc_triosy_0_52_lz => vec_rsc_triosy_0_52_lz,
      vec_rsc_triosy_0_53_lz => vec_rsc_triosy_0_53_lz,
      vec_rsc_triosy_0_54_lz => vec_rsc_triosy_0_54_lz,
      vec_rsc_triosy_0_55_lz => vec_rsc_triosy_0_55_lz,
      vec_rsc_triosy_0_56_lz => vec_rsc_triosy_0_56_lz,
      vec_rsc_triosy_0_57_lz => vec_rsc_triosy_0_57_lz,
      vec_rsc_triosy_0_58_lz => vec_rsc_triosy_0_58_lz,
      vec_rsc_triosy_0_59_lz => vec_rsc_triosy_0_59_lz,
      vec_rsc_triosy_0_60_lz => vec_rsc_triosy_0_60_lz,
      vec_rsc_triosy_0_61_lz => vec_rsc_triosy_0_61_lz,
      vec_rsc_triosy_0_62_lz => vec_rsc_triosy_0_62_lz,
      vec_rsc_triosy_0_63_lz => vec_rsc_triosy_0_63_lz,
      p_rsc_dat => inPlaceNTT_DIF_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_triosy_0_8_lz => twiddle_rsc_triosy_0_8_lz,
      twiddle_rsc_triosy_0_9_lz => twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_triosy_0_10_lz => twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_triosy_0_11_lz => twiddle_rsc_triosy_0_11_lz,
      twiddle_rsc_triosy_0_12_lz => twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_triosy_0_13_lz => twiddle_rsc_triosy_0_13_lz,
      twiddle_rsc_triosy_0_14_lz => twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_triosy_0_15_lz => twiddle_rsc_triosy_0_15_lz,
      twiddle_rsc_triosy_0_16_lz => twiddle_rsc_triosy_0_16_lz,
      twiddle_rsc_triosy_0_17_lz => twiddle_rsc_triosy_0_17_lz,
      twiddle_rsc_triosy_0_18_lz => twiddle_rsc_triosy_0_18_lz,
      twiddle_rsc_triosy_0_19_lz => twiddle_rsc_triosy_0_19_lz,
      twiddle_rsc_triosy_0_20_lz => twiddle_rsc_triosy_0_20_lz,
      twiddle_rsc_triosy_0_21_lz => twiddle_rsc_triosy_0_21_lz,
      twiddle_rsc_triosy_0_22_lz => twiddle_rsc_triosy_0_22_lz,
      twiddle_rsc_triosy_0_23_lz => twiddle_rsc_triosy_0_23_lz,
      twiddle_rsc_triosy_0_24_lz => twiddle_rsc_triosy_0_24_lz,
      twiddle_rsc_triosy_0_25_lz => twiddle_rsc_triosy_0_25_lz,
      twiddle_rsc_triosy_0_26_lz => twiddle_rsc_triosy_0_26_lz,
      twiddle_rsc_triosy_0_27_lz => twiddle_rsc_triosy_0_27_lz,
      twiddle_rsc_triosy_0_28_lz => twiddle_rsc_triosy_0_28_lz,
      twiddle_rsc_triosy_0_29_lz => twiddle_rsc_triosy_0_29_lz,
      twiddle_rsc_triosy_0_30_lz => twiddle_rsc_triosy_0_30_lz,
      twiddle_rsc_triosy_0_31_lz => twiddle_rsc_triosy_0_31_lz,
      twiddle_rsc_triosy_0_32_lz => twiddle_rsc_triosy_0_32_lz,
      twiddle_rsc_triosy_0_33_lz => twiddle_rsc_triosy_0_33_lz,
      twiddle_rsc_triosy_0_34_lz => twiddle_rsc_triosy_0_34_lz,
      twiddle_rsc_triosy_0_35_lz => twiddle_rsc_triosy_0_35_lz,
      twiddle_rsc_triosy_0_36_lz => twiddle_rsc_triosy_0_36_lz,
      twiddle_rsc_triosy_0_37_lz => twiddle_rsc_triosy_0_37_lz,
      twiddle_rsc_triosy_0_38_lz => twiddle_rsc_triosy_0_38_lz,
      twiddle_rsc_triosy_0_39_lz => twiddle_rsc_triosy_0_39_lz,
      twiddle_rsc_triosy_0_40_lz => twiddle_rsc_triosy_0_40_lz,
      twiddle_rsc_triosy_0_41_lz => twiddle_rsc_triosy_0_41_lz,
      twiddle_rsc_triosy_0_42_lz => twiddle_rsc_triosy_0_42_lz,
      twiddle_rsc_triosy_0_43_lz => twiddle_rsc_triosy_0_43_lz,
      twiddle_rsc_triosy_0_44_lz => twiddle_rsc_triosy_0_44_lz,
      twiddle_rsc_triosy_0_45_lz => twiddle_rsc_triosy_0_45_lz,
      twiddle_rsc_triosy_0_46_lz => twiddle_rsc_triosy_0_46_lz,
      twiddle_rsc_triosy_0_47_lz => twiddle_rsc_triosy_0_47_lz,
      twiddle_rsc_triosy_0_48_lz => twiddle_rsc_triosy_0_48_lz,
      twiddle_rsc_triosy_0_49_lz => twiddle_rsc_triosy_0_49_lz,
      twiddle_rsc_triosy_0_50_lz => twiddle_rsc_triosy_0_50_lz,
      twiddle_rsc_triosy_0_51_lz => twiddle_rsc_triosy_0_51_lz,
      twiddle_rsc_triosy_0_52_lz => twiddle_rsc_triosy_0_52_lz,
      twiddle_rsc_triosy_0_53_lz => twiddle_rsc_triosy_0_53_lz,
      twiddle_rsc_triosy_0_54_lz => twiddle_rsc_triosy_0_54_lz,
      twiddle_rsc_triosy_0_55_lz => twiddle_rsc_triosy_0_55_lz,
      twiddle_rsc_triosy_0_56_lz => twiddle_rsc_triosy_0_56_lz,
      twiddle_rsc_triosy_0_57_lz => twiddle_rsc_triosy_0_57_lz,
      twiddle_rsc_triosy_0_58_lz => twiddle_rsc_triosy_0_58_lz,
      twiddle_rsc_triosy_0_59_lz => twiddle_rsc_triosy_0_59_lz,
      twiddle_rsc_triosy_0_60_lz => twiddle_rsc_triosy_0_60_lz,
      twiddle_rsc_triosy_0_61_lz => twiddle_rsc_triosy_0_61_lz,
      twiddle_rsc_triosy_0_62_lz => twiddle_rsc_triosy_0_62_lz,
      twiddle_rsc_triosy_0_63_lz => twiddle_rsc_triosy_0_63_lz,
      vec_rsc_0_0_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d,
      vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d,
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d,
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d,
      vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d,
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d,
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d,
      vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d,
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_8_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d,
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d,
      vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_10_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d,
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_11_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d,
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d,
      vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_13_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d,
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_14_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d,
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d,
      vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_16_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_16_i_q_d,
      vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_17_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_17_i_q_d,
      vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_18_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_18_i_q_d,
      vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_19_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_19_i_q_d,
      vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_20_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_20_i_q_d,
      vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_21_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_21_i_q_d,
      vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_22_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_22_i_q_d,
      vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_23_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_23_i_q_d,
      vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_24_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_24_i_q_d,
      vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_25_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_25_i_q_d,
      vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_26_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_26_i_q_d,
      vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_27_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_27_i_q_d,
      vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_28_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_28_i_q_d,
      vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_29_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_29_i_q_d,
      vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_30_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_30_i_q_d,
      vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_31_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_31_i_q_d,
      vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_32_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_32_i_q_d,
      vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_33_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_33_i_q_d,
      vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_34_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_34_i_q_d,
      vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_35_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_35_i_q_d,
      vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_36_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_36_i_q_d,
      vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_37_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_37_i_q_d,
      vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_38_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_38_i_q_d,
      vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_39_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_39_i_q_d,
      vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_40_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_40_i_q_d,
      vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_41_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_41_i_q_d,
      vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_42_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_42_i_q_d,
      vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_43_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_43_i_q_d,
      vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_44_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_44_i_q_d,
      vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_45_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_45_i_q_d,
      vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_46_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_46_i_q_d,
      vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_47_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_47_i_q_d,
      vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_48_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_48_i_q_d,
      vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_49_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_49_i_q_d,
      vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_50_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_50_i_q_d,
      vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_51_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_51_i_q_d,
      vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_52_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_52_i_q_d,
      vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_53_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_53_i_q_d,
      vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_54_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_54_i_q_d,
      vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_55_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_55_i_q_d,
      vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_56_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_56_i_q_d,
      vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_57_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_57_i_q_d,
      vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_58_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_58_i_q_d,
      vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_59_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_59_i_q_d,
      vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_60_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_60_i_q_d,
      vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_61_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_61_i_q_d,
      vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_62_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_62_i_q_d,
      vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_63_i_q_d => inPlaceNTT_DIF_core_inst_vec_rsc_0_63_i_q_d,
      vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_0_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d,
      twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d,
      twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d,
      twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d,
      twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d,
      twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d,
      twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d,
      twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d,
      twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_8_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d,
      twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_9_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d,
      twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_10_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d,
      twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_11_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d,
      twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_12_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d,
      twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_13_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d,
      twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_14_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d,
      twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_15_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d,
      twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_16_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_16_i_q_d,
      twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_17_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_17_i_q_d,
      twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_18_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_18_i_q_d,
      twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_19_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_19_i_q_d,
      twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_20_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_20_i_q_d,
      twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_21_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_21_i_q_d,
      twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_22_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_22_i_q_d,
      twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_23_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_23_i_q_d,
      twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_24_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_24_i_q_d,
      twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_25_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_25_i_q_d,
      twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_26_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_26_i_q_d,
      twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_27_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_27_i_q_d,
      twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_28_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_28_i_q_d,
      twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_29_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_29_i_q_d,
      twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_30_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_30_i_q_d,
      twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_31_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_31_i_q_d,
      twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_32_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_32_i_q_d,
      twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_33_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_33_i_q_d,
      twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_34_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_34_i_q_d,
      twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_35_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_35_i_q_d,
      twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_36_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_36_i_q_d,
      twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_37_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_37_i_q_d,
      twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_38_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_38_i_q_d,
      twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_39_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_39_i_q_d,
      twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_40_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_40_i_q_d,
      twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_41_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_41_i_q_d,
      twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_42_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_42_i_q_d,
      twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_43_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_43_i_q_d,
      twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_44_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_44_i_q_d,
      twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_45_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_45_i_q_d,
      twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_46_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_46_i_q_d,
      twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_47_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_47_i_q_d,
      twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_48_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_48_i_q_d,
      twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_49_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_49_i_q_d,
      twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_50_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_50_i_q_d,
      twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_51_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_51_i_q_d,
      twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_52_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_52_i_q_d,
      twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_53_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_53_i_q_d,
      twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_54_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_54_i_q_d,
      twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_55_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_55_i_q_d,
      twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_56_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_56_i_q_d,
      twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_57_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_57_i_q_d,
      twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_58_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_58_i_q_d,
      twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_59_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_59_i_q_d,
      twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_60_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_60_i_q_d,
      twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_61_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_61_i_q_d,
      twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_62_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_62_i_q_d,
      twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_63_i_q_d => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_63_i_q_d,
      twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d => twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_d_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff,
      vec_rsc_0_0_i_radr_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff,
      vec_rsc_0_0_i_wadr_d_pff => inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff,
      vec_rsc_0_0_i_we_d_pff => vec_rsc_0_0_i_we_d_iff,
      vec_rsc_0_1_i_we_d_pff => vec_rsc_0_1_i_we_d_iff,
      vec_rsc_0_2_i_we_d_pff => vec_rsc_0_2_i_we_d_iff,
      vec_rsc_0_3_i_we_d_pff => vec_rsc_0_3_i_we_d_iff,
      vec_rsc_0_4_i_we_d_pff => vec_rsc_0_4_i_we_d_iff,
      vec_rsc_0_5_i_we_d_pff => vec_rsc_0_5_i_we_d_iff,
      vec_rsc_0_6_i_we_d_pff => vec_rsc_0_6_i_we_d_iff,
      vec_rsc_0_7_i_we_d_pff => vec_rsc_0_7_i_we_d_iff,
      vec_rsc_0_8_i_we_d_pff => vec_rsc_0_8_i_we_d_iff,
      vec_rsc_0_9_i_we_d_pff => vec_rsc_0_9_i_we_d_iff,
      vec_rsc_0_10_i_we_d_pff => vec_rsc_0_10_i_we_d_iff,
      vec_rsc_0_11_i_we_d_pff => vec_rsc_0_11_i_we_d_iff,
      vec_rsc_0_12_i_we_d_pff => vec_rsc_0_12_i_we_d_iff,
      vec_rsc_0_13_i_we_d_pff => vec_rsc_0_13_i_we_d_iff,
      vec_rsc_0_14_i_we_d_pff => vec_rsc_0_14_i_we_d_iff,
      vec_rsc_0_15_i_we_d_pff => vec_rsc_0_15_i_we_d_iff,
      vec_rsc_0_16_i_we_d_pff => vec_rsc_0_16_i_we_d_iff,
      vec_rsc_0_17_i_we_d_pff => vec_rsc_0_17_i_we_d_iff,
      vec_rsc_0_18_i_we_d_pff => vec_rsc_0_18_i_we_d_iff,
      vec_rsc_0_19_i_we_d_pff => vec_rsc_0_19_i_we_d_iff,
      vec_rsc_0_20_i_we_d_pff => vec_rsc_0_20_i_we_d_iff,
      vec_rsc_0_21_i_we_d_pff => vec_rsc_0_21_i_we_d_iff,
      vec_rsc_0_22_i_we_d_pff => vec_rsc_0_22_i_we_d_iff,
      vec_rsc_0_23_i_we_d_pff => vec_rsc_0_23_i_we_d_iff,
      vec_rsc_0_24_i_we_d_pff => vec_rsc_0_24_i_we_d_iff,
      vec_rsc_0_25_i_we_d_pff => vec_rsc_0_25_i_we_d_iff,
      vec_rsc_0_26_i_we_d_pff => vec_rsc_0_26_i_we_d_iff,
      vec_rsc_0_27_i_we_d_pff => vec_rsc_0_27_i_we_d_iff,
      vec_rsc_0_28_i_we_d_pff => vec_rsc_0_28_i_we_d_iff,
      vec_rsc_0_29_i_we_d_pff => vec_rsc_0_29_i_we_d_iff,
      vec_rsc_0_30_i_we_d_pff => vec_rsc_0_30_i_we_d_iff,
      vec_rsc_0_31_i_we_d_pff => vec_rsc_0_31_i_we_d_iff,
      vec_rsc_0_32_i_we_d_pff => vec_rsc_0_32_i_we_d_iff,
      vec_rsc_0_33_i_we_d_pff => vec_rsc_0_33_i_we_d_iff,
      vec_rsc_0_34_i_we_d_pff => vec_rsc_0_34_i_we_d_iff,
      vec_rsc_0_35_i_we_d_pff => vec_rsc_0_35_i_we_d_iff,
      vec_rsc_0_36_i_we_d_pff => vec_rsc_0_36_i_we_d_iff,
      vec_rsc_0_37_i_we_d_pff => vec_rsc_0_37_i_we_d_iff,
      vec_rsc_0_38_i_we_d_pff => vec_rsc_0_38_i_we_d_iff,
      vec_rsc_0_39_i_we_d_pff => vec_rsc_0_39_i_we_d_iff,
      vec_rsc_0_40_i_we_d_pff => vec_rsc_0_40_i_we_d_iff,
      vec_rsc_0_41_i_we_d_pff => vec_rsc_0_41_i_we_d_iff,
      vec_rsc_0_42_i_we_d_pff => vec_rsc_0_42_i_we_d_iff,
      vec_rsc_0_43_i_we_d_pff => vec_rsc_0_43_i_we_d_iff,
      vec_rsc_0_44_i_we_d_pff => vec_rsc_0_44_i_we_d_iff,
      vec_rsc_0_45_i_we_d_pff => vec_rsc_0_45_i_we_d_iff,
      vec_rsc_0_46_i_we_d_pff => vec_rsc_0_46_i_we_d_iff,
      vec_rsc_0_47_i_we_d_pff => vec_rsc_0_47_i_we_d_iff,
      vec_rsc_0_48_i_we_d_pff => vec_rsc_0_48_i_we_d_iff,
      vec_rsc_0_49_i_we_d_pff => vec_rsc_0_49_i_we_d_iff,
      vec_rsc_0_50_i_we_d_pff => vec_rsc_0_50_i_we_d_iff,
      vec_rsc_0_51_i_we_d_pff => vec_rsc_0_51_i_we_d_iff,
      vec_rsc_0_52_i_we_d_pff => vec_rsc_0_52_i_we_d_iff,
      vec_rsc_0_53_i_we_d_pff => vec_rsc_0_53_i_we_d_iff,
      vec_rsc_0_54_i_we_d_pff => vec_rsc_0_54_i_we_d_iff,
      vec_rsc_0_55_i_we_d_pff => vec_rsc_0_55_i_we_d_iff,
      vec_rsc_0_56_i_we_d_pff => vec_rsc_0_56_i_we_d_iff,
      vec_rsc_0_57_i_we_d_pff => vec_rsc_0_57_i_we_d_iff,
      vec_rsc_0_58_i_we_d_pff => vec_rsc_0_58_i_we_d_iff,
      vec_rsc_0_59_i_we_d_pff => vec_rsc_0_59_i_we_d_iff,
      vec_rsc_0_60_i_we_d_pff => vec_rsc_0_60_i_we_d_iff,
      vec_rsc_0_61_i_we_d_pff => vec_rsc_0_61_i_we_d_iff,
      vec_rsc_0_62_i_we_d_pff => vec_rsc_0_62_i_we_d_iff,
      vec_rsc_0_63_i_we_d_pff => vec_rsc_0_63_i_we_d_iff,
      twiddle_rsc_0_0_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d_pff,
      twiddle_rsc_0_1_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff,
      twiddle_rsc_0_2_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff,
      twiddle_rsc_0_4_i_radr_d_pff => inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff
    );
  inPlaceNTT_DIF_core_inst_p_rsc_dat <= p_rsc_dat;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_q_d <= vec_rsc_0_0_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_1_i_q_d <= vec_rsc_0_1_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_2_i_q_d <= vec_rsc_0_2_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_3_i_q_d <= vec_rsc_0_3_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_4_i_q_d <= vec_rsc_0_4_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_5_i_q_d <= vec_rsc_0_5_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_6_i_q_d <= vec_rsc_0_6_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_7_i_q_d <= vec_rsc_0_7_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_8_i_q_d <= vec_rsc_0_8_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_9_i_q_d <= vec_rsc_0_9_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_10_i_q_d <= vec_rsc_0_10_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_11_i_q_d <= vec_rsc_0_11_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_12_i_q_d <= vec_rsc_0_12_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_13_i_q_d <= vec_rsc_0_13_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_14_i_q_d <= vec_rsc_0_14_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_15_i_q_d <= vec_rsc_0_15_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_16_i_q_d <= vec_rsc_0_16_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_17_i_q_d <= vec_rsc_0_17_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_18_i_q_d <= vec_rsc_0_18_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_19_i_q_d <= vec_rsc_0_19_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_20_i_q_d <= vec_rsc_0_20_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_21_i_q_d <= vec_rsc_0_21_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_22_i_q_d <= vec_rsc_0_22_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_23_i_q_d <= vec_rsc_0_23_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_24_i_q_d <= vec_rsc_0_24_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_25_i_q_d <= vec_rsc_0_25_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_26_i_q_d <= vec_rsc_0_26_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_27_i_q_d <= vec_rsc_0_27_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_28_i_q_d <= vec_rsc_0_28_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_29_i_q_d <= vec_rsc_0_29_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_30_i_q_d <= vec_rsc_0_30_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_31_i_q_d <= vec_rsc_0_31_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_32_i_q_d <= vec_rsc_0_32_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_33_i_q_d <= vec_rsc_0_33_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_34_i_q_d <= vec_rsc_0_34_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_35_i_q_d <= vec_rsc_0_35_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_36_i_q_d <= vec_rsc_0_36_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_37_i_q_d <= vec_rsc_0_37_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_38_i_q_d <= vec_rsc_0_38_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_39_i_q_d <= vec_rsc_0_39_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_40_i_q_d <= vec_rsc_0_40_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_41_i_q_d <= vec_rsc_0_41_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_42_i_q_d <= vec_rsc_0_42_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_43_i_q_d <= vec_rsc_0_43_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_44_i_q_d <= vec_rsc_0_44_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_45_i_q_d <= vec_rsc_0_45_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_46_i_q_d <= vec_rsc_0_46_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_47_i_q_d <= vec_rsc_0_47_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_48_i_q_d <= vec_rsc_0_48_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_49_i_q_d <= vec_rsc_0_49_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_50_i_q_d <= vec_rsc_0_50_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_51_i_q_d <= vec_rsc_0_51_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_52_i_q_d <= vec_rsc_0_52_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_53_i_q_d <= vec_rsc_0_53_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_54_i_q_d <= vec_rsc_0_54_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_55_i_q_d <= vec_rsc_0_55_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_56_i_q_d <= vec_rsc_0_56_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_57_i_q_d <= vec_rsc_0_57_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_58_i_q_d <= vec_rsc_0_58_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_59_i_q_d <= vec_rsc_0_59_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_60_i_q_d <= vec_rsc_0_60_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_61_i_q_d <= vec_rsc_0_61_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_62_i_q_d <= vec_rsc_0_62_i_q_d;
  inPlaceNTT_DIF_core_inst_vec_rsc_0_63_i_q_d <= vec_rsc_0_63_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_q_d <= twiddle_rsc_0_0_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_q_d <= twiddle_rsc_0_1_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_q_d <= twiddle_rsc_0_2_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_3_i_q_d <= twiddle_rsc_0_3_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_q_d <= twiddle_rsc_0_4_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_5_i_q_d <= twiddle_rsc_0_5_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_6_i_q_d <= twiddle_rsc_0_6_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_7_i_q_d <= twiddle_rsc_0_7_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_8_i_q_d <= twiddle_rsc_0_8_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_9_i_q_d <= twiddle_rsc_0_9_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_10_i_q_d <= twiddle_rsc_0_10_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_11_i_q_d <= twiddle_rsc_0_11_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_12_i_q_d <= twiddle_rsc_0_12_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_13_i_q_d <= twiddle_rsc_0_13_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_14_i_q_d <= twiddle_rsc_0_14_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_15_i_q_d <= twiddle_rsc_0_15_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_16_i_q_d <= twiddle_rsc_0_16_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_17_i_q_d <= twiddle_rsc_0_17_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_18_i_q_d <= twiddle_rsc_0_18_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_19_i_q_d <= twiddle_rsc_0_19_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_20_i_q_d <= twiddle_rsc_0_20_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_21_i_q_d <= twiddle_rsc_0_21_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_22_i_q_d <= twiddle_rsc_0_22_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_23_i_q_d <= twiddle_rsc_0_23_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_24_i_q_d <= twiddle_rsc_0_24_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_25_i_q_d <= twiddle_rsc_0_25_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_26_i_q_d <= twiddle_rsc_0_26_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_27_i_q_d <= twiddle_rsc_0_27_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_28_i_q_d <= twiddle_rsc_0_28_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_29_i_q_d <= twiddle_rsc_0_29_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_30_i_q_d <= twiddle_rsc_0_30_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_31_i_q_d <= twiddle_rsc_0_31_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_32_i_q_d <= twiddle_rsc_0_32_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_33_i_q_d <= twiddle_rsc_0_33_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_34_i_q_d <= twiddle_rsc_0_34_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_35_i_q_d <= twiddle_rsc_0_35_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_36_i_q_d <= twiddle_rsc_0_36_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_37_i_q_d <= twiddle_rsc_0_37_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_38_i_q_d <= twiddle_rsc_0_38_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_39_i_q_d <= twiddle_rsc_0_39_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_40_i_q_d <= twiddle_rsc_0_40_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_41_i_q_d <= twiddle_rsc_0_41_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_42_i_q_d <= twiddle_rsc_0_42_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_43_i_q_d <= twiddle_rsc_0_43_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_44_i_q_d <= twiddle_rsc_0_44_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_45_i_q_d <= twiddle_rsc_0_45_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_46_i_q_d <= twiddle_rsc_0_46_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_47_i_q_d <= twiddle_rsc_0_47_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_48_i_q_d <= twiddle_rsc_0_48_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_49_i_q_d <= twiddle_rsc_0_49_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_50_i_q_d <= twiddle_rsc_0_50_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_51_i_q_d <= twiddle_rsc_0_51_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_52_i_q_d <= twiddle_rsc_0_52_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_53_i_q_d <= twiddle_rsc_0_53_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_54_i_q_d <= twiddle_rsc_0_54_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_55_i_q_d <= twiddle_rsc_0_55_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_56_i_q_d <= twiddle_rsc_0_56_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_57_i_q_d <= twiddle_rsc_0_57_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_58_i_q_d <= twiddle_rsc_0_58_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_59_i_q_d <= twiddle_rsc_0_59_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_60_i_q_d <= twiddle_rsc_0_60_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_61_i_q_d <= twiddle_rsc_0_61_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_62_i_q_d <= twiddle_rsc_0_62_i_q_d;
  inPlaceNTT_DIF_core_inst_twiddle_rsc_0_63_i_q_d <= twiddle_rsc_0_63_i_q_d;
  vec_rsc_0_0_i_d_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_d_d_pff;
  vec_rsc_0_0_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_radr_d_pff;
  vec_rsc_0_0_i_wadr_d_iff <= inPlaceNTT_DIF_core_inst_vec_rsc_0_0_i_wadr_d_pff;
  twiddle_rsc_0_0_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_0_i_radr_d_pff;
  twiddle_rsc_0_1_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_1_i_radr_d_pff;
  twiddle_rsc_0_2_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_2_i_radr_d_pff;
  twiddle_rsc_0_4_i_radr_d_iff <= inPlaceNTT_DIF_core_inst_twiddle_rsc_0_4_i_radr_d_pff;

END v14;



