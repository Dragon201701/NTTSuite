
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   jd4691@newnano.poly.edu
//  Generated date: Tue Jun 22 23:59:02 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_filter_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_filter_core_core_fsm (
  clk, rst, fsm_output, SHIFT_LOOP_C_0_tr0, MAC_LOOP_C_0_tr0
);
  input clk;
  input rst;
  output [4:0] fsm_output;
  reg [4:0] fsm_output;
  input SHIFT_LOOP_C_0_tr0;
  input MAC_LOOP_C_0_tr0;


  // FSM State Type Declaration for fir_filter_core_core_fsm_1
  parameter
    main_C_0 = 3'd0,
    SHIFT_LOOP_C_0 = 3'd1,
    MAC_LOOP_C_0 = 3'd2,
    main_C_1 = 3'd3,
    main_C_2 = 3'd4;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_filter_core_core_fsm_1
    case (state_var)
      SHIFT_LOOP_C_0 : begin
        fsm_output = 5'b00010;
        if ( SHIFT_LOOP_C_0_tr0 ) begin
          state_var_NS = MAC_LOOP_C_0;
        end
        else begin
          state_var_NS = SHIFT_LOOP_C_0;
        end
      end
      MAC_LOOP_C_0 : begin
        fsm_output = 5'b00100;
        if ( MAC_LOOP_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = MAC_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 5'b01000;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 5'b10000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 5'b00001;
        state_var_NS = SHIFT_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_filter_core
// ------------------------------------------------------------------


module fir_filter_core (
  clk, rst, i_sample_rsc_dat, i_sample_rsc_triosy_lz, b_rsc_dat, b_rsc_triosy_lz,
      y_rsc_dat, y_rsc_triosy_lz
);
  input clk;
  input rst;
  input [2:0] i_sample_rsc_dat;
  output i_sample_rsc_triosy_lz;
  input [1269:0] b_rsc_dat;
  output b_rsc_triosy_lz;
  output [8:0] y_rsc_dat;
  output y_rsc_triosy_lz;


  // Interconnect Declarations
  wire [2:0] i_sample_rsci_idat;
  wire [1269:0] b_rsci_idat;
  reg y_rsc_triosy_obj_ld;
  reg y_rsci_idat_8;
  reg [6:0] y_rsci_idat_7_1;
  reg y_rsci_idat_0;
  wire [4:0] fsm_output;
  wire or_dcpl_9;
  wire or_dcpl_10;
  wire or_dcpl_11;
  wire or_dcpl_12;
  wire or_dcpl_13;
  wire or_dcpl_15;
  wire or_dcpl_16;
  wire or_dcpl_17;
  wire or_dcpl_19;
  wire or_dcpl_20;
  wire or_dcpl_21;
  wire or_dcpl_22;
  wire or_dcpl_23;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire or_dcpl_28;
  wire or_dcpl_30;
  wire or_dcpl_34;
  wire or_dcpl_36;
  wire or_dcpl_40;
  wire or_dcpl_42;
  wire or_dcpl_43;
  wire or_dcpl_47;
  wire or_dcpl_48;
  wire or_dcpl_50;
  wire or_dcpl_54;
  wire or_dcpl_56;
  wire or_dcpl_60;
  wire or_dcpl_62;
  wire or_dcpl_66;
  wire or_dcpl_100;
  wire or_dcpl_101;
  wire or_dcpl_104;
  wire or_dcpl_106;
  wire or_dcpl_107;
  wire or_dcpl_110;
  reg [19:0] sum_sva;
  reg [6:0] MAC_LOOP_n_6_0_sva;
  reg reg_b_rsc_triosy_obj_ld_cse;
  wire [2:0] z_out;
  wire [6:0] z_out_2;
  wire [7:0] nl_z_out_2;
  wire [19:0] z_out_3;
  wire [20:0] nl_z_out_3;
  reg [2:0] x_0_sva;
  reg [2:0] x_63_lpi_2;
  reg [2:0] x_62_lpi_2;
  reg [2:0] x_64_lpi_2;
  reg [2:0] x_61_lpi_2;
  reg [2:0] x_65_lpi_2;
  reg [2:0] x_60_lpi_2;
  reg [2:0] x_66_lpi_2;
  reg [2:0] x_59_lpi_2;
  reg [2:0] x_67_lpi_2;
  reg [2:0] x_58_lpi_2;
  reg [2:0] x_68_lpi_2;
  reg [2:0] x_57_lpi_2;
  reg [2:0] x_69_lpi_2;
  reg [2:0] x_56_lpi_2;
  reg [2:0] x_70_lpi_2;
  reg [2:0] x_55_lpi_2;
  reg [2:0] x_71_lpi_2;
  reg [2:0] x_54_lpi_2;
  reg [2:0] x_72_lpi_2;
  reg [2:0] x_53_lpi_2;
  reg [2:0] x_73_lpi_2;
  reg [2:0] x_52_lpi_2;
  reg [2:0] x_74_lpi_2;
  reg [2:0] x_51_lpi_2;
  reg [2:0] x_75_lpi_2;
  reg [2:0] x_50_lpi_2;
  reg [2:0] x_76_lpi_2;
  reg [2:0] x_49_lpi_2;
  reg [2:0] x_77_lpi_2;
  reg [2:0] x_48_lpi_2;
  reg [2:0] x_78_lpi_2;
  reg [2:0] x_47_lpi_2;
  reg [2:0] x_79_lpi_2;
  reg [2:0] x_46_lpi_2;
  reg [2:0] x_80_lpi_2;
  reg [2:0] x_45_lpi_2;
  reg [2:0] x_81_lpi_2;
  reg [2:0] x_44_lpi_2;
  reg [2:0] x_82_lpi_2;
  reg [2:0] x_43_lpi_2;
  reg [2:0] x_83_lpi_2;
  reg [2:0] x_42_lpi_2;
  reg [2:0] x_84_lpi_2;
  reg [2:0] x_41_lpi_2;
  reg [2:0] x_85_lpi_2;
  reg [2:0] x_40_lpi_2;
  reg [2:0] x_86_lpi_2;
  reg [2:0] x_39_lpi_2;
  reg [2:0] x_87_lpi_2;
  reg [2:0] x_38_lpi_2;
  reg [2:0] x_88_lpi_2;
  reg [2:0] x_37_lpi_2;
  reg [2:0] x_89_lpi_2;
  reg [2:0] x_36_lpi_2;
  reg [2:0] x_90_lpi_2;
  reg [2:0] x_35_lpi_2;
  reg [2:0] x_91_lpi_2;
  reg [2:0] x_34_lpi_2;
  reg [2:0] x_92_lpi_2;
  reg [2:0] x_33_lpi_2;
  reg [2:0] x_93_lpi_2;
  reg [2:0] x_32_lpi_2;
  reg [2:0] x_94_lpi_2;
  reg [2:0] x_31_lpi_2;
  reg [2:0] x_95_lpi_2;
  reg [2:0] x_30_lpi_2;
  reg [2:0] x_96_lpi_2;
  reg [2:0] x_29_lpi_2;
  reg [2:0] x_97_lpi_2;
  reg [2:0] x_28_lpi_2;
  reg [2:0] x_98_lpi_2;
  reg [2:0] x_27_lpi_2;
  reg [2:0] x_99_lpi_2;
  reg [2:0] x_26_lpi_2;
  reg [2:0] x_100_lpi_2;
  reg [2:0] x_25_lpi_2;
  reg [2:0] x_101_lpi_2;
  reg [2:0] x_24_lpi_2;
  reg [2:0] x_102_lpi_2;
  reg [2:0] x_23_lpi_2;
  reg [2:0] x_103_lpi_2;
  reg [2:0] x_22_lpi_2;
  reg [2:0] x_104_lpi_2;
  reg [2:0] x_21_lpi_2;
  reg [2:0] x_105_lpi_2;
  reg [2:0] x_20_lpi_2;
  reg [2:0] x_106_lpi_2;
  reg [2:0] x_19_lpi_2;
  reg [2:0] x_107_lpi_2;
  reg [2:0] x_18_lpi_2;
  reg [2:0] x_108_lpi_2;
  reg [2:0] x_17_lpi_2;
  reg [2:0] x_109_lpi_2;
  reg [2:0] x_16_lpi_2;
  reg [2:0] x_110_lpi_2;
  reg [2:0] x_15_lpi_2;
  reg [2:0] x_111_lpi_2;
  reg [2:0] x_14_lpi_2;
  reg [2:0] x_112_lpi_2;
  reg [2:0] x_13_lpi_2;
  reg [2:0] x_113_lpi_2;
  reg [2:0] x_12_lpi_2;
  reg [2:0] x_114_lpi_2;
  reg [2:0] x_11_lpi_2;
  reg [2:0] x_115_lpi_2;
  reg [2:0] x_10_lpi_2;
  reg [2:0] x_116_lpi_2;
  reg [2:0] x_9_lpi_2;
  reg [2:0] x_117_lpi_2;
  reg [2:0] x_8_lpi_2;
  reg [2:0] x_118_lpi_2;
  reg [2:0] x_7_lpi_2;
  reg [2:0] x_119_lpi_2;
  reg [2:0] x_6_lpi_2;
  reg [2:0] x_120_lpi_2;
  reg [2:0] x_5_lpi_2;
  reg [2:0] x_121_lpi_2;
  reg [2:0] x_4_lpi_2;
  reg [2:0] x_122_lpi_2;
  reg [2:0] x_3_lpi_2;
  reg [2:0] x_123_lpi_2;
  reg [2:0] x_2_lpi_2;
  reg [2:0] x_124_lpi_2;
  reg [2:0] x_1_lpi_2;
  reg [2:0] x_125_lpi_2;
  reg [2:0] x_126_lpi_2;
  reg [2:0] i_sample_sva;
  wire nor_ovfl_sva_1;
  wire and_unfl_sva_1;
  wire z_out_1_7;

  wire[6:0] nor_5_nl;
  wire[6:0] SHIFT_LOOP_n_SHIFT_LOOP_n_mux_nl;
  wire[0:0] SHIFT_LOOP_n_or_nl;
  wire[0:0] MAC_LOOP_n_nor_nl;
  wire[7:0] SHIFT_LOOP_acc_nl;
  wire[8:0] nl_SHIFT_LOOP_acc_nl;
  wire[6:0] SHIFT_LOOP_mux_129_nl;
  wire[18:0] MAC_LOOP_mux_7_nl;
  wire[12:0] MAC_LOOP_mux_8_nl;
  wire[12:0] MAC_LOOP_mul_1_nl;
  wire[9:0] MAC_LOOP_mux_9_nl;
  wire[2:0] MAC_LOOP_mux_10_nl;
  wire[6:0] MAC_LOOP_mux_11_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [8:0] nl_y_rsci_idat;
  assign nl_y_rsci_idat = {y_rsci_idat_8 , y_rsci_idat_7_1 , y_rsci_idat_0};
  wire [0:0] nl_fir_filter_core_core_fsm_inst_SHIFT_LOOP_C_0_tr0;
  assign nl_fir_filter_core_core_fsm_inst_SHIFT_LOOP_C_0_tr0 = ~ z_out_1_7;
  wire [0:0] nl_fir_filter_core_core_fsm_inst_MAC_LOOP_C_0_tr0;
  assign nl_fir_filter_core_core_fsm_inst_MAC_LOOP_C_0_tr0 = ~ z_out_1_7;
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd3)) i_sample_rsci (
      .dat(i_sample_rsc_dat),
      .idat(i_sample_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd1270)) b_rsci (
      .dat(b_rsc_dat),
      .idat(b_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd9)) y_rsci (
      .idat(nl_y_rsci_idat[8:0]),
      .dat(y_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) i_sample_rsc_triosy_obj (
      .ld(reg_b_rsc_triosy_obj_ld_cse),
      .lz(i_sample_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) b_rsc_triosy_obj (
      .ld(reg_b_rsc_triosy_obj_ld_cse),
      .lz(b_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) y_rsc_triosy_obj (
      .ld(y_rsc_triosy_obj_ld),
      .lz(y_rsc_triosy_lz)
    );
  fir_filter_core_core_fsm fir_filter_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .SHIFT_LOOP_C_0_tr0(nl_fir_filter_core_core_fsm_inst_SHIFT_LOOP_C_0_tr0[0:0]),
      .MAC_LOOP_C_0_tr0(nl_fir_filter_core_core_fsm_inst_MAC_LOOP_C_0_tr0[0:0])
    );
  assign nor_ovfl_sva_1 = ~((z_out_3[14]) | (~((z_out_3[13:8]!=6'b000000))));
  assign and_unfl_sva_1 = (z_out_3[14]) & (~((z_out_3[13:8]==6'b111111) & ((z_out_3[7:0]!=8'b00000000))));
  assign or_dcpl_9 = ~((MAC_LOOP_n_6_0_sva[6:5]==2'b11));
  assign or_dcpl_10 = or_dcpl_9 | (MAC_LOOP_n_6_0_sva[0]);
  assign or_dcpl_11 = ~((MAC_LOOP_n_6_0_sva[4:3]==2'b11));
  assign or_dcpl_12 = ~((MAC_LOOP_n_6_0_sva[2:1]==2'b11));
  assign or_dcpl_13 = or_dcpl_12 | or_dcpl_11;
  assign or_dcpl_15 = or_dcpl_9 | (~ (MAC_LOOP_n_6_0_sva[0]));
  assign or_dcpl_16 = (MAC_LOOP_n_6_0_sva[2:1]!=2'b10);
  assign or_dcpl_17 = or_dcpl_16 | or_dcpl_11;
  assign or_dcpl_19 = (MAC_LOOP_n_6_0_sva[6:5]!=2'b00);
  assign or_dcpl_20 = or_dcpl_19 | (~ (MAC_LOOP_n_6_0_sva[0]));
  assign or_dcpl_21 = (MAC_LOOP_n_6_0_sva[4:3]!=2'b00);
  assign or_dcpl_22 = (MAC_LOOP_n_6_0_sva[2:1]!=2'b00);
  assign or_dcpl_23 = or_dcpl_22 | or_dcpl_21;
  assign or_dcpl_26 = or_dcpl_19 | (MAC_LOOP_n_6_0_sva[0]);
  assign or_dcpl_27 = (MAC_LOOP_n_6_0_sva[2:1]!=2'b01);
  assign or_dcpl_28 = or_dcpl_27 | or_dcpl_21;
  assign or_dcpl_30 = or_dcpl_27 | or_dcpl_11;
  assign or_dcpl_34 = or_dcpl_16 | or_dcpl_21;
  assign or_dcpl_36 = or_dcpl_22 | or_dcpl_11;
  assign or_dcpl_40 = or_dcpl_12 | or_dcpl_21;
  assign or_dcpl_42 = (MAC_LOOP_n_6_0_sva[4:3]!=2'b10);
  assign or_dcpl_43 = or_dcpl_12 | or_dcpl_42;
  assign or_dcpl_47 = (MAC_LOOP_n_6_0_sva[4:3]!=2'b01);
  assign or_dcpl_48 = or_dcpl_22 | or_dcpl_47;
  assign or_dcpl_50 = or_dcpl_16 | or_dcpl_42;
  assign or_dcpl_54 = or_dcpl_27 | or_dcpl_47;
  assign or_dcpl_56 = or_dcpl_27 | or_dcpl_42;
  assign or_dcpl_60 = or_dcpl_16 | or_dcpl_47;
  assign or_dcpl_62 = or_dcpl_22 | or_dcpl_42;
  assign or_dcpl_66 = or_dcpl_12 | or_dcpl_47;
  assign or_dcpl_100 = (MAC_LOOP_n_6_0_sva[6:5]!=2'b10);
  assign or_dcpl_101 = or_dcpl_100 | (~ (MAC_LOOP_n_6_0_sva[0]));
  assign or_dcpl_104 = or_dcpl_100 | (MAC_LOOP_n_6_0_sva[0]);
  assign or_dcpl_106 = (MAC_LOOP_n_6_0_sva[6:5]!=2'b01);
  assign or_dcpl_107 = or_dcpl_106 | (MAC_LOOP_n_6_0_sva[0]);
  assign or_dcpl_110 = or_dcpl_106 | (~ (MAC_LOOP_n_6_0_sva[0]));
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_0 <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      y_rsci_idat_0 <= (z_out_3[0]) | nor_ovfl_sva_1 | and_unfl_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_7_1 <= 7'b0000000;
    end
    else if ( fsm_output[3] ) begin
      y_rsci_idat_7_1 <= ~(MUX_v_7_2_2(nor_5_nl, 7'b1111111, and_unfl_sva_1));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_8 <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      y_rsci_idat_8 <= z_out_3[14];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_sample_sva <= 3'b000;
    end
    else if ( ~((fsm_output[2:1]!=2'b00)) ) begin
      i_sample_sva <= i_sample_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_126_lpi_2 <= 3'b000;
    end
    else if ( ~(or_dcpl_13 | or_dcpl_10 | (fsm_output[2])) ) begin
      x_126_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_125_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_17 | or_dcpl_15) ) begin
      x_125_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_1_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_23 | or_dcpl_20) ) begin
      x_1_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_124_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_17 | or_dcpl_10) ) begin
      x_124_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_2_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_28 | or_dcpl_26) ) begin
      x_2_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_123_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_30 | or_dcpl_15) ) begin
      x_123_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_3_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_28 | or_dcpl_20) ) begin
      x_3_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_122_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_30 | or_dcpl_10) ) begin
      x_122_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_4_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_34 | or_dcpl_26) ) begin
      x_4_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_121_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_36 | or_dcpl_15) ) begin
      x_121_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_5_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_34 | or_dcpl_20) ) begin
      x_5_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_120_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_36 | or_dcpl_10) ) begin
      x_120_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_6_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_40 | or_dcpl_26) ) begin
      x_6_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_119_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_43 | or_dcpl_15) ) begin
      x_119_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_7_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_40 | or_dcpl_20) ) begin
      x_7_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_118_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_43 | or_dcpl_10) ) begin
      x_118_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_8_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_48 | or_dcpl_26) ) begin
      x_8_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_117_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_50 | or_dcpl_15) ) begin
      x_117_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_9_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_48 | or_dcpl_20) ) begin
      x_9_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_116_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_50 | or_dcpl_10) ) begin
      x_116_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_10_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_54 | or_dcpl_26) ) begin
      x_10_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_115_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_56 | or_dcpl_15) ) begin
      x_115_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_11_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_54 | or_dcpl_20) ) begin
      x_11_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_114_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_56 | or_dcpl_10) ) begin
      x_114_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_12_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_60 | or_dcpl_26) ) begin
      x_12_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_113_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_62 | or_dcpl_15) ) begin
      x_113_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_13_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_60 | or_dcpl_20) ) begin
      x_13_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_112_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_62 | or_dcpl_10) ) begin
      x_112_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_14_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_66 | or_dcpl_26) ) begin
      x_14_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_111_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_66 | or_dcpl_15) ) begin
      x_111_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_15_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_66 | or_dcpl_20) ) begin
      x_15_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_110_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_66 | or_dcpl_10) ) begin
      x_110_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_16_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_62 | or_dcpl_26) ) begin
      x_16_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_109_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_60 | or_dcpl_15) ) begin
      x_109_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_17_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_62 | or_dcpl_20) ) begin
      x_17_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_108_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_60 | or_dcpl_10) ) begin
      x_108_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_18_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_56 | or_dcpl_26) ) begin
      x_18_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_107_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_54 | or_dcpl_15) ) begin
      x_107_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_19_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_56 | or_dcpl_20) ) begin
      x_19_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_106_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_54 | or_dcpl_10) ) begin
      x_106_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_20_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_50 | or_dcpl_26) ) begin
      x_20_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_105_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_48 | or_dcpl_15) ) begin
      x_105_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_21_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_50 | or_dcpl_20) ) begin
      x_21_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_104_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_48 | or_dcpl_10) ) begin
      x_104_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_22_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_43 | or_dcpl_26) ) begin
      x_22_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_103_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_40 | or_dcpl_15) ) begin
      x_103_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_23_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_43 | or_dcpl_20) ) begin
      x_23_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_102_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_40 | or_dcpl_10) ) begin
      x_102_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_24_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_36 | or_dcpl_26) ) begin
      x_24_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_101_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_34 | or_dcpl_15) ) begin
      x_101_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_25_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_36 | or_dcpl_20) ) begin
      x_25_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_100_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_34 | or_dcpl_10) ) begin
      x_100_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_26_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_30 | or_dcpl_26) ) begin
      x_26_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_99_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_28 | or_dcpl_15) ) begin
      x_99_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_27_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_30 | or_dcpl_20) ) begin
      x_27_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_98_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_28 | or_dcpl_10) ) begin
      x_98_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_28_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_17 | or_dcpl_26) ) begin
      x_28_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_97_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_23 | or_dcpl_15) ) begin
      x_97_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_29_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_17 | or_dcpl_20) ) begin
      x_29_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_96_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_23 | or_dcpl_10) ) begin
      x_96_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_30_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_13 | or_dcpl_26) ) begin
      x_30_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_95_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_13 | or_dcpl_101) ) begin
      x_95_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_31_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_13 | or_dcpl_20) ) begin
      x_31_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_94_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_13 | or_dcpl_104) ) begin
      x_94_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_32_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_23 | or_dcpl_107) ) begin
      x_32_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_93_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_17 | or_dcpl_101) ) begin
      x_93_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_33_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_23 | or_dcpl_110) ) begin
      x_33_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_92_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_17 | or_dcpl_104) ) begin
      x_92_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_34_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_28 | or_dcpl_107) ) begin
      x_34_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_91_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_30 | or_dcpl_101) ) begin
      x_91_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_35_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_28 | or_dcpl_110) ) begin
      x_35_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_90_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_30 | or_dcpl_104) ) begin
      x_90_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_36_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_34 | or_dcpl_107) ) begin
      x_36_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_89_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_36 | or_dcpl_101) ) begin
      x_89_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_37_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_34 | or_dcpl_110) ) begin
      x_37_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_88_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_36 | or_dcpl_104) ) begin
      x_88_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_38_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_40 | or_dcpl_107) ) begin
      x_38_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_87_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_43 | or_dcpl_101) ) begin
      x_87_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_39_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_40 | or_dcpl_110) ) begin
      x_39_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_86_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_43 | or_dcpl_104) ) begin
      x_86_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_40_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_48 | or_dcpl_107) ) begin
      x_40_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_85_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_50 | or_dcpl_101) ) begin
      x_85_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_41_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_48 | or_dcpl_110) ) begin
      x_41_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_84_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_50 | or_dcpl_104) ) begin
      x_84_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_42_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_54 | or_dcpl_107) ) begin
      x_42_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_83_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_56 | or_dcpl_101) ) begin
      x_83_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_43_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_54 | or_dcpl_110) ) begin
      x_43_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_82_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_56 | or_dcpl_104) ) begin
      x_82_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_44_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_60 | or_dcpl_107) ) begin
      x_44_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_81_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_62 | or_dcpl_101) ) begin
      x_81_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_45_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_60 | or_dcpl_110) ) begin
      x_45_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_80_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_62 | or_dcpl_104) ) begin
      x_80_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_46_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_66 | or_dcpl_107) ) begin
      x_46_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_79_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_66 | or_dcpl_101) ) begin
      x_79_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_47_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_66 | or_dcpl_110) ) begin
      x_47_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_78_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_66 | or_dcpl_104) ) begin
      x_78_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_48_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_62 | or_dcpl_107) ) begin
      x_48_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_77_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_60 | or_dcpl_101) ) begin
      x_77_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_49_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_62 | or_dcpl_110) ) begin
      x_49_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_76_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_60 | or_dcpl_104) ) begin
      x_76_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_50_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_56 | or_dcpl_107) ) begin
      x_50_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_75_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_54 | or_dcpl_101) ) begin
      x_75_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_51_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_56 | or_dcpl_110) ) begin
      x_51_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_74_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_54 | or_dcpl_104) ) begin
      x_74_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_52_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_50 | or_dcpl_107) ) begin
      x_52_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_73_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_48 | or_dcpl_101) ) begin
      x_73_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_53_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_50 | or_dcpl_110) ) begin
      x_53_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_72_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_48 | or_dcpl_104) ) begin
      x_72_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_54_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_43 | or_dcpl_107) ) begin
      x_54_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_71_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_40 | or_dcpl_101) ) begin
      x_71_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_55_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_43 | or_dcpl_110) ) begin
      x_55_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_70_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_40 | or_dcpl_104) ) begin
      x_70_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_56_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_36 | or_dcpl_107) ) begin
      x_56_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_69_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_34 | or_dcpl_101) ) begin
      x_69_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_57_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_36 | or_dcpl_110) ) begin
      x_57_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_68_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_34 | or_dcpl_104) ) begin
      x_68_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_58_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_30 | or_dcpl_107) ) begin
      x_58_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_67_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_28 | or_dcpl_101) ) begin
      x_67_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_59_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_30 | or_dcpl_110) ) begin
      x_59_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_66_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_28 | or_dcpl_104) ) begin
      x_66_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_60_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_17 | or_dcpl_107) ) begin
      x_60_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_65_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_23 | or_dcpl_101) ) begin
      x_65_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_61_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_17 | or_dcpl_110) ) begin
      x_61_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_64_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_23 | or_dcpl_104) ) begin
      x_64_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_62_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_13 | or_dcpl_107) ) begin
      x_62_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_63_lpi_2 <= 3'b000;
    end
    else if ( ~((~ (fsm_output[1])) | or_dcpl_13 | or_dcpl_110) ) begin
      x_63_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_0_sva <= 3'b000;
    end
    else if ( fsm_output[2] ) begin
      x_0_sva <= i_sample_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsc_triosy_obj_ld <= 1'b0;
      reg_b_rsc_triosy_obj_ld_cse <= 1'b0;
      MAC_LOOP_n_6_0_sva <= 7'b0000000;
      sum_sva <= 20'b00000000000000000000;
    end
    else begin
      y_rsc_triosy_obj_ld <= fsm_output[3];
      reg_b_rsc_triosy_obj_ld_cse <= (~ z_out_1_7) & (fsm_output[2]);
      MAC_LOOP_n_6_0_sva <= MUX_v_7_2_2(7'b0000000, SHIFT_LOOP_n_SHIFT_LOOP_n_mux_nl,
          MAC_LOOP_n_nor_nl);
      sum_sva <= MUX_v_20_2_2(20'b00000000000000000000, z_out_3, (fsm_output[2]));
    end
  end
  assign nor_5_nl = ~(MUX_v_7_2_2((z_out_3[7:1]), 7'b1111111, nor_ovfl_sva_1));
  assign SHIFT_LOOP_n_or_nl = (z_out_1_7 & (fsm_output[1])) | (fsm_output[2]);
  assign SHIFT_LOOP_n_SHIFT_LOOP_n_mux_nl = MUX_v_7_2_2(7'b1111110, z_out_2, SHIFT_LOOP_n_or_nl);
  assign MAC_LOOP_n_nor_nl = ~((fsm_output[4:3]!=2'b00) | ((~ z_out_1_7) & (fsm_output[1])));
  assign SHIFT_LOOP_mux_129_nl = MUX_v_7_2_2((~ z_out_2), z_out_2, fsm_output[2]);
  assign nl_SHIFT_LOOP_acc_nl = ({1'b1 , SHIFT_LOOP_mux_129_nl}) + 8'b00000001;
  assign SHIFT_LOOP_acc_nl = nl_SHIFT_LOOP_acc_nl[7:0];
  assign z_out_1_7 = readslicef_8_1_7(SHIFT_LOOP_acc_nl);
  assign nl_z_out_2 = MAC_LOOP_n_6_0_sva + conv_s2u_2_7({(fsm_output[1]) , 1'b1});
  assign z_out_2 = nl_z_out_2[6:0];
  assign MAC_LOOP_mux_7_nl = MUX_v_19_2_2((sum_sva[18:0]), (signext_19_14(sum_sva[19:6])),
      fsm_output[3]);
  assign MAC_LOOP_mux_9_nl = MUX_v_10_127_2((b_rsci_idat[9:0]), (b_rsci_idat[19:10]),
      (b_rsci_idat[29:20]), (b_rsci_idat[39:30]), (b_rsci_idat[49:40]), (b_rsci_idat[59:50]),
      (b_rsci_idat[69:60]), (b_rsci_idat[79:70]), (b_rsci_idat[89:80]), (b_rsci_idat[99:90]),
      (b_rsci_idat[109:100]), (b_rsci_idat[119:110]), (b_rsci_idat[129:120]), (b_rsci_idat[139:130]),
      (b_rsci_idat[149:140]), (b_rsci_idat[159:150]), (b_rsci_idat[169:160]), (b_rsci_idat[179:170]),
      (b_rsci_idat[189:180]), (b_rsci_idat[199:190]), (b_rsci_idat[209:200]), (b_rsci_idat[219:210]),
      (b_rsci_idat[229:220]), (b_rsci_idat[239:230]), (b_rsci_idat[249:240]), (b_rsci_idat[259:250]),
      (b_rsci_idat[269:260]), (b_rsci_idat[279:270]), (b_rsci_idat[289:280]), (b_rsci_idat[299:290]),
      (b_rsci_idat[309:300]), (b_rsci_idat[319:310]), (b_rsci_idat[329:320]), (b_rsci_idat[339:330]),
      (b_rsci_idat[349:340]), (b_rsci_idat[359:350]), (b_rsci_idat[369:360]), (b_rsci_idat[379:370]),
      (b_rsci_idat[389:380]), (b_rsci_idat[399:390]), (b_rsci_idat[409:400]), (b_rsci_idat[419:410]),
      (b_rsci_idat[429:420]), (b_rsci_idat[439:430]), (b_rsci_idat[449:440]), (b_rsci_idat[459:450]),
      (b_rsci_idat[469:460]), (b_rsci_idat[479:470]), (b_rsci_idat[489:480]), (b_rsci_idat[499:490]),
      (b_rsci_idat[509:500]), (b_rsci_idat[519:510]), (b_rsci_idat[529:520]), (b_rsci_idat[539:530]),
      (b_rsci_idat[549:540]), (b_rsci_idat[559:550]), (b_rsci_idat[569:560]), (b_rsci_idat[579:570]),
      (b_rsci_idat[589:580]), (b_rsci_idat[599:590]), (b_rsci_idat[609:600]), (b_rsci_idat[619:610]),
      (b_rsci_idat[629:620]), (b_rsci_idat[639:630]), (b_rsci_idat[649:640]), (b_rsci_idat[659:650]),
      (b_rsci_idat[669:660]), (b_rsci_idat[679:670]), (b_rsci_idat[689:680]), (b_rsci_idat[699:690]),
      (b_rsci_idat[709:700]), (b_rsci_idat[719:710]), (b_rsci_idat[729:720]), (b_rsci_idat[739:730]),
      (b_rsci_idat[749:740]), (b_rsci_idat[759:750]), (b_rsci_idat[769:760]), (b_rsci_idat[779:770]),
      (b_rsci_idat[789:780]), (b_rsci_idat[799:790]), (b_rsci_idat[809:800]), (b_rsci_idat[819:810]),
      (b_rsci_idat[829:820]), (b_rsci_idat[839:830]), (b_rsci_idat[849:840]), (b_rsci_idat[859:850]),
      (b_rsci_idat[869:860]), (b_rsci_idat[879:870]), (b_rsci_idat[889:880]), (b_rsci_idat[899:890]),
      (b_rsci_idat[909:900]), (b_rsci_idat[919:910]), (b_rsci_idat[929:920]), (b_rsci_idat[939:930]),
      (b_rsci_idat[949:940]), (b_rsci_idat[959:950]), (b_rsci_idat[969:960]), (b_rsci_idat[979:970]),
      (b_rsci_idat[989:980]), (b_rsci_idat[999:990]), (b_rsci_idat[1009:1000]), (b_rsci_idat[1019:1010]),
      (b_rsci_idat[1029:1020]), (b_rsci_idat[1039:1030]), (b_rsci_idat[1049:1040]),
      (b_rsci_idat[1059:1050]), (b_rsci_idat[1069:1060]), (b_rsci_idat[1079:1070]),
      (b_rsci_idat[1089:1080]), (b_rsci_idat[1099:1090]), (b_rsci_idat[1109:1100]),
      (b_rsci_idat[1119:1110]), (b_rsci_idat[1129:1120]), (b_rsci_idat[1139:1130]),
      (b_rsci_idat[1149:1140]), (b_rsci_idat[1159:1150]), (b_rsci_idat[1169:1160]),
      (b_rsci_idat[1179:1170]), (b_rsci_idat[1189:1180]), (b_rsci_idat[1199:1190]),
      (b_rsci_idat[1209:1200]), (b_rsci_idat[1219:1210]), (b_rsci_idat[1229:1220]),
      (b_rsci_idat[1239:1230]), (b_rsci_idat[1249:1240]), (b_rsci_idat[1259:1250]),
      (b_rsci_idat[1269:1260]), MAC_LOOP_n_6_0_sva);
  assign MAC_LOOP_mul_1_nl = conv_s2u_13_13($signed(z_out) * $signed(MAC_LOOP_mux_9_nl));
  assign MAC_LOOP_mux_8_nl = MUX_v_13_2_2(MAC_LOOP_mul_1_nl, ({12'b000000000000 ,
      (sum_sva[5])}), fsm_output[3]);
  assign nl_z_out_3 = ({(sum_sva[19]) , MAC_LOOP_mux_7_nl}) + conv_s2u_13_20(MAC_LOOP_mux_8_nl);
  assign z_out_3 = nl_z_out_3[19:0];
  assign MAC_LOOP_mux_10_nl = MUX_v_3_2_2(i_sample_sva, x_0_sva, fsm_output[1]);
  assign MAC_LOOP_mux_11_nl = MUX_v_7_2_2(MAC_LOOP_n_6_0_sva, z_out_2, fsm_output[1]);
  assign z_out = MUX_v_3_127_2(MAC_LOOP_mux_10_nl, x_1_lpi_2, x_2_lpi_2, x_3_lpi_2,
      x_4_lpi_2, x_5_lpi_2, x_6_lpi_2, x_7_lpi_2, x_8_lpi_2, x_9_lpi_2, x_10_lpi_2,
      x_11_lpi_2, x_12_lpi_2, x_13_lpi_2, x_14_lpi_2, x_15_lpi_2, x_16_lpi_2, x_17_lpi_2,
      x_18_lpi_2, x_19_lpi_2, x_20_lpi_2, x_21_lpi_2, x_22_lpi_2, x_23_lpi_2, x_24_lpi_2,
      x_25_lpi_2, x_26_lpi_2, x_27_lpi_2, x_28_lpi_2, x_29_lpi_2, x_30_lpi_2, x_31_lpi_2,
      x_32_lpi_2, x_33_lpi_2, x_34_lpi_2, x_35_lpi_2, x_36_lpi_2, x_37_lpi_2, x_38_lpi_2,
      x_39_lpi_2, x_40_lpi_2, x_41_lpi_2, x_42_lpi_2, x_43_lpi_2, x_44_lpi_2, x_45_lpi_2,
      x_46_lpi_2, x_47_lpi_2, x_48_lpi_2, x_49_lpi_2, x_50_lpi_2, x_51_lpi_2, x_52_lpi_2,
      x_53_lpi_2, x_54_lpi_2, x_55_lpi_2, x_56_lpi_2, x_57_lpi_2, x_58_lpi_2, x_59_lpi_2,
      x_60_lpi_2, x_61_lpi_2, x_62_lpi_2, x_63_lpi_2, x_64_lpi_2, x_65_lpi_2, x_66_lpi_2,
      x_67_lpi_2, x_68_lpi_2, x_69_lpi_2, x_70_lpi_2, x_71_lpi_2, x_72_lpi_2, x_73_lpi_2,
      x_74_lpi_2, x_75_lpi_2, x_76_lpi_2, x_77_lpi_2, x_78_lpi_2, x_79_lpi_2, x_80_lpi_2,
      x_81_lpi_2, x_82_lpi_2, x_83_lpi_2, x_84_lpi_2, x_85_lpi_2, x_86_lpi_2, x_87_lpi_2,
      x_88_lpi_2, x_89_lpi_2, x_90_lpi_2, x_91_lpi_2, x_92_lpi_2, x_93_lpi_2, x_94_lpi_2,
      x_95_lpi_2, x_96_lpi_2, x_97_lpi_2, x_98_lpi_2, x_99_lpi_2, x_100_lpi_2, x_101_lpi_2,
      x_102_lpi_2, x_103_lpi_2, x_104_lpi_2, x_105_lpi_2, x_106_lpi_2, x_107_lpi_2,
      x_108_lpi_2, x_109_lpi_2, x_110_lpi_2, x_111_lpi_2, x_112_lpi_2, x_113_lpi_2,
      x_114_lpi_2, x_115_lpi_2, x_116_lpi_2, x_117_lpi_2, x_118_lpi_2, x_119_lpi_2,
      x_120_lpi_2, x_121_lpi_2, x_122_lpi_2, x_123_lpi_2, x_124_lpi_2, x_125_lpi_2,
      x_126_lpi_2, MAC_LOOP_mux_11_nl);

  function automatic [9:0] MUX_v_10_127_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [9:0] input_8;
    input [9:0] input_9;
    input [9:0] input_10;
    input [9:0] input_11;
    input [9:0] input_12;
    input [9:0] input_13;
    input [9:0] input_14;
    input [9:0] input_15;
    input [9:0] input_16;
    input [9:0] input_17;
    input [9:0] input_18;
    input [9:0] input_19;
    input [9:0] input_20;
    input [9:0] input_21;
    input [9:0] input_22;
    input [9:0] input_23;
    input [9:0] input_24;
    input [9:0] input_25;
    input [9:0] input_26;
    input [9:0] input_27;
    input [9:0] input_28;
    input [9:0] input_29;
    input [9:0] input_30;
    input [9:0] input_31;
    input [9:0] input_32;
    input [9:0] input_33;
    input [9:0] input_34;
    input [9:0] input_35;
    input [9:0] input_36;
    input [9:0] input_37;
    input [9:0] input_38;
    input [9:0] input_39;
    input [9:0] input_40;
    input [9:0] input_41;
    input [9:0] input_42;
    input [9:0] input_43;
    input [9:0] input_44;
    input [9:0] input_45;
    input [9:0] input_46;
    input [9:0] input_47;
    input [9:0] input_48;
    input [9:0] input_49;
    input [9:0] input_50;
    input [9:0] input_51;
    input [9:0] input_52;
    input [9:0] input_53;
    input [9:0] input_54;
    input [9:0] input_55;
    input [9:0] input_56;
    input [9:0] input_57;
    input [9:0] input_58;
    input [9:0] input_59;
    input [9:0] input_60;
    input [9:0] input_61;
    input [9:0] input_62;
    input [9:0] input_63;
    input [9:0] input_64;
    input [9:0] input_65;
    input [9:0] input_66;
    input [9:0] input_67;
    input [9:0] input_68;
    input [9:0] input_69;
    input [9:0] input_70;
    input [9:0] input_71;
    input [9:0] input_72;
    input [9:0] input_73;
    input [9:0] input_74;
    input [9:0] input_75;
    input [9:0] input_76;
    input [9:0] input_77;
    input [9:0] input_78;
    input [9:0] input_79;
    input [9:0] input_80;
    input [9:0] input_81;
    input [9:0] input_82;
    input [9:0] input_83;
    input [9:0] input_84;
    input [9:0] input_85;
    input [9:0] input_86;
    input [9:0] input_87;
    input [9:0] input_88;
    input [9:0] input_89;
    input [9:0] input_90;
    input [9:0] input_91;
    input [9:0] input_92;
    input [9:0] input_93;
    input [9:0] input_94;
    input [9:0] input_95;
    input [9:0] input_96;
    input [9:0] input_97;
    input [9:0] input_98;
    input [9:0] input_99;
    input [9:0] input_100;
    input [9:0] input_101;
    input [9:0] input_102;
    input [9:0] input_103;
    input [9:0] input_104;
    input [9:0] input_105;
    input [9:0] input_106;
    input [9:0] input_107;
    input [9:0] input_108;
    input [9:0] input_109;
    input [9:0] input_110;
    input [9:0] input_111;
    input [9:0] input_112;
    input [9:0] input_113;
    input [9:0] input_114;
    input [9:0] input_115;
    input [9:0] input_116;
    input [9:0] input_117;
    input [9:0] input_118;
    input [9:0] input_119;
    input [9:0] input_120;
    input [9:0] input_121;
    input [9:0] input_122;
    input [9:0] input_123;
    input [9:0] input_124;
    input [9:0] input_125;
    input [9:0] input_126;
    input [6:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      7'b1000001 : begin
        result = input_65;
      end
      7'b1000010 : begin
        result = input_66;
      end
      7'b1000011 : begin
        result = input_67;
      end
      7'b1000100 : begin
        result = input_68;
      end
      7'b1000101 : begin
        result = input_69;
      end
      7'b1000110 : begin
        result = input_70;
      end
      7'b1000111 : begin
        result = input_71;
      end
      7'b1001000 : begin
        result = input_72;
      end
      7'b1001001 : begin
        result = input_73;
      end
      7'b1001010 : begin
        result = input_74;
      end
      7'b1001011 : begin
        result = input_75;
      end
      7'b1001100 : begin
        result = input_76;
      end
      7'b1001101 : begin
        result = input_77;
      end
      7'b1001110 : begin
        result = input_78;
      end
      7'b1001111 : begin
        result = input_79;
      end
      7'b1010000 : begin
        result = input_80;
      end
      7'b1010001 : begin
        result = input_81;
      end
      7'b1010010 : begin
        result = input_82;
      end
      7'b1010011 : begin
        result = input_83;
      end
      7'b1010100 : begin
        result = input_84;
      end
      7'b1010101 : begin
        result = input_85;
      end
      7'b1010110 : begin
        result = input_86;
      end
      7'b1010111 : begin
        result = input_87;
      end
      7'b1011000 : begin
        result = input_88;
      end
      7'b1011001 : begin
        result = input_89;
      end
      7'b1011010 : begin
        result = input_90;
      end
      7'b1011011 : begin
        result = input_91;
      end
      7'b1011100 : begin
        result = input_92;
      end
      7'b1011101 : begin
        result = input_93;
      end
      7'b1011110 : begin
        result = input_94;
      end
      7'b1011111 : begin
        result = input_95;
      end
      7'b1100000 : begin
        result = input_96;
      end
      7'b1100001 : begin
        result = input_97;
      end
      7'b1100010 : begin
        result = input_98;
      end
      7'b1100011 : begin
        result = input_99;
      end
      7'b1100100 : begin
        result = input_100;
      end
      7'b1100101 : begin
        result = input_101;
      end
      7'b1100110 : begin
        result = input_102;
      end
      7'b1100111 : begin
        result = input_103;
      end
      7'b1101000 : begin
        result = input_104;
      end
      7'b1101001 : begin
        result = input_105;
      end
      7'b1101010 : begin
        result = input_106;
      end
      7'b1101011 : begin
        result = input_107;
      end
      7'b1101100 : begin
        result = input_108;
      end
      7'b1101101 : begin
        result = input_109;
      end
      7'b1101110 : begin
        result = input_110;
      end
      7'b1101111 : begin
        result = input_111;
      end
      7'b1110000 : begin
        result = input_112;
      end
      7'b1110001 : begin
        result = input_113;
      end
      7'b1110010 : begin
        result = input_114;
      end
      7'b1110011 : begin
        result = input_115;
      end
      7'b1110100 : begin
        result = input_116;
      end
      7'b1110101 : begin
        result = input_117;
      end
      7'b1110110 : begin
        result = input_118;
      end
      7'b1110111 : begin
        result = input_119;
      end
      7'b1111000 : begin
        result = input_120;
      end
      7'b1111001 : begin
        result = input_121;
      end
      7'b1111010 : begin
        result = input_122;
      end
      7'b1111011 : begin
        result = input_123;
      end
      7'b1111100 : begin
        result = input_124;
      end
      7'b1111101 : begin
        result = input_125;
      end
      default : begin
        result = input_126;
      end
    endcase
    MUX_v_10_127_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input [0:0] sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [18:0] MUX_v_19_2_2;
    input [18:0] input_0;
    input [18:0] input_1;
    input [0:0] sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_127_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] input_8;
    input [2:0] input_9;
    input [2:0] input_10;
    input [2:0] input_11;
    input [2:0] input_12;
    input [2:0] input_13;
    input [2:0] input_14;
    input [2:0] input_15;
    input [2:0] input_16;
    input [2:0] input_17;
    input [2:0] input_18;
    input [2:0] input_19;
    input [2:0] input_20;
    input [2:0] input_21;
    input [2:0] input_22;
    input [2:0] input_23;
    input [2:0] input_24;
    input [2:0] input_25;
    input [2:0] input_26;
    input [2:0] input_27;
    input [2:0] input_28;
    input [2:0] input_29;
    input [2:0] input_30;
    input [2:0] input_31;
    input [2:0] input_32;
    input [2:0] input_33;
    input [2:0] input_34;
    input [2:0] input_35;
    input [2:0] input_36;
    input [2:0] input_37;
    input [2:0] input_38;
    input [2:0] input_39;
    input [2:0] input_40;
    input [2:0] input_41;
    input [2:0] input_42;
    input [2:0] input_43;
    input [2:0] input_44;
    input [2:0] input_45;
    input [2:0] input_46;
    input [2:0] input_47;
    input [2:0] input_48;
    input [2:0] input_49;
    input [2:0] input_50;
    input [2:0] input_51;
    input [2:0] input_52;
    input [2:0] input_53;
    input [2:0] input_54;
    input [2:0] input_55;
    input [2:0] input_56;
    input [2:0] input_57;
    input [2:0] input_58;
    input [2:0] input_59;
    input [2:0] input_60;
    input [2:0] input_61;
    input [2:0] input_62;
    input [2:0] input_63;
    input [2:0] input_64;
    input [2:0] input_65;
    input [2:0] input_66;
    input [2:0] input_67;
    input [2:0] input_68;
    input [2:0] input_69;
    input [2:0] input_70;
    input [2:0] input_71;
    input [2:0] input_72;
    input [2:0] input_73;
    input [2:0] input_74;
    input [2:0] input_75;
    input [2:0] input_76;
    input [2:0] input_77;
    input [2:0] input_78;
    input [2:0] input_79;
    input [2:0] input_80;
    input [2:0] input_81;
    input [2:0] input_82;
    input [2:0] input_83;
    input [2:0] input_84;
    input [2:0] input_85;
    input [2:0] input_86;
    input [2:0] input_87;
    input [2:0] input_88;
    input [2:0] input_89;
    input [2:0] input_90;
    input [2:0] input_91;
    input [2:0] input_92;
    input [2:0] input_93;
    input [2:0] input_94;
    input [2:0] input_95;
    input [2:0] input_96;
    input [2:0] input_97;
    input [2:0] input_98;
    input [2:0] input_99;
    input [2:0] input_100;
    input [2:0] input_101;
    input [2:0] input_102;
    input [2:0] input_103;
    input [2:0] input_104;
    input [2:0] input_105;
    input [2:0] input_106;
    input [2:0] input_107;
    input [2:0] input_108;
    input [2:0] input_109;
    input [2:0] input_110;
    input [2:0] input_111;
    input [2:0] input_112;
    input [2:0] input_113;
    input [2:0] input_114;
    input [2:0] input_115;
    input [2:0] input_116;
    input [2:0] input_117;
    input [2:0] input_118;
    input [2:0] input_119;
    input [2:0] input_120;
    input [2:0] input_121;
    input [2:0] input_122;
    input [2:0] input_123;
    input [2:0] input_124;
    input [2:0] input_125;
    input [2:0] input_126;
    input [6:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      7'b1000001 : begin
        result = input_65;
      end
      7'b1000010 : begin
        result = input_66;
      end
      7'b1000011 : begin
        result = input_67;
      end
      7'b1000100 : begin
        result = input_68;
      end
      7'b1000101 : begin
        result = input_69;
      end
      7'b1000110 : begin
        result = input_70;
      end
      7'b1000111 : begin
        result = input_71;
      end
      7'b1001000 : begin
        result = input_72;
      end
      7'b1001001 : begin
        result = input_73;
      end
      7'b1001010 : begin
        result = input_74;
      end
      7'b1001011 : begin
        result = input_75;
      end
      7'b1001100 : begin
        result = input_76;
      end
      7'b1001101 : begin
        result = input_77;
      end
      7'b1001110 : begin
        result = input_78;
      end
      7'b1001111 : begin
        result = input_79;
      end
      7'b1010000 : begin
        result = input_80;
      end
      7'b1010001 : begin
        result = input_81;
      end
      7'b1010010 : begin
        result = input_82;
      end
      7'b1010011 : begin
        result = input_83;
      end
      7'b1010100 : begin
        result = input_84;
      end
      7'b1010101 : begin
        result = input_85;
      end
      7'b1010110 : begin
        result = input_86;
      end
      7'b1010111 : begin
        result = input_87;
      end
      7'b1011000 : begin
        result = input_88;
      end
      7'b1011001 : begin
        result = input_89;
      end
      7'b1011010 : begin
        result = input_90;
      end
      7'b1011011 : begin
        result = input_91;
      end
      7'b1011100 : begin
        result = input_92;
      end
      7'b1011101 : begin
        result = input_93;
      end
      7'b1011110 : begin
        result = input_94;
      end
      7'b1011111 : begin
        result = input_95;
      end
      7'b1100000 : begin
        result = input_96;
      end
      7'b1100001 : begin
        result = input_97;
      end
      7'b1100010 : begin
        result = input_98;
      end
      7'b1100011 : begin
        result = input_99;
      end
      7'b1100100 : begin
        result = input_100;
      end
      7'b1100101 : begin
        result = input_101;
      end
      7'b1100110 : begin
        result = input_102;
      end
      7'b1100111 : begin
        result = input_103;
      end
      7'b1101000 : begin
        result = input_104;
      end
      7'b1101001 : begin
        result = input_105;
      end
      7'b1101010 : begin
        result = input_106;
      end
      7'b1101011 : begin
        result = input_107;
      end
      7'b1101100 : begin
        result = input_108;
      end
      7'b1101101 : begin
        result = input_109;
      end
      7'b1101110 : begin
        result = input_110;
      end
      7'b1101111 : begin
        result = input_111;
      end
      7'b1110000 : begin
        result = input_112;
      end
      7'b1110001 : begin
        result = input_113;
      end
      7'b1110010 : begin
        result = input_114;
      end
      7'b1110011 : begin
        result = input_115;
      end
      7'b1110100 : begin
        result = input_116;
      end
      7'b1110101 : begin
        result = input_117;
      end
      7'b1110110 : begin
        result = input_118;
      end
      7'b1110111 : begin
        result = input_119;
      end
      7'b1111000 : begin
        result = input_120;
      end
      7'b1111001 : begin
        result = input_121;
      end
      7'b1111010 : begin
        result = input_122;
      end
      7'b1111011 : begin
        result = input_123;
      end
      7'b1111100 : begin
        result = input_124;
      end
      7'b1111101 : begin
        result = input_125;
      end
      default : begin
        result = input_126;
      end
    endcase
    MUX_v_3_127_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] signext_19_14;
    input [13:0] vector;
  begin
    signext_19_14= {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [6:0] conv_s2u_2_7 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_7 = {{5{vector[1]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_13_13 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_13 = vector;
  end
  endfunction


  function automatic [19:0] conv_s2u_13_20 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_20 = {{7{vector[12]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_filter
// ------------------------------------------------------------------


module fir_filter (
  clk, rst, i_sample_rsc_dat, i_sample_rsc_triosy_lz, b_rsc_dat, b_rsc_triosy_lz,
      y_rsc_dat, y_rsc_triosy_lz
);
  input clk;
  input rst;
  input [2:0] i_sample_rsc_dat;
  output i_sample_rsc_triosy_lz;
  input [1269:0] b_rsc_dat;
  output b_rsc_triosy_lz;
  output [8:0] y_rsc_dat;
  output y_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  fir_filter_core fir_filter_core_inst (
      .clk(clk),
      .rst(rst),
      .i_sample_rsc_dat(i_sample_rsc_dat),
      .i_sample_rsc_triosy_lz(i_sample_rsc_triosy_lz),
      .b_rsc_dat(b_rsc_dat),
      .b_rsc_triosy_lz(b_rsc_triosy_lz),
      .y_rsc_dat(y_rsc_dat),
      .y_rsc_triosy_lz(y_rsc_triosy_lz)
    );
endmodule



