
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_out_dreg_pkg_v2 IS

COMPONENT mgc_out_dreg_v2
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_out_dreg_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_out_dreg_v2 IS
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    d        : IN  std_logic_vector(width-1 DOWNTO 0);
    z        : OUT std_logic_vector(width-1 DOWNTO 0)
  );
END mgc_out_dreg_v2;

ARCHITECTURE beh OF mgc_out_dreg_v2 IS
BEGIN

  z <= d;

END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_rem IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END mgc_rem;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_rem IS
BEGIN
  z <= std_logic_vector(unsigned(a) rem unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) rem   signed(b));
END beh;

--------> ../td_ccore_solutions/modulo_dev_bb61c76201db0c9669a47462bb7d006361ff_0/rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Tue Jul 20 15:24:30 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    modulo_dev_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_dev_core IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_dev_core;

ARCHITECTURE v1 OF modulo_dev_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL base_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat : STD_LOGIC;
  SIGNAL rem_13_cmp_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_1_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_2_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_3_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_4_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_5_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_6_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_7_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_8_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_9_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_10_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_11_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_1_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_2_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_3_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_4_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_5_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_6_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_7_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_8_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_9_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_10_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_11_b_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_1_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_2_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_3_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_4_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_5_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_6_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_7_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_8_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_9_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_10_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_13_cmp_11_a_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL acc_tmp : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL acc_1_tmp : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_dcpl_1 : STD_LOGIC;
  SIGNAL and_dcpl_2 : STD_LOGIC;
  SIGNAL and_dcpl_3 : STD_LOGIC;
  SIGNAL and_dcpl_4 : STD_LOGIC;
  SIGNAL and_dcpl_6 : STD_LOGIC;
  SIGNAL and_dcpl_8 : STD_LOGIC;
  SIGNAL and_dcpl_9 : STD_LOGIC;
  SIGNAL and_dcpl_11 : STD_LOGIC;
  SIGNAL and_dcpl_13 : STD_LOGIC;
  SIGNAL and_dcpl_18 : STD_LOGIC;
  SIGNAL and_dcpl_23 : STD_LOGIC;
  SIGNAL and_dcpl_28 : STD_LOGIC;
  SIGNAL and_dcpl_29 : STD_LOGIC;
  SIGNAL and_dcpl_30 : STD_LOGIC;
  SIGNAL and_dcpl_31 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_35 : STD_LOGIC;
  SIGNAL and_dcpl_36 : STD_LOGIC;
  SIGNAL and_dcpl_38 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_56 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_62 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_77 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_87 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_90 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_104 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_114 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL and_dcpl_121 : STD_LOGIC;
  SIGNAL and_dcpl_126 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_137 : STD_LOGIC;
  SIGNAL and_dcpl_138 : STD_LOGIC;
  SIGNAL and_dcpl_139 : STD_LOGIC;
  SIGNAL and_dcpl_141 : STD_LOGIC;
  SIGNAL and_dcpl_143 : STD_LOGIC;
  SIGNAL and_dcpl_144 : STD_LOGIC;
  SIGNAL and_dcpl_146 : STD_LOGIC;
  SIGNAL and_dcpl_148 : STD_LOGIC;
  SIGNAL and_dcpl_153 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_163 : STD_LOGIC;
  SIGNAL and_dcpl_164 : STD_LOGIC;
  SIGNAL and_dcpl_165 : STD_LOGIC;
  SIGNAL and_dcpl_166 : STD_LOGIC;
  SIGNAL and_dcpl_168 : STD_LOGIC;
  SIGNAL and_dcpl_170 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_180 : STD_LOGIC;
  SIGNAL and_dcpl_185 : STD_LOGIC;
  SIGNAL and_dcpl_190 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL and_dcpl_193 : STD_LOGIC;
  SIGNAL and_dcpl_195 : STD_LOGIC;
  SIGNAL and_dcpl_197 : STD_LOGIC;
  SIGNAL and_dcpl_198 : STD_LOGIC;
  SIGNAL and_dcpl_200 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL and_dcpl_212 : STD_LOGIC;
  SIGNAL and_dcpl_217 : STD_LOGIC;
  SIGNAL and_dcpl_218 : STD_LOGIC;
  SIGNAL and_dcpl_219 : STD_LOGIC;
  SIGNAL and_dcpl_220 : STD_LOGIC;
  SIGNAL and_dcpl_222 : STD_LOGIC;
  SIGNAL and_dcpl_224 : STD_LOGIC;
  SIGNAL and_dcpl_225 : STD_LOGIC;
  SIGNAL and_dcpl_227 : STD_LOGIC;
  SIGNAL and_dcpl_229 : STD_LOGIC;
  SIGNAL and_dcpl_234 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_244 : STD_LOGIC;
  SIGNAL and_dcpl_245 : STD_LOGIC;
  SIGNAL and_dcpl_246 : STD_LOGIC;
  SIGNAL and_dcpl_247 : STD_LOGIC;
  SIGNAL and_dcpl_249 : STD_LOGIC;
  SIGNAL and_dcpl_251 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL and_dcpl_254 : STD_LOGIC;
  SIGNAL and_dcpl_256 : STD_LOGIC;
  SIGNAL and_dcpl_261 : STD_LOGIC;
  SIGNAL and_dcpl_266 : STD_LOGIC;
  SIGNAL and_dcpl_271 : STD_LOGIC;
  SIGNAL and_dcpl_272 : STD_LOGIC;
  SIGNAL and_dcpl_274 : STD_LOGIC;
  SIGNAL and_dcpl_276 : STD_LOGIC;
  SIGNAL and_dcpl_278 : STD_LOGIC;
  SIGNAL and_dcpl_280 : STD_LOGIC;
  SIGNAL and_dcpl_285 : STD_LOGIC;
  SIGNAL and_dcpl_291 : STD_LOGIC;
  SIGNAL and_dcpl_292 : STD_LOGIC;
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL and_dcpl_294 : STD_LOGIC;
  SIGNAL and_dcpl_295 : STD_LOGIC;
  SIGNAL and_dcpl_296 : STD_LOGIC;
  SIGNAL and_dcpl_298 : STD_LOGIC;
  SIGNAL not_tmp_54 : STD_LOGIC;
  SIGNAL or_tmp_2 : STD_LOGIC;
  SIGNAL and_dcpl_300 : STD_LOGIC;
  SIGNAL and_dcpl_301 : STD_LOGIC;
  SIGNAL and_dcpl_302 : STD_LOGIC;
  SIGNAL and_dcpl_304 : STD_LOGIC;
  SIGNAL and_tmp : STD_LOGIC;
  SIGNAL and_dcpl_306 : STD_LOGIC;
  SIGNAL and_dcpl_307 : STD_LOGIC;
  SIGNAL and_dcpl_308 : STD_LOGIC;
  SIGNAL and_dcpl_310 : STD_LOGIC;
  SIGNAL and_tmp_2 : STD_LOGIC;
  SIGNAL and_dcpl_312 : STD_LOGIC;
  SIGNAL and_dcpl_313 : STD_LOGIC;
  SIGNAL and_dcpl_314 : STD_LOGIC;
  SIGNAL and_dcpl_316 : STD_LOGIC;
  SIGNAL and_tmp_5 : STD_LOGIC;
  SIGNAL and_dcpl_318 : STD_LOGIC;
  SIGNAL and_tmp_9 : STD_LOGIC;
  SIGNAL and_dcpl_324 : STD_LOGIC;
  SIGNAL and_tmp_13 : STD_LOGIC;
  SIGNAL and_dcpl_330 : STD_LOGIC;
  SIGNAL mux_tmp_19 : STD_LOGIC;
  SIGNAL and_tmp_17 : STD_LOGIC;
  SIGNAL and_dcpl_336 : STD_LOGIC;
  SIGNAL mux_tmp_22 : STD_LOGIC;
  SIGNAL mux_tmp_23 : STD_LOGIC;
  SIGNAL and_tmp_21 : STD_LOGIC;
  SIGNAL and_dcpl_342 : STD_LOGIC;
  SIGNAL mux_tmp_26 : STD_LOGIC;
  SIGNAL mux_tmp_27 : STD_LOGIC;
  SIGNAL mux_tmp_28 : STD_LOGIC;
  SIGNAL and_tmp_25 : STD_LOGIC;
  SIGNAL and_dcpl_348 : STD_LOGIC;
  SIGNAL and_tmp_35 : STD_LOGIC;
  SIGNAL and_dcpl_355 : STD_LOGIC;
  SIGNAL and_dcpl_356 : STD_LOGIC;
  SIGNAL and_dcpl_358 : STD_LOGIC;
  SIGNAL or_tmp_80 : STD_LOGIC;
  SIGNAL and_dcpl_360 : STD_LOGIC;
  SIGNAL and_dcpl_362 : STD_LOGIC;
  SIGNAL mux_tmp_32 : STD_LOGIC;
  SIGNAL and_dcpl_364 : STD_LOGIC;
  SIGNAL and_dcpl_366 : STD_LOGIC;
  SIGNAL mux_tmp_34 : STD_LOGIC;
  SIGNAL mux_tmp_35 : STD_LOGIC;
  SIGNAL and_dcpl_368 : STD_LOGIC;
  SIGNAL and_dcpl_370 : STD_LOGIC;
  SIGNAL mux_tmp_37 : STD_LOGIC;
  SIGNAL mux_tmp_38 : STD_LOGIC;
  SIGNAL mux_tmp_39 : STD_LOGIC;
  SIGNAL and_dcpl_372 : STD_LOGIC;
  SIGNAL mux_tmp_41 : STD_LOGIC;
  SIGNAL mux_tmp_42 : STD_LOGIC;
  SIGNAL mux_tmp_43 : STD_LOGIC;
  SIGNAL mux_tmp_44 : STD_LOGIC;
  SIGNAL and_dcpl_376 : STD_LOGIC;
  SIGNAL mux_tmp_46 : STD_LOGIC;
  SIGNAL mux_tmp_47 : STD_LOGIC;
  SIGNAL mux_tmp_48 : STD_LOGIC;
  SIGNAL mux_tmp_49 : STD_LOGIC;
  SIGNAL mux_tmp_50 : STD_LOGIC;
  SIGNAL and_dcpl_379 : STD_LOGIC;
  SIGNAL mux_tmp_52 : STD_LOGIC;
  SIGNAL mux_tmp_53 : STD_LOGIC;
  SIGNAL mux_tmp_54 : STD_LOGIC;
  SIGNAL mux_tmp_55 : STD_LOGIC;
  SIGNAL mux_tmp_56 : STD_LOGIC;
  SIGNAL mux_tmp_57 : STD_LOGIC;
  SIGNAL and_dcpl_382 : STD_LOGIC;
  SIGNAL mux_tmp_59 : STD_LOGIC;
  SIGNAL mux_tmp_60 : STD_LOGIC;
  SIGNAL mux_tmp_61 : STD_LOGIC;
  SIGNAL mux_tmp_62 : STD_LOGIC;
  SIGNAL mux_tmp_63 : STD_LOGIC;
  SIGNAL mux_tmp_64 : STD_LOGIC;
  SIGNAL mux_tmp_65 : STD_LOGIC;
  SIGNAL and_dcpl_385 : STD_LOGIC;
  SIGNAL mux_tmp_67 : STD_LOGIC;
  SIGNAL mux_tmp_68 : STD_LOGIC;
  SIGNAL mux_tmp_69 : STD_LOGIC;
  SIGNAL mux_tmp_70 : STD_LOGIC;
  SIGNAL mux_tmp_71 : STD_LOGIC;
  SIGNAL mux_tmp_72 : STD_LOGIC;
  SIGNAL mux_tmp_73 : STD_LOGIC;
  SIGNAL mux_tmp_74 : STD_LOGIC;
  SIGNAL and_dcpl_388 : STD_LOGIC;
  SIGNAL and_tmp_44 : STD_LOGIC;
  SIGNAL mux_tmp_76 : STD_LOGIC;
  SIGNAL and_dcpl_393 : STD_LOGIC;
  SIGNAL and_dcpl_394 : STD_LOGIC;
  SIGNAL and_dcpl_395 : STD_LOGIC;
  SIGNAL or_tmp_185 : STD_LOGIC;
  SIGNAL and_dcpl_397 : STD_LOGIC;
  SIGNAL and_dcpl_398 : STD_LOGIC;
  SIGNAL and_tmp_45 : STD_LOGIC;
  SIGNAL and_dcpl_400 : STD_LOGIC;
  SIGNAL and_dcpl_401 : STD_LOGIC;
  SIGNAL and_tmp_47 : STD_LOGIC;
  SIGNAL and_dcpl_403 : STD_LOGIC;
  SIGNAL and_dcpl_404 : STD_LOGIC;
  SIGNAL and_tmp_50 : STD_LOGIC;
  SIGNAL and_dcpl_406 : STD_LOGIC;
  SIGNAL and_tmp_54 : STD_LOGIC;
  SIGNAL and_dcpl_409 : STD_LOGIC;
  SIGNAL and_tmp_58 : STD_LOGIC;
  SIGNAL and_dcpl_413 : STD_LOGIC;
  SIGNAL mux_tmp_84 : STD_LOGIC;
  SIGNAL and_tmp_62 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL mux_tmp_87 : STD_LOGIC;
  SIGNAL mux_tmp_88 : STD_LOGIC;
  SIGNAL and_tmp_66 : STD_LOGIC;
  SIGNAL and_dcpl_421 : STD_LOGIC;
  SIGNAL mux_tmp_91 : STD_LOGIC;
  SIGNAL mux_tmp_92 : STD_LOGIC;
  SIGNAL mux_tmp_93 : STD_LOGIC;
  SIGNAL and_tmp_70 : STD_LOGIC;
  SIGNAL and_dcpl_425 : STD_LOGIC;
  SIGNAL and_tmp_80 : STD_LOGIC;
  SIGNAL and_dcpl_430 : STD_LOGIC;
  SIGNAL and_dcpl_431 : STD_LOGIC;
  SIGNAL or_tmp_263 : STD_LOGIC;
  SIGNAL and_dcpl_433 : STD_LOGIC;
  SIGNAL mux_tmp_97 : STD_LOGIC;
  SIGNAL and_dcpl_435 : STD_LOGIC;
  SIGNAL mux_tmp_99 : STD_LOGIC;
  SIGNAL mux_tmp_100 : STD_LOGIC;
  SIGNAL and_dcpl_437 : STD_LOGIC;
  SIGNAL mux_tmp_102 : STD_LOGIC;
  SIGNAL mux_tmp_103 : STD_LOGIC;
  SIGNAL mux_tmp_104 : STD_LOGIC;
  SIGNAL and_dcpl_439 : STD_LOGIC;
  SIGNAL mux_tmp_106 : STD_LOGIC;
  SIGNAL mux_tmp_107 : STD_LOGIC;
  SIGNAL mux_tmp_108 : STD_LOGIC;
  SIGNAL mux_tmp_109 : STD_LOGIC;
  SIGNAL and_dcpl_442 : STD_LOGIC;
  SIGNAL mux_tmp_111 : STD_LOGIC;
  SIGNAL mux_tmp_112 : STD_LOGIC;
  SIGNAL mux_tmp_113 : STD_LOGIC;
  SIGNAL mux_tmp_114 : STD_LOGIC;
  SIGNAL mux_tmp_115 : STD_LOGIC;
  SIGNAL and_dcpl_445 : STD_LOGIC;
  SIGNAL mux_tmp_117 : STD_LOGIC;
  SIGNAL mux_tmp_118 : STD_LOGIC;
  SIGNAL mux_tmp_119 : STD_LOGIC;
  SIGNAL mux_tmp_120 : STD_LOGIC;
  SIGNAL mux_tmp_121 : STD_LOGIC;
  SIGNAL mux_tmp_122 : STD_LOGIC;
  SIGNAL and_dcpl_448 : STD_LOGIC;
  SIGNAL mux_tmp_124 : STD_LOGIC;
  SIGNAL mux_tmp_125 : STD_LOGIC;
  SIGNAL mux_tmp_126 : STD_LOGIC;
  SIGNAL mux_tmp_127 : STD_LOGIC;
  SIGNAL mux_tmp_128 : STD_LOGIC;
  SIGNAL mux_tmp_129 : STD_LOGIC;
  SIGNAL mux_tmp_130 : STD_LOGIC;
  SIGNAL and_dcpl_451 : STD_LOGIC;
  SIGNAL mux_tmp_132 : STD_LOGIC;
  SIGNAL mux_tmp_133 : STD_LOGIC;
  SIGNAL mux_tmp_134 : STD_LOGIC;
  SIGNAL mux_tmp_135 : STD_LOGIC;
  SIGNAL mux_tmp_136 : STD_LOGIC;
  SIGNAL mux_tmp_137 : STD_LOGIC;
  SIGNAL mux_tmp_138 : STD_LOGIC;
  SIGNAL mux_tmp_139 : STD_LOGIC;
  SIGNAL and_dcpl_454 : STD_LOGIC;
  SIGNAL and_tmp_89 : STD_LOGIC;
  SIGNAL mux_tmp_141 : STD_LOGIC;
  SIGNAL and_dcpl_460 : STD_LOGIC;
  SIGNAL and_dcpl_461 : STD_LOGIC;
  SIGNAL and_dcpl_462 : STD_LOGIC;
  SIGNAL and_dcpl_463 : STD_LOGIC;
  SIGNAL not_tmp_332 : STD_LOGIC;
  SIGNAL or_tmp_368 : STD_LOGIC;
  SIGNAL and_dcpl_465 : STD_LOGIC;
  SIGNAL and_dcpl_466 : STD_LOGIC;
  SIGNAL and_dcpl_467 : STD_LOGIC;
  SIGNAL and_tmp_90 : STD_LOGIC;
  SIGNAL and_dcpl_469 : STD_LOGIC;
  SIGNAL and_dcpl_470 : STD_LOGIC;
  SIGNAL and_dcpl_471 : STD_LOGIC;
  SIGNAL and_tmp_92 : STD_LOGIC;
  SIGNAL and_dcpl_473 : STD_LOGIC;
  SIGNAL and_dcpl_474 : STD_LOGIC;
  SIGNAL and_dcpl_475 : STD_LOGIC;
  SIGNAL and_tmp_95 : STD_LOGIC;
  SIGNAL and_dcpl_477 : STD_LOGIC;
  SIGNAL and_tmp_99 : STD_LOGIC;
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL and_tmp_103 : STD_LOGIC;
  SIGNAL and_dcpl_483 : STD_LOGIC;
  SIGNAL mux_tmp_149 : STD_LOGIC;
  SIGNAL and_tmp_107 : STD_LOGIC;
  SIGNAL and_dcpl_486 : STD_LOGIC;
  SIGNAL mux_tmp_152 : STD_LOGIC;
  SIGNAL mux_tmp_153 : STD_LOGIC;
  SIGNAL and_tmp_111 : STD_LOGIC;
  SIGNAL and_dcpl_489 : STD_LOGIC;
  SIGNAL mux_tmp_156 : STD_LOGIC;
  SIGNAL mux_tmp_157 : STD_LOGIC;
  SIGNAL mux_tmp_158 : STD_LOGIC;
  SIGNAL and_tmp_115 : STD_LOGIC;
  SIGNAL and_dcpl_492 : STD_LOGIC;
  SIGNAL and_tmp_125 : STD_LOGIC;
  SIGNAL and_dcpl_498 : STD_LOGIC;
  SIGNAL or_tmp_446 : STD_LOGIC;
  SIGNAL and_dcpl_500 : STD_LOGIC;
  SIGNAL mux_tmp_162 : STD_LOGIC;
  SIGNAL and_dcpl_502 : STD_LOGIC;
  SIGNAL mux_tmp_164 : STD_LOGIC;
  SIGNAL mux_tmp_165 : STD_LOGIC;
  SIGNAL and_dcpl_504 : STD_LOGIC;
  SIGNAL mux_tmp_167 : STD_LOGIC;
  SIGNAL mux_tmp_168 : STD_LOGIC;
  SIGNAL mux_tmp_169 : STD_LOGIC;
  SIGNAL and_dcpl_506 : STD_LOGIC;
  SIGNAL mux_tmp_171 : STD_LOGIC;
  SIGNAL mux_tmp_172 : STD_LOGIC;
  SIGNAL mux_tmp_173 : STD_LOGIC;
  SIGNAL mux_tmp_174 : STD_LOGIC;
  SIGNAL and_dcpl_508 : STD_LOGIC;
  SIGNAL mux_tmp_176 : STD_LOGIC;
  SIGNAL mux_tmp_177 : STD_LOGIC;
  SIGNAL mux_tmp_178 : STD_LOGIC;
  SIGNAL mux_tmp_179 : STD_LOGIC;
  SIGNAL mux_tmp_180 : STD_LOGIC;
  SIGNAL and_dcpl_510 : STD_LOGIC;
  SIGNAL mux_tmp_182 : STD_LOGIC;
  SIGNAL mux_tmp_183 : STD_LOGIC;
  SIGNAL mux_tmp_184 : STD_LOGIC;
  SIGNAL mux_tmp_185 : STD_LOGIC;
  SIGNAL mux_tmp_186 : STD_LOGIC;
  SIGNAL mux_tmp_187 : STD_LOGIC;
  SIGNAL and_dcpl_512 : STD_LOGIC;
  SIGNAL mux_tmp_189 : STD_LOGIC;
  SIGNAL mux_tmp_190 : STD_LOGIC;
  SIGNAL mux_tmp_191 : STD_LOGIC;
  SIGNAL mux_tmp_192 : STD_LOGIC;
  SIGNAL mux_tmp_193 : STD_LOGIC;
  SIGNAL mux_tmp_194 : STD_LOGIC;
  SIGNAL mux_tmp_195 : STD_LOGIC;
  SIGNAL and_dcpl_514 : STD_LOGIC;
  SIGNAL mux_tmp_197 : STD_LOGIC;
  SIGNAL mux_tmp_198 : STD_LOGIC;
  SIGNAL mux_tmp_199 : STD_LOGIC;
  SIGNAL mux_tmp_200 : STD_LOGIC;
  SIGNAL mux_tmp_201 : STD_LOGIC;
  SIGNAL mux_tmp_202 : STD_LOGIC;
  SIGNAL mux_tmp_203 : STD_LOGIC;
  SIGNAL mux_tmp_204 : STD_LOGIC;
  SIGNAL and_dcpl_516 : STD_LOGIC;
  SIGNAL and_tmp_134 : STD_LOGIC;
  SIGNAL mux_tmp_206 : STD_LOGIC;
  SIGNAL and_dcpl_520 : STD_LOGIC;
  SIGNAL and_dcpl_521 : STD_LOGIC;
  SIGNAL or_tmp_551 : STD_LOGIC;
  SIGNAL and_dcpl_523 : STD_LOGIC;
  SIGNAL and_dcpl_524 : STD_LOGIC;
  SIGNAL and_tmp_135 : STD_LOGIC;
  SIGNAL and_dcpl_526 : STD_LOGIC;
  SIGNAL and_dcpl_527 : STD_LOGIC;
  SIGNAL and_tmp_137 : STD_LOGIC;
  SIGNAL and_dcpl_529 : STD_LOGIC;
  SIGNAL and_dcpl_530 : STD_LOGIC;
  SIGNAL and_tmp_140 : STD_LOGIC;
  SIGNAL and_dcpl_532 : STD_LOGIC;
  SIGNAL and_tmp_144 : STD_LOGIC;
  SIGNAL and_dcpl_534 : STD_LOGIC;
  SIGNAL and_tmp_148 : STD_LOGIC;
  SIGNAL and_dcpl_536 : STD_LOGIC;
  SIGNAL mux_tmp_214 : STD_LOGIC;
  SIGNAL and_tmp_152 : STD_LOGIC;
  SIGNAL and_dcpl_538 : STD_LOGIC;
  SIGNAL mux_tmp_217 : STD_LOGIC;
  SIGNAL mux_tmp_218 : STD_LOGIC;
  SIGNAL and_tmp_156 : STD_LOGIC;
  SIGNAL and_dcpl_540 : STD_LOGIC;
  SIGNAL mux_tmp_221 : STD_LOGIC;
  SIGNAL mux_tmp_222 : STD_LOGIC;
  SIGNAL mux_tmp_223 : STD_LOGIC;
  SIGNAL and_tmp_160 : STD_LOGIC;
  SIGNAL and_dcpl_542 : STD_LOGIC;
  SIGNAL and_tmp_170 : STD_LOGIC;
  SIGNAL and_dcpl_546 : STD_LOGIC;
  SIGNAL or_tmp_629 : STD_LOGIC;
  SIGNAL and_dcpl_548 : STD_LOGIC;
  SIGNAL mux_tmp_227 : STD_LOGIC;
  SIGNAL and_dcpl_550 : STD_LOGIC;
  SIGNAL mux_tmp_229 : STD_LOGIC;
  SIGNAL mux_tmp_230 : STD_LOGIC;
  SIGNAL and_dcpl_552 : STD_LOGIC;
  SIGNAL mux_tmp_232 : STD_LOGIC;
  SIGNAL mux_tmp_233 : STD_LOGIC;
  SIGNAL mux_tmp_234 : STD_LOGIC;
  SIGNAL and_dcpl_554 : STD_LOGIC;
  SIGNAL mux_tmp_236 : STD_LOGIC;
  SIGNAL mux_tmp_237 : STD_LOGIC;
  SIGNAL mux_tmp_238 : STD_LOGIC;
  SIGNAL mux_tmp_239 : STD_LOGIC;
  SIGNAL and_dcpl_556 : STD_LOGIC;
  SIGNAL mux_tmp_241 : STD_LOGIC;
  SIGNAL mux_tmp_242 : STD_LOGIC;
  SIGNAL mux_tmp_243 : STD_LOGIC;
  SIGNAL mux_tmp_244 : STD_LOGIC;
  SIGNAL mux_tmp_245 : STD_LOGIC;
  SIGNAL and_dcpl_558 : STD_LOGIC;
  SIGNAL mux_tmp_247 : STD_LOGIC;
  SIGNAL mux_tmp_248 : STD_LOGIC;
  SIGNAL mux_tmp_249 : STD_LOGIC;
  SIGNAL mux_tmp_250 : STD_LOGIC;
  SIGNAL mux_tmp_251 : STD_LOGIC;
  SIGNAL mux_tmp_252 : STD_LOGIC;
  SIGNAL and_dcpl_560 : STD_LOGIC;
  SIGNAL mux_tmp_254 : STD_LOGIC;
  SIGNAL mux_tmp_255 : STD_LOGIC;
  SIGNAL mux_tmp_256 : STD_LOGIC;
  SIGNAL mux_tmp_257 : STD_LOGIC;
  SIGNAL mux_tmp_258 : STD_LOGIC;
  SIGNAL mux_tmp_259 : STD_LOGIC;
  SIGNAL mux_tmp_260 : STD_LOGIC;
  SIGNAL and_dcpl_562 : STD_LOGIC;
  SIGNAL mux_tmp_262 : STD_LOGIC;
  SIGNAL mux_tmp_263 : STD_LOGIC;
  SIGNAL mux_tmp_264 : STD_LOGIC;
  SIGNAL mux_tmp_265 : STD_LOGIC;
  SIGNAL mux_tmp_266 : STD_LOGIC;
  SIGNAL mux_tmp_267 : STD_LOGIC;
  SIGNAL mux_tmp_268 : STD_LOGIC;
  SIGNAL mux_tmp_269 : STD_LOGIC;
  SIGNAL and_dcpl_564 : STD_LOGIC;
  SIGNAL and_tmp_179 : STD_LOGIC;
  SIGNAL mux_tmp_271 : STD_LOGIC;
  SIGNAL and_dcpl_568 : STD_LOGIC;
  SIGNAL and_dcpl_569 : STD_LOGIC;
  SIGNAL and_dcpl_570 : STD_LOGIC;
  SIGNAL and_dcpl_571 : STD_LOGIC;
  SIGNAL or_tmp_733 : STD_LOGIC;
  SIGNAL and_dcpl_573 : STD_LOGIC;
  SIGNAL and_dcpl_574 : STD_LOGIC;
  SIGNAL and_dcpl_575 : STD_LOGIC;
  SIGNAL and_tmp_180 : STD_LOGIC;
  SIGNAL and_dcpl_577 : STD_LOGIC;
  SIGNAL and_dcpl_578 : STD_LOGIC;
  SIGNAL and_dcpl_579 : STD_LOGIC;
  SIGNAL and_tmp_182 : STD_LOGIC;
  SIGNAL and_dcpl_581 : STD_LOGIC;
  SIGNAL and_dcpl_582 : STD_LOGIC;
  SIGNAL and_dcpl_583 : STD_LOGIC;
  SIGNAL and_tmp_185 : STD_LOGIC;
  SIGNAL and_dcpl_585 : STD_LOGIC;
  SIGNAL and_tmp_189 : STD_LOGIC;
  SIGNAL and_dcpl_589 : STD_LOGIC;
  SIGNAL and_tmp_193 : STD_LOGIC;
  SIGNAL and_dcpl_593 : STD_LOGIC;
  SIGNAL mux_tmp_279 : STD_LOGIC;
  SIGNAL and_tmp_197 : STD_LOGIC;
  SIGNAL and_dcpl_597 : STD_LOGIC;
  SIGNAL mux_tmp_282 : STD_LOGIC;
  SIGNAL mux_tmp_283 : STD_LOGIC;
  SIGNAL and_tmp_201 : STD_LOGIC;
  SIGNAL and_dcpl_601 : STD_LOGIC;
  SIGNAL mux_tmp_286 : STD_LOGIC;
  SIGNAL mux_tmp_287 : STD_LOGIC;
  SIGNAL mux_tmp_288 : STD_LOGIC;
  SIGNAL and_tmp_205 : STD_LOGIC;
  SIGNAL and_dcpl_605 : STD_LOGIC;
  SIGNAL or_tmp_808 : STD_LOGIC;
  SIGNAL mux_tmp_291 : STD_LOGIC;
  SIGNAL mux_tmp_292 : STD_LOGIC;
  SIGNAL mux_tmp_293 : STD_LOGIC;
  SIGNAL mux_tmp_294 : STD_LOGIC;
  SIGNAL mux_tmp_295 : STD_LOGIC;
  SIGNAL mux_tmp_296 : STD_LOGIC;
  SIGNAL mux_tmp_297 : STD_LOGIC;
  SIGNAL mux_tmp_298 : STD_LOGIC;
  SIGNAL and_tmp_206 : STD_LOGIC;
  SIGNAL and_dcpl_610 : STD_LOGIC;
  SIGNAL or_tmp_820 : STD_LOGIC;
  SIGNAL and_dcpl_612 : STD_LOGIC;
  SIGNAL mux_tmp_301 : STD_LOGIC;
  SIGNAL and_dcpl_614 : STD_LOGIC;
  SIGNAL mux_tmp_303 : STD_LOGIC;
  SIGNAL mux_tmp_304 : STD_LOGIC;
  SIGNAL and_dcpl_616 : STD_LOGIC;
  SIGNAL mux_tmp_306 : STD_LOGIC;
  SIGNAL mux_tmp_307 : STD_LOGIC;
  SIGNAL mux_tmp_308 : STD_LOGIC;
  SIGNAL and_dcpl_618 : STD_LOGIC;
  SIGNAL mux_tmp_310 : STD_LOGIC;
  SIGNAL mux_tmp_311 : STD_LOGIC;
  SIGNAL mux_tmp_312 : STD_LOGIC;
  SIGNAL mux_tmp_313 : STD_LOGIC;
  SIGNAL and_dcpl_622 : STD_LOGIC;
  SIGNAL mux_tmp_315 : STD_LOGIC;
  SIGNAL mux_tmp_316 : STD_LOGIC;
  SIGNAL mux_tmp_317 : STD_LOGIC;
  SIGNAL mux_tmp_318 : STD_LOGIC;
  SIGNAL mux_tmp_319 : STD_LOGIC;
  SIGNAL and_dcpl_625 : STD_LOGIC;
  SIGNAL mux_tmp_321 : STD_LOGIC;
  SIGNAL mux_tmp_322 : STD_LOGIC;
  SIGNAL mux_tmp_323 : STD_LOGIC;
  SIGNAL mux_tmp_324 : STD_LOGIC;
  SIGNAL mux_tmp_325 : STD_LOGIC;
  SIGNAL mux_tmp_326 : STD_LOGIC;
  SIGNAL and_dcpl_628 : STD_LOGIC;
  SIGNAL mux_tmp_328 : STD_LOGIC;
  SIGNAL mux_tmp_329 : STD_LOGIC;
  SIGNAL mux_tmp_330 : STD_LOGIC;
  SIGNAL mux_tmp_331 : STD_LOGIC;
  SIGNAL mux_tmp_332 : STD_LOGIC;
  SIGNAL mux_tmp_333 : STD_LOGIC;
  SIGNAL mux_tmp_334 : STD_LOGIC;
  SIGNAL and_dcpl_631 : STD_LOGIC;
  SIGNAL mux_tmp_336 : STD_LOGIC;
  SIGNAL mux_tmp_337 : STD_LOGIC;
  SIGNAL mux_tmp_338 : STD_LOGIC;
  SIGNAL mux_tmp_339 : STD_LOGIC;
  SIGNAL mux_tmp_340 : STD_LOGIC;
  SIGNAL mux_tmp_341 : STD_LOGIC;
  SIGNAL mux_tmp_342 : STD_LOGIC;
  SIGNAL mux_tmp_343 : STD_LOGIC;
  SIGNAL and_dcpl_634 : STD_LOGIC;
  SIGNAL or_tmp_921 : STD_LOGIC;
  SIGNAL mux_tmp_345 : STD_LOGIC;
  SIGNAL mux_tmp_346 : STD_LOGIC;
  SIGNAL mux_tmp_347 : STD_LOGIC;
  SIGNAL mux_tmp_348 : STD_LOGIC;
  SIGNAL mux_tmp_349 : STD_LOGIC;
  SIGNAL mux_tmp_350 : STD_LOGIC;
  SIGNAL mux_tmp_351 : STD_LOGIC;
  SIGNAL mux_tmp_352 : STD_LOGIC;
  SIGNAL mux_tmp_353 : STD_LOGIC;
  SIGNAL mux_tmp_354 : STD_LOGIC;
  SIGNAL and_dcpl_638 : STD_LOGIC;
  SIGNAL and_dcpl_639 : STD_LOGIC;
  SIGNAL or_tmp_934 : STD_LOGIC;
  SIGNAL and_dcpl_641 : STD_LOGIC;
  SIGNAL and_dcpl_642 : STD_LOGIC;
  SIGNAL and_tmp_207 : STD_LOGIC;
  SIGNAL and_dcpl_644 : STD_LOGIC;
  SIGNAL and_dcpl_645 : STD_LOGIC;
  SIGNAL and_tmp_209 : STD_LOGIC;
  SIGNAL and_dcpl_647 : STD_LOGIC;
  SIGNAL and_dcpl_648 : STD_LOGIC;
  SIGNAL and_tmp_212 : STD_LOGIC;
  SIGNAL and_dcpl_650 : STD_LOGIC;
  SIGNAL and_tmp_216 : STD_LOGIC;
  SIGNAL and_dcpl_653 : STD_LOGIC;
  SIGNAL and_tmp_220 : STD_LOGIC;
  SIGNAL and_dcpl_657 : STD_LOGIC;
  SIGNAL mux_tmp_362 : STD_LOGIC;
  SIGNAL and_tmp_224 : STD_LOGIC;
  SIGNAL and_dcpl_661 : STD_LOGIC;
  SIGNAL mux_tmp_365 : STD_LOGIC;
  SIGNAL mux_tmp_366 : STD_LOGIC;
  SIGNAL and_tmp_228 : STD_LOGIC;
  SIGNAL and_dcpl_665 : STD_LOGIC;
  SIGNAL mux_tmp_369 : STD_LOGIC;
  SIGNAL mux_tmp_370 : STD_LOGIC;
  SIGNAL mux_tmp_371 : STD_LOGIC;
  SIGNAL and_tmp_232 : STD_LOGIC;
  SIGNAL and_dcpl_669 : STD_LOGIC;
  SIGNAL or_tmp_1009 : STD_LOGIC;
  SIGNAL mux_tmp_374 : STD_LOGIC;
  SIGNAL mux_tmp_375 : STD_LOGIC;
  SIGNAL mux_tmp_376 : STD_LOGIC;
  SIGNAL mux_tmp_377 : STD_LOGIC;
  SIGNAL mux_tmp_378 : STD_LOGIC;
  SIGNAL mux_tmp_379 : STD_LOGIC;
  SIGNAL mux_tmp_380 : STD_LOGIC;
  SIGNAL mux_tmp_381 : STD_LOGIC;
  SIGNAL and_tmp_233 : STD_LOGIC;
  SIGNAL and_dcpl_673 : STD_LOGIC;
  SIGNAL or_tmp_1021 : STD_LOGIC;
  SIGNAL and_dcpl_675 : STD_LOGIC;
  SIGNAL mux_tmp_384 : STD_LOGIC;
  SIGNAL and_dcpl_677 : STD_LOGIC;
  SIGNAL mux_tmp_386 : STD_LOGIC;
  SIGNAL mux_tmp_387 : STD_LOGIC;
  SIGNAL and_dcpl_679 : STD_LOGIC;
  SIGNAL mux_tmp_389 : STD_LOGIC;
  SIGNAL mux_tmp_390 : STD_LOGIC;
  SIGNAL mux_tmp_391 : STD_LOGIC;
  SIGNAL and_dcpl_681 : STD_LOGIC;
  SIGNAL mux_tmp_393 : STD_LOGIC;
  SIGNAL mux_tmp_394 : STD_LOGIC;
  SIGNAL mux_tmp_395 : STD_LOGIC;
  SIGNAL mux_tmp_396 : STD_LOGIC;
  SIGNAL and_dcpl_684 : STD_LOGIC;
  SIGNAL mux_tmp_398 : STD_LOGIC;
  SIGNAL mux_tmp_399 : STD_LOGIC;
  SIGNAL mux_tmp_400 : STD_LOGIC;
  SIGNAL mux_tmp_401 : STD_LOGIC;
  SIGNAL mux_tmp_402 : STD_LOGIC;
  SIGNAL and_dcpl_687 : STD_LOGIC;
  SIGNAL mux_tmp_404 : STD_LOGIC;
  SIGNAL mux_tmp_405 : STD_LOGIC;
  SIGNAL mux_tmp_406 : STD_LOGIC;
  SIGNAL mux_tmp_407 : STD_LOGIC;
  SIGNAL mux_tmp_408 : STD_LOGIC;
  SIGNAL mux_tmp_409 : STD_LOGIC;
  SIGNAL and_dcpl_690 : STD_LOGIC;
  SIGNAL mux_tmp_411 : STD_LOGIC;
  SIGNAL mux_tmp_412 : STD_LOGIC;
  SIGNAL mux_tmp_413 : STD_LOGIC;
  SIGNAL mux_tmp_414 : STD_LOGIC;
  SIGNAL mux_tmp_415 : STD_LOGIC;
  SIGNAL mux_tmp_416 : STD_LOGIC;
  SIGNAL mux_tmp_417 : STD_LOGIC;
  SIGNAL and_dcpl_693 : STD_LOGIC;
  SIGNAL mux_tmp_419 : STD_LOGIC;
  SIGNAL mux_tmp_420 : STD_LOGIC;
  SIGNAL mux_tmp_421 : STD_LOGIC;
  SIGNAL mux_tmp_422 : STD_LOGIC;
  SIGNAL mux_tmp_423 : STD_LOGIC;
  SIGNAL mux_tmp_424 : STD_LOGIC;
  SIGNAL mux_tmp_425 : STD_LOGIC;
  SIGNAL mux_tmp_426 : STD_LOGIC;
  SIGNAL and_dcpl_696 : STD_LOGIC;
  SIGNAL or_tmp_1122 : STD_LOGIC;
  SIGNAL mux_tmp_428 : STD_LOGIC;
  SIGNAL mux_tmp_429 : STD_LOGIC;
  SIGNAL mux_tmp_430 : STD_LOGIC;
  SIGNAL mux_tmp_431 : STD_LOGIC;
  SIGNAL mux_tmp_432 : STD_LOGIC;
  SIGNAL mux_tmp_433 : STD_LOGIC;
  SIGNAL mux_tmp_434 : STD_LOGIC;
  SIGNAL mux_tmp_435 : STD_LOGIC;
  SIGNAL mux_tmp_436 : STD_LOGIC;
  SIGNAL mux_tmp_437 : STD_LOGIC;
  SIGNAL rem_12cyc_st_10_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_10_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_9_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_9_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_8_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_8_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_7_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_7_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_6_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_6_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_5_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_5_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_4_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_4_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_3_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_3_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_2_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_2_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_12_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL result_sva_duc : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12cyc_st_12_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL asn_itm_12 : STD_LOGIC;
  SIGNAL main_stage_0_13 : STD_LOGIC;
  SIGNAL main_stage_0_3 : STD_LOGIC;
  SIGNAL asn_itm_1 : STD_LOGIC;
  SIGNAL main_stage_0_2 : STD_LOGIC;
  SIGNAL main_stage_0_4 : STD_LOGIC;
  SIGNAL asn_itm_2 : STD_LOGIC;
  SIGNAL main_stage_0_5 : STD_LOGIC;
  SIGNAL asn_itm_3 : STD_LOGIC;
  SIGNAL main_stage_0_6 : STD_LOGIC;
  SIGNAL asn_itm_4 : STD_LOGIC;
  SIGNAL asn_itm_5 : STD_LOGIC;
  SIGNAL main_stage_0_8 : STD_LOGIC;
  SIGNAL asn_itm_7 : STD_LOGIC;
  SIGNAL main_stage_0_9 : STD_LOGIC;
  SIGNAL asn_itm_8 : STD_LOGIC;
  SIGNAL main_stage_0_10 : STD_LOGIC;
  SIGNAL asn_itm_9 : STD_LOGIC;
  SIGNAL main_stage_0_7 : STD_LOGIC;
  SIGNAL asn_itm_6 : STD_LOGIC;
  SIGNAL main_stage_0_11 : STD_LOGIC;
  SIGNAL asn_itm_10 : STD_LOGIC;
  SIGNAL and_1173_cse : STD_LOGIC;
  SIGNAL and_1175_cse : STD_LOGIC;
  SIGNAL and_1177_cse : STD_LOGIC;
  SIGNAL and_1179_cse : STD_LOGIC;
  SIGNAL and_1181_cse : STD_LOGIC;
  SIGNAL and_1183_cse : STD_LOGIC;
  SIGNAL and_1185_cse : STD_LOGIC;
  SIGNAL and_1187_cse : STD_LOGIC;
  SIGNAL and_1189_cse : STD_LOGIC;
  SIGNAL and_1191_cse : STD_LOGIC;
  SIGNAL and_1193_cse : STD_LOGIC;
  SIGNAL and_1195_cse : STD_LOGIC;
  SIGNAL and_1197_cse : STD_LOGIC;
  SIGNAL or_1_cse : STD_LOGIC;
  SIGNAL or_6_cse : STD_LOGIC;
  SIGNAL or_10_cse : STD_LOGIC;
  SIGNAL or_15_cse : STD_LOGIC;
  SIGNAL or_21_cse : STD_LOGIC;
  SIGNAL or_28_cse : STD_LOGIC;
  SIGNAL or_37_cse : STD_LOGIC;
  SIGNAL or_48_cse : STD_LOGIC;
  SIGNAL or_83_cse : STD_LOGIC;
  SIGNAL nand_276_cse : STD_LOGIC;
  SIGNAL or_88_cse : STD_LOGIC;
  SIGNAL nand_274_cse : STD_LOGIC;
  SIGNAL or_93_cse : STD_LOGIC;
  SIGNAL nand_271_cse : STD_LOGIC;
  SIGNAL or_100_cse : STD_LOGIC;
  SIGNAL nand_267_cse : STD_LOGIC;
  SIGNAL or_109_cse : STD_LOGIC;
  SIGNAL or_120_cse : STD_LOGIC;
  SIGNAL or_133_cse : STD_LOGIC;
  SIGNAL or_148_cse : STD_LOGIC;
  SIGNAL or_190_cse : STD_LOGIC;
  SIGNAL or_195_cse : STD_LOGIC;
  SIGNAL or_199_cse : STD_LOGIC;
  SIGNAL or_204_cse : STD_LOGIC;
  SIGNAL or_210_cse : STD_LOGIC;
  SIGNAL or_217_cse : STD_LOGIC;
  SIGNAL or_226_cse : STD_LOGIC;
  SIGNAL or_237_cse : STD_LOGIC;
  SIGNAL or_270_cse : STD_LOGIC;
  SIGNAL or_275_cse : STD_LOGIC;
  SIGNAL or_280_cse : STD_LOGIC;
  SIGNAL or_287_cse : STD_LOGIC;
  SIGNAL or_296_cse : STD_LOGIC;
  SIGNAL or_307_cse : STD_LOGIC;
  SIGNAL or_320_cse : STD_LOGIC;
  SIGNAL or_335_cse : STD_LOGIC;
  SIGNAL nand_281_cse : STD_LOGIC;
  SIGNAL or_377_cse : STD_LOGIC;
  SIGNAL or_382_cse : STD_LOGIC;
  SIGNAL or_386_cse : STD_LOGIC;
  SIGNAL or_391_cse : STD_LOGIC;
  SIGNAL or_397_cse : STD_LOGIC;
  SIGNAL nand_215_cse : STD_LOGIC;
  SIGNAL or_404_cse : STD_LOGIC;
  SIGNAL nand_212_cse : STD_LOGIC;
  SIGNAL or_413_cse : STD_LOGIC;
  SIGNAL nand_208_cse : STD_LOGIC;
  SIGNAL or_424_cse : STD_LOGIC;
  SIGNAL or_458_cse : STD_LOGIC;
  SIGNAL or_463_cse : STD_LOGIC;
  SIGNAL nand_198_cse : STD_LOGIC;
  SIGNAL or_468_cse : STD_LOGIC;
  SIGNAL or_475_cse : STD_LOGIC;
  SIGNAL nand_189_cse : STD_LOGIC;
  SIGNAL or_484_cse : STD_LOGIC;
  SIGNAL or_495_cse : STD_LOGIC;
  SIGNAL or_508_cse : STD_LOGIC;
  SIGNAL nand_203_cse : STD_LOGIC;
  SIGNAL or_523_cse : STD_LOGIC;
  SIGNAL nand_250_cse : STD_LOGIC;
  SIGNAL or_564_cse : STD_LOGIC;
  SIGNAL or_569_cse : STD_LOGIC;
  SIGNAL or_573_cse : STD_LOGIC;
  SIGNAL or_578_cse : STD_LOGIC;
  SIGNAL or_584_cse : STD_LOGIC;
  SIGNAL or_591_cse : STD_LOGIC;
  SIGNAL or_600_cse : STD_LOGIC;
  SIGNAL or_611_cse : STD_LOGIC;
  SIGNAL or_643_cse : STD_LOGIC;
  SIGNAL or_648_cse : STD_LOGIC;
  SIGNAL or_653_cse : STD_LOGIC;
  SIGNAL or_660_cse : STD_LOGIC;
  SIGNAL or_669_cse : STD_LOGIC;
  SIGNAL or_680_cse : STD_LOGIC;
  SIGNAL or_693_cse : STD_LOGIC;
  SIGNAL or_708_cse : STD_LOGIC;
  SIGNAL or_748_cse : STD_LOGIC;
  SIGNAL or_753_cse : STD_LOGIC;
  SIGNAL or_757_cse : STD_LOGIC;
  SIGNAL or_762_cse : STD_LOGIC;
  SIGNAL or_768_cse : STD_LOGIC;
  SIGNAL or_775_cse : STD_LOGIC;
  SIGNAL or_784_cse : STD_LOGIC;
  SIGNAL or_795_cse : STD_LOGIC;
  SIGNAL or_837_cse : STD_LOGIC;
  SIGNAL nand_84_cse : STD_LOGIC;
  SIGNAL or_842_cse : STD_LOGIC;
  SIGNAL or_847_cse : STD_LOGIC;
  SIGNAL nand_79_cse : STD_LOGIC;
  SIGNAL or_854_cse : STD_LOGIC;
  SIGNAL or_863_cse : STD_LOGIC;
  SIGNAL or_874_cse : STD_LOGIC;
  SIGNAL or_887_cse : STD_LOGIC;
  SIGNAL or_902_cse : STD_LOGIC;
  SIGNAL or_952_cse : STD_LOGIC;
  SIGNAL or_957_cse : STD_LOGIC;
  SIGNAL or_961_cse : STD_LOGIC;
  SIGNAL or_966_cse : STD_LOGIC;
  SIGNAL or_972_cse : STD_LOGIC;
  SIGNAL or_979_cse : STD_LOGIC;
  SIGNAL or_988_cse : STD_LOGIC;
  SIGNAL or_999_cse : STD_LOGIC;
  SIGNAL nand_57_cse : STD_LOGIC;
  SIGNAL or_1045_cse : STD_LOGIC;
  SIGNAL or_1050_cse : STD_LOGIC;
  SIGNAL or_1057_cse : STD_LOGIC;
  SIGNAL or_1066_cse : STD_LOGIC;
  SIGNAL nand_36_cse : STD_LOGIC;
  SIGNAL nand_29_cse : STD_LOGIC;
  SIGNAL nand_21_cse : STD_LOGIC;
  SIGNAL nand_222_cse : STD_LOGIC;
  SIGNAL nand_223_cse : STD_LOGIC;
  SIGNAL main_stage_0_12 : STD_LOGIC;
  SIGNAL m_buf_sva_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_2 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_3 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_4 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_5 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_6 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_7 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_8 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_9 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_10 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_11 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_buf_sva_12 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL asn_itm_11 : STD_LOGIC;
  SIGNAL mut_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_1_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_2_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_3_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_4_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_5_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_6_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_7_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_8_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_9_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_10_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_11_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_12_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_13_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_14_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_15_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_16_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_17_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_18_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_19_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_20_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_21_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_22_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_2_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_3_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_4_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_5_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_6_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_7_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_8_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_9_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_10_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mut_23_11_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL rem_12cyc_st_11_3_2 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL rem_12cyc_st_11_1_0 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL result_sva_duc_mx0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_1203_cse : STD_LOGIC;
  SIGNAL and_1205_cse : STD_LOGIC;
  SIGNAL and_1207_cse : STD_LOGIC;
  SIGNAL and_1209_cse : STD_LOGIC;
  SIGNAL and_1211_cse : STD_LOGIC;
  SIGNAL and_1213_cse : STD_LOGIC;
  SIGNAL and_1215_cse : STD_LOGIC;
  SIGNAL and_1217_cse : STD_LOGIC;
  SIGNAL and_1219_cse : STD_LOGIC;
  SIGNAL and_1221_cse : STD_LOGIC;
  SIGNAL and_1223_cse : STD_LOGIC;
  SIGNAL and_1225_cse : STD_LOGIC;
  SIGNAL and_1227_cse : STD_LOGIC;
  SIGNAL and_1229_cse : STD_LOGIC;
  SIGNAL and_1231_cse : STD_LOGIC;
  SIGNAL and_1233_cse : STD_LOGIC;
  SIGNAL and_1235_cse : STD_LOGIC;
  SIGNAL and_1237_cse : STD_LOGIC;
  SIGNAL and_1239_cse : STD_LOGIC;
  SIGNAL and_1241_cse : STD_LOGIC;
  SIGNAL and_1243_cse : STD_LOGIC;
  SIGNAL and_1245_cse : STD_LOGIC;
  SIGNAL and_1247_cse : STD_LOGIC;
  SIGNAL and_1249_cse : STD_LOGIC;
  SIGNAL and_1251_cse : STD_LOGIC;
  SIGNAL and_1253_cse : STD_LOGIC;
  SIGNAL and_1255_cse : STD_LOGIC;
  SIGNAL and_1257_cse : STD_LOGIC;
  SIGNAL and_1259_cse : STD_LOGIC;
  SIGNAL and_1261_cse : STD_LOGIC;
  SIGNAL and_1263_cse : STD_LOGIC;
  SIGNAL and_1265_cse : STD_LOGIC;
  SIGNAL and_1267_cse : STD_LOGIC;
  SIGNAL and_1269_cse : STD_LOGIC;
  SIGNAL and_1271_cse : STD_LOGIC;
  SIGNAL and_1273_cse : STD_LOGIC;
  SIGNAL and_1275_cse : STD_LOGIC;
  SIGNAL and_1277_cse : STD_LOGIC;
  SIGNAL and_1279_cse : STD_LOGIC;
  SIGNAL and_1281_cse : STD_LOGIC;
  SIGNAL and_1283_cse : STD_LOGIC;
  SIGNAL and_1285_cse : STD_LOGIC;
  SIGNAL and_1287_cse : STD_LOGIC;
  SIGNAL and_1289_cse : STD_LOGIC;
  SIGNAL and_1291_cse : STD_LOGIC;
  SIGNAL and_1293_cse : STD_LOGIC;
  SIGNAL and_1295_cse : STD_LOGIC;
  SIGNAL and_1297_cse : STD_LOGIC;
  SIGNAL and_1299_cse : STD_LOGIC;
  SIGNAL and_1301_cse : STD_LOGIC;
  SIGNAL and_1303_cse : STD_LOGIC;
  SIGNAL and_1305_cse : STD_LOGIC;
  SIGNAL and_1307_cse : STD_LOGIC;
  SIGNAL and_1309_cse : STD_LOGIC;
  SIGNAL and_1311_cse : STD_LOGIC;
  SIGNAL and_1313_cse : STD_LOGIC;
  SIGNAL and_1315_cse : STD_LOGIC;
  SIGNAL and_1317_cse : STD_LOGIC;
  SIGNAL and_1319_cse : STD_LOGIC;
  SIGNAL and_1321_cse : STD_LOGIC;
  SIGNAL and_1323_cse : STD_LOGIC;
  SIGNAL and_1325_cse : STD_LOGIC;
  SIGNAL and_1327_cse : STD_LOGIC;
  SIGNAL and_1329_cse : STD_LOGIC;
  SIGNAL and_1331_cse : STD_LOGIC;
  SIGNAL and_1333_cse : STD_LOGIC;
  SIGNAL and_1335_cse : STD_LOGIC;
  SIGNAL and_1337_cse : STD_LOGIC;
  SIGNAL and_1339_cse : STD_LOGIC;
  SIGNAL and_1341_cse : STD_LOGIC;
  SIGNAL and_1343_cse : STD_LOGIC;
  SIGNAL and_1345_cse : STD_LOGIC;
  SIGNAL and_1347_cse : STD_LOGIC;
  SIGNAL and_1349_cse : STD_LOGIC;
  SIGNAL and_1351_cse : STD_LOGIC;
  SIGNAL and_1353_cse : STD_LOGIC;
  SIGNAL and_1355_cse : STD_LOGIC;
  SIGNAL and_1357_cse : STD_LOGIC;
  SIGNAL and_1359_cse : STD_LOGIC;
  SIGNAL and_1361_cse : STD_LOGIC;
  SIGNAL and_1363_cse : STD_LOGIC;
  SIGNAL and_1365_cse : STD_LOGIC;
  SIGNAL and_1367_cse : STD_LOGIC;
  SIGNAL and_1369_cse : STD_LOGIC;
  SIGNAL and_1371_cse : STD_LOGIC;
  SIGNAL and_1373_cse : STD_LOGIC;
  SIGNAL and_1375_cse : STD_LOGIC;
  SIGNAL and_1377_cse : STD_LOGIC;
  SIGNAL and_1379_cse : STD_LOGIC;
  SIGNAL and_1381_cse : STD_LOGIC;
  SIGNAL and_1383_cse : STD_LOGIC;
  SIGNAL and_1385_cse : STD_LOGIC;
  SIGNAL and_1387_cse : STD_LOGIC;
  SIGNAL and_1389_cse : STD_LOGIC;
  SIGNAL and_1391_cse : STD_LOGIC;
  SIGNAL and_1393_cse : STD_LOGIC;
  SIGNAL and_1395_cse : STD_LOGIC;
  SIGNAL and_1397_cse : STD_LOGIC;
  SIGNAL and_1399_cse : STD_LOGIC;
  SIGNAL and_1401_cse : STD_LOGIC;
  SIGNAL and_1403_cse : STD_LOGIC;
  SIGNAL and_1405_cse : STD_LOGIC;
  SIGNAL and_1407_cse : STD_LOGIC;
  SIGNAL and_1409_cse : STD_LOGIC;
  SIGNAL and_1411_cse : STD_LOGIC;
  SIGNAL and_1413_cse : STD_LOGIC;
  SIGNAL and_1415_cse : STD_LOGIC;
  SIGNAL and_1417_cse : STD_LOGIC;
  SIGNAL and_1419_cse : STD_LOGIC;
  SIGNAL and_1421_cse : STD_LOGIC;
  SIGNAL and_1423_cse : STD_LOGIC;
  SIGNAL and_1425_cse : STD_LOGIC;
  SIGNAL and_1427_cse : STD_LOGIC;
  SIGNAL and_1429_cse : STD_LOGIC;
  SIGNAL and_1431_cse : STD_LOGIC;
  SIGNAL and_1433_cse : STD_LOGIC;
  SIGNAL and_1435_cse : STD_LOGIC;
  SIGNAL and_1437_cse : STD_LOGIC;
  SIGNAL and_1439_cse : STD_LOGIC;
  SIGNAL and_1441_cse : STD_LOGIC;
  SIGNAL and_1443_cse : STD_LOGIC;
  SIGNAL and_1445_cse : STD_LOGIC;
  SIGNAL and_1447_cse : STD_LOGIC;
  SIGNAL and_1449_cse : STD_LOGIC;
  SIGNAL and_1451_cse : STD_LOGIC;
  SIGNAL and_1453_cse : STD_LOGIC;
  SIGNAL and_1455_cse : STD_LOGIC;
  SIGNAL and_1457_cse : STD_LOGIC;
  SIGNAL and_1459_cse : STD_LOGIC;
  SIGNAL and_1461_cse : STD_LOGIC;
  SIGNAL and_1463_cse : STD_LOGIC;

  SIGNAL qelse_acc_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mux_13_nl : STD_LOGIC;
  SIGNAL mux_12_nl : STD_LOGIC;
  SIGNAL mux_11_nl : STD_LOGIC;
  SIGNAL mux_10_nl : STD_LOGIC;
  SIGNAL mux_9_nl : STD_LOGIC;
  SIGNAL mux_8_nl : STD_LOGIC;
  SIGNAL mux_7_nl : STD_LOGIC;
  SIGNAL mux_6_nl : STD_LOGIC;
  SIGNAL mux_5_nl : STD_LOGIC;
  SIGNAL mux_4_nl : STD_LOGIC;
  SIGNAL mux_3_nl : STD_LOGIC;
  SIGNAL mux_2_nl : STD_LOGIC;
  SIGNAL and_273_nl : STD_LOGIC;
  SIGNAL and_275_nl : STD_LOGIC;
  SIGNAL and_277_nl : STD_LOGIC;
  SIGNAL and_279_nl : STD_LOGIC;
  SIGNAL and_281_nl : STD_LOGIC;
  SIGNAL and_282_nl : STD_LOGIC;
  SIGNAL and_283_nl : STD_LOGIC;
  SIGNAL and_284_nl : STD_LOGIC;
  SIGNAL and_286_nl : STD_LOGIC;
  SIGNAL and_287_nl : STD_LOGIC;
  SIGNAL and_288_nl : STD_LOGIC;
  SIGNAL and_289_nl : STD_LOGIC;
  SIGNAL and_290_nl : STD_LOGIC;
  SIGNAL xor_nl : STD_LOGIC;
  SIGNAL nor_nl : STD_LOGIC;
  SIGNAL mux_14_nl : STD_LOGIC;
  SIGNAL nor_518_nl : STD_LOGIC;
  SIGNAL mux_15_nl : STD_LOGIC;
  SIGNAL nor_517_nl : STD_LOGIC;
  SIGNAL mux_16_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL mux_17_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL mux_18_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL mux_19_nl : STD_LOGIC;
  SIGNAL nor_512_nl : STD_LOGIC;
  SIGNAL mux_20_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL mux_22_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL mux_23_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL nor_506_nl : STD_LOGIC;
  SIGNAL mux_26_nl : STD_LOGIC;
  SIGNAL nor_507_nl : STD_LOGIC;
  SIGNAL mux_27_nl : STD_LOGIC;
  SIGNAL nor_508_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL or_61_nl : STD_LOGIC;
  SIGNAL nor_501_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL mux_31_nl : STD_LOGIC;
  SIGNAL nor_503_nl : STD_LOGIC;
  SIGNAL mux_32_nl : STD_LOGIC;
  SIGNAL nor_504_nl : STD_LOGIC;
  SIGNAL mux_33_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL and_1168_nl : STD_LOGIC;
  SIGNAL mux_35_nl : STD_LOGIC;
  SIGNAL nor_498_nl : STD_LOGIC;
  SIGNAL and_1166_nl : STD_LOGIC;
  SIGNAL and_1167_nl : STD_LOGIC;
  SIGNAL mux_38_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL and_1163_nl : STD_LOGIC;
  SIGNAL and_1164_nl : STD_LOGIC;
  SIGNAL and_1165_nl : STD_LOGIC;
  SIGNAL mux_42_nl : STD_LOGIC;
  SIGNAL nor_496_nl : STD_LOGIC;
  SIGNAL and_1159_nl : STD_LOGIC;
  SIGNAL and_1160_nl : STD_LOGIC;
  SIGNAL and_1161_nl : STD_LOGIC;
  SIGNAL and_1162_nl : STD_LOGIC;
  SIGNAL mux_47_nl : STD_LOGIC;
  SIGNAL nor_495_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL and_1155_nl : STD_LOGIC;
  SIGNAL and_1156_nl : STD_LOGIC;
  SIGNAL and_1157_nl : STD_LOGIC;
  SIGNAL and_1158_nl : STD_LOGIC;
  SIGNAL mux_53_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL nor_491_nl : STD_LOGIC;
  SIGNAL and_1151_nl : STD_LOGIC;
  SIGNAL and_1152_nl : STD_LOGIC;
  SIGNAL and_1153_nl : STD_LOGIC;
  SIGNAL and_1154_nl : STD_LOGIC;
  SIGNAL mux_60_nl : STD_LOGIC;
  SIGNAL nor_492_nl : STD_LOGIC;
  SIGNAL nor_486_nl : STD_LOGIC;
  SIGNAL nor_487_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL and_1147_nl : STD_LOGIC;
  SIGNAL and_1148_nl : STD_LOGIC;
  SIGNAL and_1149_nl : STD_LOGIC;
  SIGNAL and_1150_nl : STD_LOGIC;
  SIGNAL mux_68_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL nor_481_nl : STD_LOGIC;
  SIGNAL or_165_nl : STD_LOGIC;
  SIGNAL nor_482_nl : STD_LOGIC;
  SIGNAL nor_483_nl : STD_LOGIC;
  SIGNAL nor_484_nl : STD_LOGIC;
  SIGNAL and_1143_nl : STD_LOGIC;
  SIGNAL and_1144_nl : STD_LOGIC;
  SIGNAL and_1145_nl : STD_LOGIC;
  SIGNAL and_1146_nl : STD_LOGIC;
  SIGNAL mux_77_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL nor_480_nl : STD_LOGIC;
  SIGNAL or_175_nl : STD_LOGIC;
  SIGNAL mux_79_nl : STD_LOGIC;
  SIGNAL nor_479_nl : STD_LOGIC;
  SIGNAL mux_80_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL mux_81_nl : STD_LOGIC;
  SIGNAL nor_477_nl : STD_LOGIC;
  SIGNAL mux_82_nl : STD_LOGIC;
  SIGNAL nor_476_nl : STD_LOGIC;
  SIGNAL mux_83_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL mux_84_nl : STD_LOGIC;
  SIGNAL nor_473_nl : STD_LOGIC;
  SIGNAL mux_85_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL mux_87_nl : STD_LOGIC;
  SIGNAL nor_471_nl : STD_LOGIC;
  SIGNAL mux_88_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL nor_467_nl : STD_LOGIC;
  SIGNAL mux_91_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL mux_92_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL nor_461_nl : STD_LOGIC;
  SIGNAL or_250_nl : STD_LOGIC;
  SIGNAL nor_462_nl : STD_LOGIC;
  SIGNAL nor_463_nl : STD_LOGIC;
  SIGNAL mux_96_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL mux_97_nl : STD_LOGIC;
  SIGNAL nor_465_nl : STD_LOGIC;
  SIGNAL mux_98_nl : STD_LOGIC;
  SIGNAL nor_460_nl : STD_LOGIC;
  SIGNAL and_1142_nl : STD_LOGIC;
  SIGNAL mux_100_nl : STD_LOGIC;
  SIGNAL nor_459_nl : STD_LOGIC;
  SIGNAL and_1140_nl : STD_LOGIC;
  SIGNAL and_1141_nl : STD_LOGIC;
  SIGNAL mux_103_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL and_1137_nl : STD_LOGIC;
  SIGNAL and_1138_nl : STD_LOGIC;
  SIGNAL and_1139_nl : STD_LOGIC;
  SIGNAL mux_107_nl : STD_LOGIC;
  SIGNAL nor_457_nl : STD_LOGIC;
  SIGNAL and_1133_nl : STD_LOGIC;
  SIGNAL and_1134_nl : STD_LOGIC;
  SIGNAL and_1135_nl : STD_LOGIC;
  SIGNAL and_1136_nl : STD_LOGIC;
  SIGNAL mux_112_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL and_1129_nl : STD_LOGIC;
  SIGNAL and_1130_nl : STD_LOGIC;
  SIGNAL and_1131_nl : STD_LOGIC;
  SIGNAL and_1132_nl : STD_LOGIC;
  SIGNAL mux_118_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL nor_451_nl : STD_LOGIC;
  SIGNAL nor_452_nl : STD_LOGIC;
  SIGNAL and_1125_nl : STD_LOGIC;
  SIGNAL and_1126_nl : STD_LOGIC;
  SIGNAL and_1127_nl : STD_LOGIC;
  SIGNAL and_1128_nl : STD_LOGIC;
  SIGNAL mux_125_nl : STD_LOGIC;
  SIGNAL nor_453_nl : STD_LOGIC;
  SIGNAL nor_447_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL nor_449_nl : STD_LOGIC;
  SIGNAL and_1121_nl : STD_LOGIC;
  SIGNAL and_1122_nl : STD_LOGIC;
  SIGNAL and_1123_nl : STD_LOGIC;
  SIGNAL and_1124_nl : STD_LOGIC;
  SIGNAL mux_133_nl : STD_LOGIC;
  SIGNAL nor_450_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL or_352_nl : STD_LOGIC;
  SIGNAL nor_443_nl : STD_LOGIC;
  SIGNAL nor_444_nl : STD_LOGIC;
  SIGNAL nor_445_nl : STD_LOGIC;
  SIGNAL and_1117_nl : STD_LOGIC;
  SIGNAL and_1118_nl : STD_LOGIC;
  SIGNAL and_1119_nl : STD_LOGIC;
  SIGNAL and_1120_nl : STD_LOGIC;
  SIGNAL mux_142_nl : STD_LOGIC;
  SIGNAL nor_446_nl : STD_LOGIC;
  SIGNAL and_1116_nl : STD_LOGIC;
  SIGNAL or_362_nl : STD_LOGIC;
  SIGNAL mux_144_nl : STD_LOGIC;
  SIGNAL and_1172_nl : STD_LOGIC;
  SIGNAL mux_145_nl : STD_LOGIC;
  SIGNAL and_1114_nl : STD_LOGIC;
  SIGNAL mux_146_nl : STD_LOGIC;
  SIGNAL and_1113_nl : STD_LOGIC;
  SIGNAL mux_147_nl : STD_LOGIC;
  SIGNAL and_1112_nl : STD_LOGIC;
  SIGNAL mux_148_nl : STD_LOGIC;
  SIGNAL and_1111_nl : STD_LOGIC;
  SIGNAL mux_149_nl : STD_LOGIC;
  SIGNAL and_1109_nl : STD_LOGIC;
  SIGNAL mux_150_nl : STD_LOGIC;
  SIGNAL and_1110_nl : STD_LOGIC;
  SIGNAL and_1106_nl : STD_LOGIC;
  SIGNAL mux_152_nl : STD_LOGIC;
  SIGNAL and_1107_nl : STD_LOGIC;
  SIGNAL mux_153_nl : STD_LOGIC;
  SIGNAL and_1108_nl : STD_LOGIC;
  SIGNAL and_1102_nl : STD_LOGIC;
  SIGNAL and_1103_nl : STD_LOGIC;
  SIGNAL mux_156_nl : STD_LOGIC;
  SIGNAL and_1104_nl : STD_LOGIC;
  SIGNAL mux_157_nl : STD_LOGIC;
  SIGNAL and_1105_nl : STD_LOGIC;
  SIGNAL and_1097_nl : STD_LOGIC;
  SIGNAL or_437_nl : STD_LOGIC;
  SIGNAL and_1098_nl : STD_LOGIC;
  SIGNAL and_1099_nl : STD_LOGIC;
  SIGNAL mux_161_nl : STD_LOGIC;
  SIGNAL and_1100_nl : STD_LOGIC;
  SIGNAL mux_162_nl : STD_LOGIC;
  SIGNAL and_1101_nl : STD_LOGIC;
  SIGNAL mux_163_nl : STD_LOGIC;
  SIGNAL and_1171_nl : STD_LOGIC;
  SIGNAL and_1094_nl : STD_LOGIC;
  SIGNAL mux_165_nl : STD_LOGIC;
  SIGNAL and_1095_nl : STD_LOGIC;
  SIGNAL and_1091_nl : STD_LOGIC;
  SIGNAL and_1092_nl : STD_LOGIC;
  SIGNAL mux_168_nl : STD_LOGIC;
  SIGNAL and_1093_nl : STD_LOGIC;
  SIGNAL and_1087_nl : STD_LOGIC;
  SIGNAL and_1088_nl : STD_LOGIC;
  SIGNAL and_1089_nl : STD_LOGIC;
  SIGNAL mux_172_nl : STD_LOGIC;
  SIGNAL and_1090_nl : STD_LOGIC;
  SIGNAL and_1082_nl : STD_LOGIC;
  SIGNAL and_1083_nl : STD_LOGIC;
  SIGNAL and_1084_nl : STD_LOGIC;
  SIGNAL and_1085_nl : STD_LOGIC;
  SIGNAL mux_177_nl : STD_LOGIC;
  SIGNAL and_1086_nl : STD_LOGIC;
  SIGNAL and_1076_nl : STD_LOGIC;
  SIGNAL and_1077_nl : STD_LOGIC;
  SIGNAL and_1078_nl : STD_LOGIC;
  SIGNAL and_1079_nl : STD_LOGIC;
  SIGNAL and_1080_nl : STD_LOGIC;
  SIGNAL mux_183_nl : STD_LOGIC;
  SIGNAL and_1081_nl : STD_LOGIC;
  SIGNAL and_1069_nl : STD_LOGIC;
  SIGNAL and_1070_nl : STD_LOGIC;
  SIGNAL and_1071_nl : STD_LOGIC;
  SIGNAL and_1072_nl : STD_LOGIC;
  SIGNAL and_1073_nl : STD_LOGIC;
  SIGNAL and_1074_nl : STD_LOGIC;
  SIGNAL mux_190_nl : STD_LOGIC;
  SIGNAL and_1075_nl : STD_LOGIC;
  SIGNAL and_1061_nl : STD_LOGIC;
  SIGNAL and_1062_nl : STD_LOGIC;
  SIGNAL and_1063_nl : STD_LOGIC;
  SIGNAL and_1064_nl : STD_LOGIC;
  SIGNAL and_1065_nl : STD_LOGIC;
  SIGNAL and_1066_nl : STD_LOGIC;
  SIGNAL and_1067_nl : STD_LOGIC;
  SIGNAL mux_198_nl : STD_LOGIC;
  SIGNAL and_1068_nl : STD_LOGIC;
  SIGNAL and_1052_nl : STD_LOGIC;
  SIGNAL or_540_nl : STD_LOGIC;
  SIGNAL and_1053_nl : STD_LOGIC;
  SIGNAL and_1054_nl : STD_LOGIC;
  SIGNAL and_1055_nl : STD_LOGIC;
  SIGNAL and_1056_nl : STD_LOGIC;
  SIGNAL and_1057_nl : STD_LOGIC;
  SIGNAL and_1058_nl : STD_LOGIC;
  SIGNAL and_1059_nl : STD_LOGIC;
  SIGNAL mux_207_nl : STD_LOGIC;
  SIGNAL and_1060_nl : STD_LOGIC;
  SIGNAL nor_439_nl : STD_LOGIC;
  SIGNAL or_550_nl : STD_LOGIC;
  SIGNAL mux_209_nl : STD_LOGIC;
  SIGNAL and_1170_nl : STD_LOGIC;
  SIGNAL mux_210_nl : STD_LOGIC;
  SIGNAL and_1050_nl : STD_LOGIC;
  SIGNAL mux_211_nl : STD_LOGIC;
  SIGNAL and_1049_nl : STD_LOGIC;
  SIGNAL mux_212_nl : STD_LOGIC;
  SIGNAL and_1048_nl : STD_LOGIC;
  SIGNAL mux_213_nl : STD_LOGIC;
  SIGNAL and_1047_nl : STD_LOGIC;
  SIGNAL mux_214_nl : STD_LOGIC;
  SIGNAL and_1045_nl : STD_LOGIC;
  SIGNAL mux_215_nl : STD_LOGIC;
  SIGNAL and_1046_nl : STD_LOGIC;
  SIGNAL and_1042_nl : STD_LOGIC;
  SIGNAL mux_217_nl : STD_LOGIC;
  SIGNAL and_1043_nl : STD_LOGIC;
  SIGNAL mux_218_nl : STD_LOGIC;
  SIGNAL and_1044_nl : STD_LOGIC;
  SIGNAL and_1038_nl : STD_LOGIC;
  SIGNAL and_1039_nl : STD_LOGIC;
  SIGNAL mux_221_nl : STD_LOGIC;
  SIGNAL and_1040_nl : STD_LOGIC;
  SIGNAL mux_222_nl : STD_LOGIC;
  SIGNAL and_1041_nl : STD_LOGIC;
  SIGNAL and_1033_nl : STD_LOGIC;
  SIGNAL or_624_nl : STD_LOGIC;
  SIGNAL and_1034_nl : STD_LOGIC;
  SIGNAL and_1035_nl : STD_LOGIC;
  SIGNAL mux_226_nl : STD_LOGIC;
  SIGNAL and_1036_nl : STD_LOGIC;
  SIGNAL mux_227_nl : STD_LOGIC;
  SIGNAL and_1037_nl : STD_LOGIC;
  SIGNAL mux_228_nl : STD_LOGIC;
  SIGNAL and_1169_nl : STD_LOGIC;
  SIGNAL and_1030_nl : STD_LOGIC;
  SIGNAL mux_230_nl : STD_LOGIC;
  SIGNAL and_1031_nl : STD_LOGIC;
  SIGNAL and_1027_nl : STD_LOGIC;
  SIGNAL and_1028_nl : STD_LOGIC;
  SIGNAL mux_233_nl : STD_LOGIC;
  SIGNAL and_1029_nl : STD_LOGIC;
  SIGNAL and_1023_nl : STD_LOGIC;
  SIGNAL and_1024_nl : STD_LOGIC;
  SIGNAL and_1025_nl : STD_LOGIC;
  SIGNAL mux_237_nl : STD_LOGIC;
  SIGNAL and_1026_nl : STD_LOGIC;
  SIGNAL and_1018_nl : STD_LOGIC;
  SIGNAL and_1019_nl : STD_LOGIC;
  SIGNAL and_1020_nl : STD_LOGIC;
  SIGNAL and_1021_nl : STD_LOGIC;
  SIGNAL mux_242_nl : STD_LOGIC;
  SIGNAL and_1022_nl : STD_LOGIC;
  SIGNAL and_1012_nl : STD_LOGIC;
  SIGNAL and_1013_nl : STD_LOGIC;
  SIGNAL and_1014_nl : STD_LOGIC;
  SIGNAL and_1015_nl : STD_LOGIC;
  SIGNAL and_1016_nl : STD_LOGIC;
  SIGNAL mux_248_nl : STD_LOGIC;
  SIGNAL and_1017_nl : STD_LOGIC;
  SIGNAL and_1005_nl : STD_LOGIC;
  SIGNAL and_1006_nl : STD_LOGIC;
  SIGNAL and_1007_nl : STD_LOGIC;
  SIGNAL and_1008_nl : STD_LOGIC;
  SIGNAL and_1009_nl : STD_LOGIC;
  SIGNAL and_1010_nl : STD_LOGIC;
  SIGNAL mux_255_nl : STD_LOGIC;
  SIGNAL and_1011_nl : STD_LOGIC;
  SIGNAL and_997_nl : STD_LOGIC;
  SIGNAL and_998_nl : STD_LOGIC;
  SIGNAL and_999_nl : STD_LOGIC;
  SIGNAL and_1000_nl : STD_LOGIC;
  SIGNAL and_1001_nl : STD_LOGIC;
  SIGNAL and_1002_nl : STD_LOGIC;
  SIGNAL and_1003_nl : STD_LOGIC;
  SIGNAL mux_263_nl : STD_LOGIC;
  SIGNAL and_1004_nl : STD_LOGIC;
  SIGNAL and_988_nl : STD_LOGIC;
  SIGNAL or_725_nl : STD_LOGIC;
  SIGNAL and_989_nl : STD_LOGIC;
  SIGNAL and_990_nl : STD_LOGIC;
  SIGNAL and_991_nl : STD_LOGIC;
  SIGNAL and_992_nl : STD_LOGIC;
  SIGNAL and_993_nl : STD_LOGIC;
  SIGNAL and_994_nl : STD_LOGIC;
  SIGNAL and_995_nl : STD_LOGIC;
  SIGNAL mux_272_nl : STD_LOGIC;
  SIGNAL and_996_nl : STD_LOGIC;
  SIGNAL and_987_nl : STD_LOGIC;
  SIGNAL or_735_nl : STD_LOGIC;
  SIGNAL mux_274_nl : STD_LOGIC;
  SIGNAL nor_436_nl : STD_LOGIC;
  SIGNAL mux_275_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL mux_276_nl : STD_LOGIC;
  SIGNAL nor_434_nl : STD_LOGIC;
  SIGNAL mux_277_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL mux_278_nl : STD_LOGIC;
  SIGNAL nor_432_nl : STD_LOGIC;
  SIGNAL mux_279_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL mux_280_nl : STD_LOGIC;
  SIGNAL nor_431_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL mux_282_nl : STD_LOGIC;
  SIGNAL nor_428_nl : STD_LOGIC;
  SIGNAL mux_283_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL nor_423_nl : STD_LOGIC;
  SIGNAL nor_424_nl : STD_LOGIC;
  SIGNAL mux_286_nl : STD_LOGIC;
  SIGNAL nor_425_nl : STD_LOGIC;
  SIGNAL mux_287_nl : STD_LOGIC;
  SIGNAL nor_426_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL or_808_nl : STD_LOGIC;
  SIGNAL nor_419_nl : STD_LOGIC;
  SIGNAL nor_420_nl : STD_LOGIC;
  SIGNAL mux_291_nl : STD_LOGIC;
  SIGNAL nor_421_nl : STD_LOGIC;
  SIGNAL mux_292_nl : STD_LOGIC;
  SIGNAL nor_422_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL or_823_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL or_822_nl : STD_LOGIC;
  SIGNAL nor_411_nl : STD_LOGIC;
  SIGNAL or_821_nl : STD_LOGIC;
  SIGNAL nor_412_nl : STD_LOGIC;
  SIGNAL or_820_nl : STD_LOGIC;
  SIGNAL nor_413_nl : STD_LOGIC;
  SIGNAL or_819_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL or_818_nl : STD_LOGIC;
  SIGNAL nor_415_nl : STD_LOGIC;
  SIGNAL or_817_nl : STD_LOGIC;
  SIGNAL nor_416_nl : STD_LOGIC;
  SIGNAL or_816_nl : STD_LOGIC;
  SIGNAL mux_301_nl : STD_LOGIC;
  SIGNAL nor_417_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL mux_302_nl : STD_LOGIC;
  SIGNAL nor_408_nl : STD_LOGIC;
  SIGNAL and_986_nl : STD_LOGIC;
  SIGNAL mux_304_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL and_984_nl : STD_LOGIC;
  SIGNAL and_985_nl : STD_LOGIC;
  SIGNAL mux_307_nl : STD_LOGIC;
  SIGNAL nor_406_nl : STD_LOGIC;
  SIGNAL and_981_nl : STD_LOGIC;
  SIGNAL and_982_nl : STD_LOGIC;
  SIGNAL and_983_nl : STD_LOGIC;
  SIGNAL mux_311_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL and_977_nl : STD_LOGIC;
  SIGNAL and_978_nl : STD_LOGIC;
  SIGNAL and_979_nl : STD_LOGIC;
  SIGNAL and_980_nl : STD_LOGIC;
  SIGNAL mux_316_nl : STD_LOGIC;
  SIGNAL nor_404_nl : STD_LOGIC;
  SIGNAL nor_402_nl : STD_LOGIC;
  SIGNAL and_973_nl : STD_LOGIC;
  SIGNAL and_974_nl : STD_LOGIC;
  SIGNAL and_975_nl : STD_LOGIC;
  SIGNAL and_976_nl : STD_LOGIC;
  SIGNAL mux_322_nl : STD_LOGIC;
  SIGNAL nor_403_nl : STD_LOGIC;
  SIGNAL nor_399_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL and_969_nl : STD_LOGIC;
  SIGNAL and_970_nl : STD_LOGIC;
  SIGNAL and_971_nl : STD_LOGIC;
  SIGNAL and_972_nl : STD_LOGIC;
  SIGNAL mux_329_nl : STD_LOGIC;
  SIGNAL nor_401_nl : STD_LOGIC;
  SIGNAL nor_395_nl : STD_LOGIC;
  SIGNAL nor_396_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL and_965_nl : STD_LOGIC;
  SIGNAL and_966_nl : STD_LOGIC;
  SIGNAL and_967_nl : STD_LOGIC;
  SIGNAL and_968_nl : STD_LOGIC;
  SIGNAL mux_337_nl : STD_LOGIC;
  SIGNAL nor_398_nl : STD_LOGIC;
  SIGNAL nor_390_nl : STD_LOGIC;
  SIGNAL or_919_nl : STD_LOGIC;
  SIGNAL nor_391_nl : STD_LOGIC;
  SIGNAL nor_392_nl : STD_LOGIC;
  SIGNAL nor_393_nl : STD_LOGIC;
  SIGNAL and_961_nl : STD_LOGIC;
  SIGNAL and_962_nl : STD_LOGIC;
  SIGNAL and_963_nl : STD_LOGIC;
  SIGNAL and_964_nl : STD_LOGIC;
  SIGNAL mux_346_nl : STD_LOGIC;
  SIGNAL nor_394_nl : STD_LOGIC;
  SIGNAL nor_380_nl : STD_LOGIC;
  SIGNAL or_938_nl : STD_LOGIC;
  SIGNAL nor_381_nl : STD_LOGIC;
  SIGNAL or_937_nl : STD_LOGIC;
  SIGNAL nor_382_nl : STD_LOGIC;
  SIGNAL or_936_nl : STD_LOGIC;
  SIGNAL nor_383_nl : STD_LOGIC;
  SIGNAL or_935_nl : STD_LOGIC;
  SIGNAL nor_384_nl : STD_LOGIC;
  SIGNAL or_934_nl : STD_LOGIC;
  SIGNAL nor_385_nl : STD_LOGIC;
  SIGNAL or_933_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL or_932_nl : STD_LOGIC;
  SIGNAL nor_387_nl : STD_LOGIC;
  SIGNAL or_931_nl : STD_LOGIC;
  SIGNAL nor_388_nl : STD_LOGIC;
  SIGNAL or_930_nl : STD_LOGIC;
  SIGNAL nor_389_nl : STD_LOGIC;
  SIGNAL or_929_nl : STD_LOGIC;
  SIGNAL mux_357_nl : STD_LOGIC;
  SIGNAL nor_379_nl : STD_LOGIC;
  SIGNAL mux_358_nl : STD_LOGIC;
  SIGNAL nor_378_nl : STD_LOGIC;
  SIGNAL mux_359_nl : STD_LOGIC;
  SIGNAL nor_377_nl : STD_LOGIC;
  SIGNAL mux_360_nl : STD_LOGIC;
  SIGNAL nor_376_nl : STD_LOGIC;
  SIGNAL mux_361_nl : STD_LOGIC;
  SIGNAL nor_375_nl : STD_LOGIC;
  SIGNAL mux_362_nl : STD_LOGIC;
  SIGNAL nor_373_nl : STD_LOGIC;
  SIGNAL mux_363_nl : STD_LOGIC;
  SIGNAL nor_374_nl : STD_LOGIC;
  SIGNAL nor_370_nl : STD_LOGIC;
  SIGNAL mux_365_nl : STD_LOGIC;
  SIGNAL nor_371_nl : STD_LOGIC;
  SIGNAL mux_366_nl : STD_LOGIC;
  SIGNAL nor_372_nl : STD_LOGIC;
  SIGNAL nor_366_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL mux_369_nl : STD_LOGIC;
  SIGNAL nor_368_nl : STD_LOGIC;
  SIGNAL mux_370_nl : STD_LOGIC;
  SIGNAL nor_369_nl : STD_LOGIC;
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL or_1012_nl : STD_LOGIC;
  SIGNAL nor_362_nl : STD_LOGIC;
  SIGNAL nor_363_nl : STD_LOGIC;
  SIGNAL mux_374_nl : STD_LOGIC;
  SIGNAL nor_364_nl : STD_LOGIC;
  SIGNAL mux_375_nl : STD_LOGIC;
  SIGNAL nor_365_nl : STD_LOGIC;
  SIGNAL nor_352_nl : STD_LOGIC;
  SIGNAL or_1027_nl : STD_LOGIC;
  SIGNAL nor_353_nl : STD_LOGIC;
  SIGNAL or_1026_nl : STD_LOGIC;
  SIGNAL nor_354_nl : STD_LOGIC;
  SIGNAL or_1025_nl : STD_LOGIC;
  SIGNAL nor_355_nl : STD_LOGIC;
  SIGNAL or_1024_nl : STD_LOGIC;
  SIGNAL nor_356_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL nor_357_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL nor_358_nl : STD_LOGIC;
  SIGNAL or_1021_nl : STD_LOGIC;
  SIGNAL nor_359_nl : STD_LOGIC;
  SIGNAL or_1020_nl : STD_LOGIC;
  SIGNAL mux_384_nl : STD_LOGIC;
  SIGNAL nor_360_nl : STD_LOGIC;
  SIGNAL or_1019_nl : STD_LOGIC;
  SIGNAL mux_385_nl : STD_LOGIC;
  SIGNAL nor_351_nl : STD_LOGIC;
  SIGNAL and_960_nl : STD_LOGIC;
  SIGNAL mux_387_nl : STD_LOGIC;
  SIGNAL nor_350_nl : STD_LOGIC;
  SIGNAL and_958_nl : STD_LOGIC;
  SIGNAL and_959_nl : STD_LOGIC;
  SIGNAL mux_390_nl : STD_LOGIC;
  SIGNAL nor_349_nl : STD_LOGIC;
  SIGNAL and_955_nl : STD_LOGIC;
  SIGNAL and_956_nl : STD_LOGIC;
  SIGNAL and_957_nl : STD_LOGIC;
  SIGNAL mux_394_nl : STD_LOGIC;
  SIGNAL nor_348_nl : STD_LOGIC;
  SIGNAL and_951_nl : STD_LOGIC;
  SIGNAL and_952_nl : STD_LOGIC;
  SIGNAL and_953_nl : STD_LOGIC;
  SIGNAL and_954_nl : STD_LOGIC;
  SIGNAL mux_399_nl : STD_LOGIC;
  SIGNAL nor_347_nl : STD_LOGIC;
  SIGNAL nor_345_nl : STD_LOGIC;
  SIGNAL and_947_nl : STD_LOGIC;
  SIGNAL and_948_nl : STD_LOGIC;
  SIGNAL and_949_nl : STD_LOGIC;
  SIGNAL and_950_nl : STD_LOGIC;
  SIGNAL mux_405_nl : STD_LOGIC;
  SIGNAL nor_346_nl : STD_LOGIC;
  SIGNAL nor_342_nl : STD_LOGIC;
  SIGNAL nor_343_nl : STD_LOGIC;
  SIGNAL and_943_nl : STD_LOGIC;
  SIGNAL and_944_nl : STD_LOGIC;
  SIGNAL and_945_nl : STD_LOGIC;
  SIGNAL and_946_nl : STD_LOGIC;
  SIGNAL mux_412_nl : STD_LOGIC;
  SIGNAL nor_344_nl : STD_LOGIC;
  SIGNAL nor_338_nl : STD_LOGIC;
  SIGNAL nor_339_nl : STD_LOGIC;
  SIGNAL nor_340_nl : STD_LOGIC;
  SIGNAL and_939_nl : STD_LOGIC;
  SIGNAL and_940_nl : STD_LOGIC;
  SIGNAL and_941_nl : STD_LOGIC;
  SIGNAL and_942_nl : STD_LOGIC;
  SIGNAL mux_420_nl : STD_LOGIC;
  SIGNAL nor_341_nl : STD_LOGIC;
  SIGNAL nor_333_nl : STD_LOGIC;
  SIGNAL nand_12_nl : STD_LOGIC;
  SIGNAL nor_334_nl : STD_LOGIC;
  SIGNAL nor_335_nl : STD_LOGIC;
  SIGNAL nor_336_nl : STD_LOGIC;
  SIGNAL and_935_nl : STD_LOGIC;
  SIGNAL and_936_nl : STD_LOGIC;
  SIGNAL and_937_nl : STD_LOGIC;
  SIGNAL and_938_nl : STD_LOGIC;
  SIGNAL mux_429_nl : STD_LOGIC;
  SIGNAL nor_337_nl : STD_LOGIC;
  SIGNAL nor_324_nl : STD_LOGIC;
  SIGNAL nand_1_nl : STD_LOGIC;
  SIGNAL nor_325_nl : STD_LOGIC;
  SIGNAL nand_2_nl : STD_LOGIC;
  SIGNAL nor_326_nl : STD_LOGIC;
  SIGNAL nand_3_nl : STD_LOGIC;
  SIGNAL nor_327_nl : STD_LOGIC;
  SIGNAL nand_4_nl : STD_LOGIC;
  SIGNAL nor_328_nl : STD_LOGIC;
  SIGNAL nand_5_nl : STD_LOGIC;
  SIGNAL nor_329_nl : STD_LOGIC;
  SIGNAL nand_6_nl : STD_LOGIC;
  SIGNAL nor_330_nl : STD_LOGIC;
  SIGNAL nand_7_nl : STD_LOGIC;
  SIGNAL nor_331_nl : STD_LOGIC;
  SIGNAL nand_8_nl : STD_LOGIC;
  SIGNAL nor_332_nl : STD_LOGIC;
  SIGNAL nand_9_nl : STD_LOGIC;
  SIGNAL and_934_nl : STD_LOGIC;
  SIGNAL nand_11_nl : STD_LOGIC;
  SIGNAL base_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL base_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL m_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL m_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL return_rsci_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL return_rsci_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL ccs_ccore_start_rsci_dat : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL ccs_ccore_start_rsci_idat_1 : STD_LOGIC_VECTOR (0 DOWNTO 0);

  SIGNAL rem_13_cmp_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_1_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_1_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_1_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_2_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_2_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_2_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_3_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_3_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_3_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_4_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_4_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_4_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_5_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_5_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_5_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_6_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_6_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_6_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_7_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_7_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_7_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_8_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_8_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_8_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_9_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_9_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_9_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_10_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_10_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_10_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL rem_13_cmp_11_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_11_b : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL rem_13_cmp_11_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_v_64_11_2(input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_13_2(input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(12 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  base_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 1,
      width => 64
      )
    PORT MAP(
      dat => base_rsci_dat,
      idat => base_rsci_idat_1
    );
  base_rsci_dat <= base_rsc_dat;
  base_rsci_idat <= base_rsci_idat_1;

  m_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 64
      )
    PORT MAP(
      dat => m_rsci_dat,
      idat => m_rsci_idat_1
    );
  m_rsci_dat <= m_rsc_dat;
  m_rsci_idat <= m_rsci_idat_1;

  return_rsci : work.mgc_out_dreg_pkg_v2.mgc_out_dreg_v2
    GENERIC MAP(
      rscid => 3,
      width => 64
      )
    PORT MAP(
      d => return_rsci_d_1,
      z => return_rsci_z
    );
  return_rsci_d_1 <= return_rsci_d;
  return_rsc_z <= return_rsci_z;

  ccs_ccore_start_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 7,
      width => 1
      )
    PORT MAP(
      dat => ccs_ccore_start_rsci_dat,
      idat => ccs_ccore_start_rsci_idat_1
    );
  ccs_ccore_start_rsci_dat(0) <= ccs_ccore_start_rsc_dat;
  ccs_ccore_start_rsci_idat <= ccs_ccore_start_rsci_idat_1(0);

  rem_13_cmp : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_a,
      b => rem_13_cmp_b,
      z => rem_13_cmp_z_1
    );
  rem_13_cmp_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_a_63_0),65));
  rem_13_cmp_b <= '0' & rem_13_cmp_b_63_0;
  rem_13_cmp_z <= rem_13_cmp_z_1;

  rem_13_cmp_1 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_1_a,
      b => rem_13_cmp_1_b,
      z => rem_13_cmp_1_z_1
    );
  rem_13_cmp_1_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_1_a_63_0),65));
  rem_13_cmp_1_b <= '0' & rem_13_cmp_1_b_63_0;
  rem_13_cmp_1_z <= rem_13_cmp_1_z_1;

  rem_13_cmp_2 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_2_a,
      b => rem_13_cmp_2_b,
      z => rem_13_cmp_2_z_1
    );
  rem_13_cmp_2_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_2_a_63_0),65));
  rem_13_cmp_2_b <= '0' & rem_13_cmp_2_b_63_0;
  rem_13_cmp_2_z <= rem_13_cmp_2_z_1;

  rem_13_cmp_3 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_3_a,
      b => rem_13_cmp_3_b,
      z => rem_13_cmp_3_z_1
    );
  rem_13_cmp_3_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_3_a_63_0),65));
  rem_13_cmp_3_b <= '0' & rem_13_cmp_3_b_63_0;
  rem_13_cmp_3_z <= rem_13_cmp_3_z_1;

  rem_13_cmp_4 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_4_a,
      b => rem_13_cmp_4_b,
      z => rem_13_cmp_4_z_1
    );
  rem_13_cmp_4_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_4_a_63_0),65));
  rem_13_cmp_4_b <= '0' & rem_13_cmp_4_b_63_0;
  rem_13_cmp_4_z <= rem_13_cmp_4_z_1;

  rem_13_cmp_5 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_5_a,
      b => rem_13_cmp_5_b,
      z => rem_13_cmp_5_z_1
    );
  rem_13_cmp_5_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_5_a_63_0),65));
  rem_13_cmp_5_b <= '0' & rem_13_cmp_5_b_63_0;
  rem_13_cmp_5_z <= rem_13_cmp_5_z_1;

  rem_13_cmp_6 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_6_a,
      b => rem_13_cmp_6_b,
      z => rem_13_cmp_6_z_1
    );
  rem_13_cmp_6_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_6_a_63_0),65));
  rem_13_cmp_6_b <= '0' & rem_13_cmp_6_b_63_0;
  rem_13_cmp_6_z <= rem_13_cmp_6_z_1;

  rem_13_cmp_7 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_7_a,
      b => rem_13_cmp_7_b,
      z => rem_13_cmp_7_z_1
    );
  rem_13_cmp_7_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_7_a_63_0),65));
  rem_13_cmp_7_b <= '0' & rem_13_cmp_7_b_63_0;
  rem_13_cmp_7_z <= rem_13_cmp_7_z_1;

  rem_13_cmp_8 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_8_a,
      b => rem_13_cmp_8_b,
      z => rem_13_cmp_8_z_1
    );
  rem_13_cmp_8_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_8_a_63_0),65));
  rem_13_cmp_8_b <= '0' & rem_13_cmp_8_b_63_0;
  rem_13_cmp_8_z <= rem_13_cmp_8_z_1;

  rem_13_cmp_9 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_9_a,
      b => rem_13_cmp_9_b,
      z => rem_13_cmp_9_z_1
    );
  rem_13_cmp_9_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_9_a_63_0),65));
  rem_13_cmp_9_b <= '0' & rem_13_cmp_9_b_63_0;
  rem_13_cmp_9_z <= rem_13_cmp_9_z_1;

  rem_13_cmp_10 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_10_a,
      b => rem_13_cmp_10_b,
      z => rem_13_cmp_10_z_1
    );
  rem_13_cmp_10_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_10_a_63_0),65));
  rem_13_cmp_10_b <= '0' & rem_13_cmp_10_b_63_0;
  rem_13_cmp_10_z <= rem_13_cmp_10_z_1;

  rem_13_cmp_11 : work.mgc_comps.mgc_rem
    GENERIC MAP(
      width_a => 65,
      width_b => 65,
      signd => 1
      )
    PORT MAP(
      a => rem_13_cmp_11_a,
      b => rem_13_cmp_11_b,
      z => rem_13_cmp_11_z_1
    );
  rem_13_cmp_11_a <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(rem_13_cmp_11_a_63_0),65));
  rem_13_cmp_11_b <= '0' & rem_13_cmp_11_b_63_0;
  rem_13_cmp_11_z <= rem_13_cmp_11_z_1;

  and_1203_cse <= ccs_ccore_en AND main_stage_0_12 AND asn_itm_11;
  and_1173_cse <= ccs_ccore_en AND (and_dcpl_294 OR and_dcpl_300 OR and_dcpl_306
      OR and_dcpl_312 OR and_dcpl_318 OR and_dcpl_324 OR and_dcpl_330 OR and_dcpl_336
      OR and_dcpl_342 OR and_dcpl_348 OR and_tmp_35);
  and_1175_cse <= ccs_ccore_en AND (and_dcpl_356 OR and_dcpl_360 OR and_dcpl_364
      OR and_dcpl_368 OR and_dcpl_372 OR and_dcpl_376 OR and_dcpl_379 OR and_dcpl_382
      OR and_dcpl_385 OR and_dcpl_388 OR mux_tmp_76);
  and_1177_cse <= ccs_ccore_en AND (and_dcpl_394 OR and_dcpl_397 OR and_dcpl_400
      OR and_dcpl_403 OR and_dcpl_406 OR and_dcpl_409 OR and_dcpl_413 OR and_dcpl_417
      OR and_dcpl_421 OR and_dcpl_425 OR and_tmp_80);
  and_1179_cse <= ccs_ccore_en AND (and_dcpl_431 OR and_dcpl_433 OR and_dcpl_435
      OR and_dcpl_437 OR and_dcpl_439 OR and_dcpl_442 OR and_dcpl_445 OR and_dcpl_448
      OR and_dcpl_451 OR and_dcpl_454 OR mux_tmp_141);
  and_1181_cse <= ccs_ccore_en AND (and_dcpl_461 OR and_dcpl_465 OR and_dcpl_469
      OR and_dcpl_473 OR and_dcpl_477 OR and_dcpl_480 OR and_dcpl_483 OR and_dcpl_486
      OR and_dcpl_489 OR and_dcpl_492 OR and_tmp_125);
  and_1183_cse <= ccs_ccore_en AND (and_dcpl_498 OR and_dcpl_500 OR and_dcpl_502
      OR and_dcpl_504 OR and_dcpl_506 OR and_dcpl_508 OR and_dcpl_510 OR and_dcpl_512
      OR and_dcpl_514 OR and_dcpl_516 OR mux_tmp_206);
  and_1185_cse <= ccs_ccore_en AND (and_dcpl_520 OR and_dcpl_523 OR and_dcpl_526
      OR and_dcpl_529 OR and_dcpl_532 OR and_dcpl_534 OR and_dcpl_536 OR and_dcpl_538
      OR and_dcpl_540 OR and_dcpl_542 OR and_tmp_170);
  and_1187_cse <= ccs_ccore_en AND (and_dcpl_546 OR and_dcpl_548 OR and_dcpl_550
      OR and_dcpl_552 OR and_dcpl_554 OR and_dcpl_556 OR and_dcpl_558 OR and_dcpl_560
      OR and_dcpl_562 OR and_dcpl_564 OR mux_tmp_271);
  and_1189_cse <= ccs_ccore_en AND (and_dcpl_569 OR and_dcpl_573 OR and_dcpl_577
      OR and_dcpl_581 OR and_dcpl_585 OR and_dcpl_589 OR and_dcpl_593 OR and_dcpl_597
      OR and_dcpl_601 OR and_dcpl_605 OR and_tmp_206);
  and_1191_cse <= ccs_ccore_en AND (and_dcpl_610 OR and_dcpl_612 OR and_dcpl_614
      OR and_dcpl_616 OR and_dcpl_618 OR and_dcpl_622 OR and_dcpl_625 OR and_dcpl_628
      OR and_dcpl_631 OR and_dcpl_634 OR mux_tmp_354);
  and_1193_cse <= ccs_ccore_en AND (and_dcpl_638 OR and_dcpl_641 OR and_dcpl_644
      OR and_dcpl_647 OR and_dcpl_650 OR and_dcpl_653 OR and_dcpl_657 OR and_dcpl_661
      OR and_dcpl_665 OR and_dcpl_669 OR and_tmp_233);
  and_1195_cse <= ccs_ccore_en AND (and_dcpl_673 OR and_dcpl_675 OR and_dcpl_677
      OR and_dcpl_679 OR and_dcpl_681 OR and_dcpl_684 OR and_dcpl_687 OR and_dcpl_690
      OR and_dcpl_693 OR and_dcpl_696 OR mux_tmp_437);
  and_1205_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_2;
  and_1207_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_6;
  and_1209_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_9;
  and_1211_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_11;
  and_1213_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_2;
  and_1215_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_6;
  and_1217_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_9;
  and_1219_cse <= ccs_ccore_en AND and_dcpl_13 AND and_dcpl_11;
  and_1221_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_1223_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_18 AND (rem_12cyc_st_10_1_0(0));
  and_1225_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_23 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_1227_cse <= ccs_ccore_en AND and_dcpl_4 AND and_dcpl_23 AND (rem_12cyc_st_10_1_0(0));
  and_1229_cse <= ccs_ccore_en AND and_dcpl_3;
  and_1231_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_29;
  and_1233_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_33;
  and_1235_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_36;
  and_1237_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_38;
  and_1239_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_29;
  and_1241_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_33;
  and_1243_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_36;
  and_1245_cse <= ccs_ccore_en AND and_dcpl_40 AND and_dcpl_38;
  and_1247_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_45 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_1249_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_45 AND (rem_12cyc_st_9_1_0(0));
  and_1251_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_50 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_1253_cse <= ccs_ccore_en AND and_dcpl_31 AND and_dcpl_50 AND (rem_12cyc_st_9_1_0(0));
  and_1255_cse <= ccs_ccore_en AND and_dcpl_30;
  and_1257_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_56;
  and_1259_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_60;
  and_1261_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_63;
  and_1263_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_65;
  and_1265_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_56;
  and_1267_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_60;
  and_1269_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_63;
  and_1271_cse <= ccs_ccore_en AND and_dcpl_67 AND and_dcpl_65;
  and_1273_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_72 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_1275_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_72 AND (rem_12cyc_st_8_1_0(0));
  and_1277_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_77 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_1279_cse <= ccs_ccore_en AND and_dcpl_58 AND and_dcpl_77 AND (rem_12cyc_st_8_1_0(0));
  and_1281_cse <= ccs_ccore_en AND and_dcpl_57;
  and_1283_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_83;
  and_1285_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_87;
  and_1287_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_90;
  and_1289_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_92;
  and_1291_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_83;
  and_1293_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_87;
  and_1295_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_90;
  and_1297_cse <= ccs_ccore_en AND and_dcpl_94 AND and_dcpl_92;
  and_1299_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_99 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_1301_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_99 AND (rem_12cyc_st_7_1_0(0));
  and_1303_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_104 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_1305_cse <= ccs_ccore_en AND and_dcpl_85 AND and_dcpl_104 AND (rem_12cyc_st_7_1_0(0));
  and_1307_cse <= ccs_ccore_en AND and_dcpl_84;
  and_1309_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_110;
  and_1311_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_115;
  and_1313_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_117;
  and_1315_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_119;
  and_1317_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_110;
  and_1319_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_115;
  and_1321_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_117;
  and_1323_cse <= ccs_ccore_en AND and_dcpl_121 AND and_dcpl_119;
  and_1325_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_126 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_1327_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_129 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_1329_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_126 AND (rem_12cyc_st_6_1_0(1));
  and_1331_cse <= ccs_ccore_en AND and_dcpl_112 AND and_dcpl_129 AND (rem_12cyc_st_6_1_0(1));
  and_1333_cse <= ccs_ccore_en AND and_dcpl_111;
  and_1335_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_137;
  and_1337_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_141;
  and_1339_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_144;
  and_1341_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_146;
  and_1343_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_137;
  and_1345_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_141;
  and_1347_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_144;
  and_1349_cse <= ccs_ccore_en AND and_dcpl_148 AND and_dcpl_146;
  and_1351_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_153 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_1353_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_153 AND (rem_12cyc_st_5_1_0(0));
  and_1355_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_158 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_1357_cse <= ccs_ccore_en AND and_dcpl_139 AND and_dcpl_158 AND (rem_12cyc_st_5_1_0(0));
  and_1359_cse <= ccs_ccore_en AND and_dcpl_138;
  and_1361_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_164;
  and_1363_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_168;
  and_1365_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_171;
  and_1367_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_173;
  and_1369_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_175 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_1371_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_175 AND (rem_12cyc_st_4_1_0(0));
  and_1373_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_180 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_1375_cse <= ccs_ccore_en AND and_dcpl_166 AND and_dcpl_180 AND (rem_12cyc_st_4_1_0(0));
  and_1377_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_164;
  and_1379_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_168;
  and_1381_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_171;
  and_1383_cse <= ccs_ccore_en AND and_dcpl_185 AND and_dcpl_173;
  and_1385_cse <= ccs_ccore_en AND and_dcpl_165;
  and_1387_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_191;
  and_1389_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_195;
  and_1391_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_198;
  and_1393_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_200;
  and_1395_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_191;
  and_1397_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_195;
  and_1399_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_198;
  and_1401_cse <= ccs_ccore_en AND and_dcpl_202 AND and_dcpl_200;
  and_1403_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_207 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_1405_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_207 AND (rem_12cyc_st_3_1_0(0));
  and_1407_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_212 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_1409_cse <= ccs_ccore_en AND and_dcpl_193 AND and_dcpl_212 AND (rem_12cyc_st_3_1_0(0));
  and_1411_cse <= ccs_ccore_en AND and_dcpl_192;
  and_1413_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_218;
  and_1415_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_222;
  and_1417_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_225;
  and_1419_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_227;
  and_1421_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_229 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_1423_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_229 AND (rem_12cyc_st_2_1_0(0));
  and_1425_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_234 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_1427_cse <= ccs_ccore_en AND and_dcpl_220 AND and_dcpl_234 AND (rem_12cyc_st_2_1_0(0));
  and_1429_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_218;
  and_1431_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_222;
  and_1433_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_225;
  and_1435_cse <= ccs_ccore_en AND and_dcpl_239 AND and_dcpl_227;
  and_1437_cse <= ccs_ccore_en AND and_dcpl_219;
  and_1439_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_245;
  and_1441_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_249;
  and_1443_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_252;
  and_1445_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_254;
  and_1447_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_245;
  and_1449_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_249;
  and_1451_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_252;
  and_1453_cse <= ccs_ccore_en AND and_dcpl_256 AND and_dcpl_254;
  and_1455_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_261 AND (NOT (rem_12cyc_1_0(0)));
  and_1457_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_261 AND (rem_12cyc_1_0(0));
  and_1459_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_266 AND (NOT (rem_12cyc_1_0(0)));
  and_1461_cse <= ccs_ccore_en AND and_dcpl_247 AND and_dcpl_266 AND (rem_12cyc_1_0(0));
  and_1463_cse <= ccs_ccore_en AND and_dcpl_246;
  and_1197_cse <= ccs_ccore_en AND ccs_ccore_start_rsci_idat;
  and_273_nl <= and_dcpl_272 AND and_dcpl_271;
  and_275_nl <= and_dcpl_272 AND and_dcpl_274;
  and_277_nl <= and_dcpl_272 AND and_dcpl_276;
  and_279_nl <= and_dcpl_272 AND and_dcpl_278;
  and_281_nl <= and_dcpl_280 AND and_dcpl_271;
  and_282_nl <= and_dcpl_280 AND and_dcpl_274;
  and_283_nl <= and_dcpl_280 AND and_dcpl_276;
  and_284_nl <= and_dcpl_280 AND and_dcpl_278;
  and_286_nl <= and_dcpl_285 AND and_dcpl_271;
  and_287_nl <= and_dcpl_285 AND and_dcpl_274;
  and_288_nl <= and_dcpl_285 AND and_dcpl_276;
  and_289_nl <= and_dcpl_285 AND and_dcpl_278;
  and_290_nl <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("11"));
  result_sva_duc_mx0 <= MUX1HOT_v_64_13_2((rem_13_cmp_1_z(63 DOWNTO 0)), (rem_13_cmp_2_z(63
      DOWNTO 0)), (rem_13_cmp_3_z(63 DOWNTO 0)), (rem_13_cmp_4_z(63 DOWNTO 0)), (rem_13_cmp_5_z(63
      DOWNTO 0)), (rem_13_cmp_6_z(63 DOWNTO 0)), (rem_13_cmp_7_z(63 DOWNTO 0)), (rem_13_cmp_8_z(63
      DOWNTO 0)), (rem_13_cmp_9_z(63 DOWNTO 0)), (rem_13_cmp_10_z(63 DOWNTO 0)),
      (rem_13_cmp_11_z(63 DOWNTO 0)), (rem_13_cmp_z(63 DOWNTO 0)), result_sva_duc,
      STD_LOGIC_VECTOR'( and_273_nl & and_275_nl & and_277_nl & and_279_nl & and_281_nl
      & and_282_nl & and_283_nl & and_284_nl & and_286_nl & and_287_nl & and_288_nl
      & and_289_nl & and_290_nl));
  acc_1_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(rem_12cyc_3_2 & rem_12cyc_1_0)
      + UNSIGNED'( "0001"), 4));
  xor_nl <= (acc_1_tmp(2)) XOR (acc_1_tmp(3));
  nor_nl <= NOT(CONV_SL_1_1(acc_1_tmp(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")));
  acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(xor_nl, 1),
      2) + CONV_UNSIGNED(CONV_UNSIGNED(nor_nl, 1), 2), 2));
  and_dcpl_1 <= NOT((rem_12cyc_st_10_3_2(1)) OR (rem_12cyc_st_10_1_0(1)));
  and_dcpl_2 <= and_dcpl_1 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_dcpl_3 <= main_stage_0_11 AND asn_itm_10;
  and_dcpl_4 <= and_dcpl_3 AND (NOT (rem_12cyc_st_10_3_2(0)));
  and_dcpl_6 <= and_dcpl_1 AND (rem_12cyc_st_10_1_0(0));
  and_dcpl_8 <= (NOT (rem_12cyc_st_10_3_2(1))) AND (rem_12cyc_st_10_1_0(1));
  and_dcpl_9 <= and_dcpl_8 AND (NOT (rem_12cyc_st_10_1_0(0)));
  and_dcpl_11 <= and_dcpl_8 AND (rem_12cyc_st_10_1_0(0));
  and_dcpl_13 <= and_dcpl_3 AND (rem_12cyc_st_10_3_2(0));
  and_dcpl_18 <= (rem_12cyc_st_10_3_2(1)) AND (NOT (rem_12cyc_st_10_1_0(1)));
  and_dcpl_23 <= (rem_12cyc_st_10_3_2(1)) AND (rem_12cyc_st_10_1_0(1));
  and_dcpl_28 <= NOT((rem_12cyc_st_9_3_2(1)) OR (rem_12cyc_st_9_1_0(1)));
  and_dcpl_29 <= and_dcpl_28 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_dcpl_30 <= main_stage_0_10 AND asn_itm_9;
  and_dcpl_31 <= and_dcpl_30 AND (NOT (rem_12cyc_st_9_3_2(0)));
  and_dcpl_33 <= and_dcpl_28 AND (rem_12cyc_st_9_1_0(0));
  and_dcpl_35 <= (NOT (rem_12cyc_st_9_3_2(1))) AND (rem_12cyc_st_9_1_0(1));
  and_dcpl_36 <= and_dcpl_35 AND (NOT (rem_12cyc_st_9_1_0(0)));
  and_dcpl_38 <= and_dcpl_35 AND (rem_12cyc_st_9_1_0(0));
  and_dcpl_40 <= and_dcpl_30 AND (rem_12cyc_st_9_3_2(0));
  and_dcpl_45 <= (rem_12cyc_st_9_3_2(1)) AND (NOT (rem_12cyc_st_9_1_0(1)));
  and_dcpl_50 <= (rem_12cyc_st_9_3_2(1)) AND (rem_12cyc_st_9_1_0(1));
  and_dcpl_55 <= NOT((rem_12cyc_st_8_3_2(1)) OR (rem_12cyc_st_8_1_0(1)));
  and_dcpl_56 <= and_dcpl_55 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_dcpl_57 <= main_stage_0_9 AND asn_itm_8;
  and_dcpl_58 <= and_dcpl_57 AND (NOT (rem_12cyc_st_8_3_2(0)));
  and_dcpl_60 <= and_dcpl_55 AND (rem_12cyc_st_8_1_0(0));
  and_dcpl_62 <= (NOT (rem_12cyc_st_8_3_2(1))) AND (rem_12cyc_st_8_1_0(1));
  and_dcpl_63 <= and_dcpl_62 AND (NOT (rem_12cyc_st_8_1_0(0)));
  and_dcpl_65 <= and_dcpl_62 AND (rem_12cyc_st_8_1_0(0));
  and_dcpl_67 <= and_dcpl_57 AND (rem_12cyc_st_8_3_2(0));
  and_dcpl_72 <= (rem_12cyc_st_8_3_2(1)) AND (NOT (rem_12cyc_st_8_1_0(1)));
  and_dcpl_77 <= (rem_12cyc_st_8_3_2(1)) AND (rem_12cyc_st_8_1_0(1));
  and_dcpl_82 <= NOT((rem_12cyc_st_7_3_2(1)) OR (rem_12cyc_st_7_1_0(1)));
  and_dcpl_83 <= and_dcpl_82 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_dcpl_84 <= main_stage_0_8 AND asn_itm_7;
  and_dcpl_85 <= and_dcpl_84 AND (NOT (rem_12cyc_st_7_3_2(0)));
  and_dcpl_87 <= and_dcpl_82 AND (rem_12cyc_st_7_1_0(0));
  and_dcpl_89 <= (NOT (rem_12cyc_st_7_3_2(1))) AND (rem_12cyc_st_7_1_0(1));
  and_dcpl_90 <= and_dcpl_89 AND (NOT (rem_12cyc_st_7_1_0(0)));
  and_dcpl_92 <= and_dcpl_89 AND (rem_12cyc_st_7_1_0(0));
  and_dcpl_94 <= and_dcpl_84 AND (rem_12cyc_st_7_3_2(0));
  and_dcpl_99 <= (rem_12cyc_st_7_3_2(1)) AND (NOT (rem_12cyc_st_7_1_0(1)));
  and_dcpl_104 <= (rem_12cyc_st_7_3_2(1)) AND (rem_12cyc_st_7_1_0(1));
  and_dcpl_109 <= NOT((rem_12cyc_st_6_3_2(1)) OR (rem_12cyc_st_6_1_0(0)));
  and_dcpl_110 <= and_dcpl_109 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_dcpl_111 <= main_stage_0_7 AND asn_itm_6;
  and_dcpl_112 <= and_dcpl_111 AND (NOT (rem_12cyc_st_6_3_2(0)));
  and_dcpl_114 <= (NOT (rem_12cyc_st_6_3_2(1))) AND (rem_12cyc_st_6_1_0(0));
  and_dcpl_115 <= and_dcpl_114 AND (NOT (rem_12cyc_st_6_1_0(1)));
  and_dcpl_117 <= and_dcpl_109 AND (rem_12cyc_st_6_1_0(1));
  and_dcpl_119 <= and_dcpl_114 AND (rem_12cyc_st_6_1_0(1));
  and_dcpl_121 <= and_dcpl_111 AND (rem_12cyc_st_6_3_2(0));
  and_dcpl_126 <= (rem_12cyc_st_6_3_2(1)) AND (NOT (rem_12cyc_st_6_1_0(0)));
  and_dcpl_129 <= (rem_12cyc_st_6_3_2(1)) AND (rem_12cyc_st_6_1_0(0));
  and_dcpl_136 <= NOT((rem_12cyc_st_5_3_2(1)) OR (rem_12cyc_st_5_1_0(1)));
  and_dcpl_137 <= and_dcpl_136 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_dcpl_138 <= main_stage_0_6 AND asn_itm_5;
  and_dcpl_139 <= and_dcpl_138 AND (NOT (rem_12cyc_st_5_3_2(0)));
  and_dcpl_141 <= and_dcpl_136 AND (rem_12cyc_st_5_1_0(0));
  and_dcpl_143 <= (NOT (rem_12cyc_st_5_3_2(1))) AND (rem_12cyc_st_5_1_0(1));
  and_dcpl_144 <= and_dcpl_143 AND (NOT (rem_12cyc_st_5_1_0(0)));
  and_dcpl_146 <= and_dcpl_143 AND (rem_12cyc_st_5_1_0(0));
  and_dcpl_148 <= and_dcpl_138 AND (rem_12cyc_st_5_3_2(0));
  and_dcpl_153 <= (rem_12cyc_st_5_3_2(1)) AND (NOT (rem_12cyc_st_5_1_0(1)));
  and_dcpl_158 <= (rem_12cyc_st_5_3_2(1)) AND (rem_12cyc_st_5_1_0(1));
  and_dcpl_163 <= NOT((rem_12cyc_st_4_3_2(0)) OR (rem_12cyc_st_4_1_0(1)));
  and_dcpl_164 <= and_dcpl_163 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_dcpl_165 <= main_stage_0_5 AND asn_itm_4;
  and_dcpl_166 <= and_dcpl_165 AND (NOT (rem_12cyc_st_4_3_2(1)));
  and_dcpl_168 <= and_dcpl_163 AND (rem_12cyc_st_4_1_0(0));
  and_dcpl_170 <= (NOT (rem_12cyc_st_4_3_2(0))) AND (rem_12cyc_st_4_1_0(1));
  and_dcpl_171 <= and_dcpl_170 AND (NOT (rem_12cyc_st_4_1_0(0)));
  and_dcpl_173 <= and_dcpl_170 AND (rem_12cyc_st_4_1_0(0));
  and_dcpl_175 <= (rem_12cyc_st_4_3_2(0)) AND (NOT (rem_12cyc_st_4_1_0(1)));
  and_dcpl_180 <= (rem_12cyc_st_4_3_2(0)) AND (rem_12cyc_st_4_1_0(1));
  and_dcpl_185 <= and_dcpl_165 AND (rem_12cyc_st_4_3_2(1));
  and_dcpl_190 <= NOT((rem_12cyc_st_3_3_2(1)) OR (rem_12cyc_st_3_1_0(1)));
  and_dcpl_191 <= and_dcpl_190 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_dcpl_192 <= main_stage_0_4 AND asn_itm_3;
  and_dcpl_193 <= and_dcpl_192 AND (NOT (rem_12cyc_st_3_3_2(0)));
  and_dcpl_195 <= and_dcpl_190 AND (rem_12cyc_st_3_1_0(0));
  and_dcpl_197 <= (NOT (rem_12cyc_st_3_3_2(1))) AND (rem_12cyc_st_3_1_0(1));
  and_dcpl_198 <= and_dcpl_197 AND (NOT (rem_12cyc_st_3_1_0(0)));
  and_dcpl_200 <= and_dcpl_197 AND (rem_12cyc_st_3_1_0(0));
  and_dcpl_202 <= and_dcpl_192 AND (rem_12cyc_st_3_3_2(0));
  and_dcpl_207 <= (rem_12cyc_st_3_3_2(1)) AND (NOT (rem_12cyc_st_3_1_0(1)));
  and_dcpl_212 <= (rem_12cyc_st_3_3_2(1)) AND (rem_12cyc_st_3_1_0(1));
  and_dcpl_217 <= NOT((rem_12cyc_st_2_3_2(0)) OR (rem_12cyc_st_2_1_0(1)));
  and_dcpl_218 <= and_dcpl_217 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_dcpl_219 <= main_stage_0_3 AND asn_itm_2;
  and_dcpl_220 <= and_dcpl_219 AND (NOT (rem_12cyc_st_2_3_2(1)));
  and_dcpl_222 <= and_dcpl_217 AND (rem_12cyc_st_2_1_0(0));
  and_dcpl_224 <= (NOT (rem_12cyc_st_2_3_2(0))) AND (rem_12cyc_st_2_1_0(1));
  and_dcpl_225 <= and_dcpl_224 AND (NOT (rem_12cyc_st_2_1_0(0)));
  and_dcpl_227 <= and_dcpl_224 AND (rem_12cyc_st_2_1_0(0));
  and_dcpl_229 <= (rem_12cyc_st_2_3_2(0)) AND (NOT (rem_12cyc_st_2_1_0(1)));
  and_dcpl_234 <= (rem_12cyc_st_2_3_2(0)) AND (rem_12cyc_st_2_1_0(1));
  and_dcpl_239 <= and_dcpl_219 AND (rem_12cyc_st_2_3_2(1));
  and_dcpl_244 <= NOT((rem_12cyc_3_2(1)) OR (rem_12cyc_1_0(1)));
  and_dcpl_245 <= and_dcpl_244 AND (NOT (rem_12cyc_1_0(0)));
  and_dcpl_246 <= main_stage_0_2 AND asn_itm_1;
  and_dcpl_247 <= and_dcpl_246 AND (NOT (rem_12cyc_3_2(0)));
  and_dcpl_249 <= and_dcpl_244 AND (rem_12cyc_1_0(0));
  and_dcpl_251 <= (NOT (rem_12cyc_3_2(1))) AND (rem_12cyc_1_0(1));
  and_dcpl_252 <= and_dcpl_251 AND (NOT (rem_12cyc_1_0(0)));
  and_dcpl_254 <= and_dcpl_251 AND (rem_12cyc_1_0(0));
  and_dcpl_256 <= and_dcpl_246 AND (rem_12cyc_3_2(0));
  and_dcpl_261 <= (rem_12cyc_3_2(1)) AND (NOT (rem_12cyc_1_0(1)));
  and_dcpl_266 <= (rem_12cyc_3_2(1)) AND (rem_12cyc_1_0(1));
  and_dcpl_271 <= NOT(CONV_SL_1_1(rem_12cyc_st_12_1_0/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_272 <= NOT(CONV_SL_1_1(rem_12cyc_st_12_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_274 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("01"));
  and_dcpl_276 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("10"));
  and_dcpl_278 <= CONV_SL_1_1(rem_12cyc_st_12_1_0=STD_LOGIC_VECTOR'("11"));
  and_dcpl_280 <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_285 <= CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_291 <= NOT(CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_292 <= ccs_ccore_start_rsci_idat AND (NOT (acc_tmp(0)));
  and_dcpl_293 <= and_dcpl_292 AND (NOT (acc_tmp(1)));
  and_dcpl_294 <= and_dcpl_293 AND and_dcpl_291;
  and_dcpl_295 <= NOT(CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_296 <= and_dcpl_295 AND (NOT (rem_12cyc_st_2_1_0(1)));
  and_dcpl_298 <= (NOT (rem_12cyc_st_2_1_0(0))) AND main_stage_0_3 AND asn_itm_2;
  not_tmp_54 <= NOT(asn_itm_1 AND main_stage_0_2);
  or_tmp_2 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_1_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_518_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_2));
  mux_14_nl <= MUX_s_1_2_2(nor_518_nl, or_tmp_2, or_1_cse);
  and_dcpl_300 <= mux_14_nl AND and_dcpl_298 AND and_dcpl_296;
  and_dcpl_301 <= NOT(CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_302 <= and_dcpl_301 AND (NOT (rem_12cyc_st_3_1_0(1)));
  and_dcpl_304 <= (NOT (rem_12cyc_st_3_1_0(0))) AND main_stage_0_4 AND asn_itm_3;
  or_6_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp <= or_6_cse AND or_tmp_2;
  nor_517_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp));
  mux_15_nl <= MUX_s_1_2_2(nor_517_nl, and_tmp, or_1_cse);
  and_dcpl_306 <= mux_15_nl AND and_dcpl_304 AND and_dcpl_302;
  and_dcpl_307 <= NOT(CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_308 <= and_dcpl_307 AND (NOT (rem_12cyc_st_4_1_0(1)));
  and_dcpl_310 <= (NOT (rem_12cyc_st_4_1_0(0))) AND main_stage_0_5 AND asn_itm_4;
  or_10_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_2 <= or_6_cse AND or_10_cse AND or_tmp_2;
  nor_516_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_2));
  mux_16_nl <= MUX_s_1_2_2(nor_516_nl, and_tmp_2, or_1_cse);
  and_dcpl_312 <= mux_16_nl AND and_dcpl_310 AND and_dcpl_308;
  and_dcpl_313 <= NOT(CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_314 <= and_dcpl_313 AND (NOT (rem_12cyc_st_5_1_0(1)));
  and_dcpl_316 <= (NOT (rem_12cyc_st_5_1_0(0))) AND main_stage_0_6 AND asn_itm_5;
  or_15_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_5 <= or_6_cse AND or_10_cse AND or_15_cse AND or_tmp_2;
  nor_515_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_5));
  mux_17_nl <= MUX_s_1_2_2(nor_515_nl, and_tmp_5, or_1_cse);
  and_dcpl_318 <= mux_17_nl AND and_dcpl_316 AND and_dcpl_314;
  or_21_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_9 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND or_tmp_2;
  nor_514_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_9));
  mux_18_nl <= MUX_s_1_2_2(nor_514_nl, and_tmp_9, or_1_cse);
  and_dcpl_324 <= mux_18_nl AND and_dcpl_112 AND and_dcpl_110;
  or_28_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_512_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_2));
  mux_19_nl <= MUX_s_1_2_2(nor_512_nl, or_tmp_2, or_28_cse);
  and_tmp_13 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_19_nl;
  nor_513_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_13));
  mux_20_nl <= MUX_s_1_2_2(nor_513_nl, and_tmp_13, or_1_cse);
  and_dcpl_330 <= mux_20_nl AND and_dcpl_85 AND and_dcpl_83;
  or_37_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_509_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_2));
  mux_tmp_19 <= MUX_s_1_2_2(nor_509_nl, or_tmp_2, or_37_cse);
  nor_510_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_19));
  mux_22_nl <= MUX_s_1_2_2(nor_510_nl, mux_tmp_19, or_28_cse);
  and_tmp_17 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_22_nl;
  nor_511_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_17));
  mux_23_nl <= MUX_s_1_2_2(nor_511_nl, and_tmp_17, or_1_cse);
  and_dcpl_336 <= mux_23_nl AND and_dcpl_58 AND and_dcpl_56;
  or_48_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_505_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_2));
  mux_tmp_22 <= MUX_s_1_2_2(nor_505_nl, or_tmp_2, or_48_cse);
  nor_506_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_22));
  mux_tmp_23 <= MUX_s_1_2_2(nor_506_nl, mux_tmp_22, or_37_cse);
  nor_507_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_23));
  mux_26_nl <= MUX_s_1_2_2(nor_507_nl, mux_tmp_23, or_28_cse);
  and_tmp_21 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_26_nl;
  nor_508_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_21));
  mux_27_nl <= MUX_s_1_2_2(nor_508_nl, and_tmp_21, or_1_cse);
  and_dcpl_342 <= mux_27_nl AND and_dcpl_31 AND and_dcpl_29;
  nor_500_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_2));
  or_61_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_26 <= MUX_s_1_2_2(nor_500_nl, or_tmp_2, or_61_nl);
  nor_501_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_26));
  mux_tmp_27 <= MUX_s_1_2_2(nor_501_nl, mux_tmp_26, or_48_cse);
  nor_502_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_27));
  mux_tmp_28 <= MUX_s_1_2_2(nor_502_nl, mux_tmp_27, or_37_cse);
  nor_503_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_28));
  mux_31_nl <= MUX_s_1_2_2(nor_503_nl, mux_tmp_28, or_28_cse);
  and_tmp_25 <= or_6_cse AND or_10_cse AND or_15_cse AND or_21_cse AND mux_31_nl;
  nor_504_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_25));
  mux_32_nl <= MUX_s_1_2_2(nor_504_nl, and_tmp_25, or_1_cse);
  and_dcpl_348 <= mux_32_nl AND and_dcpl_4 AND and_dcpl_2;
  and_tmp_35 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_8)
      OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND or_6_cse AND
      or_10_cse AND or_15_cse AND or_21_cse AND ((NOT main_stage_0_7) OR (NOT asn_itm_6)
      OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00")))
      AND ((NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_355 <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_356 <= and_dcpl_293 AND and_dcpl_355;
  and_dcpl_358 <= (rem_12cyc_st_2_1_0(0)) AND main_stage_0_3 AND asn_itm_2;
  or_tmp_80 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_83_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_499_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_80));
  mux_33_nl <= MUX_s_1_2_2(nor_499_nl, or_tmp_80, or_83_cse);
  and_dcpl_360 <= mux_33_nl AND and_dcpl_358 AND and_dcpl_296;
  and_dcpl_362 <= (rem_12cyc_st_3_1_0(0)) AND main_stage_0_4 AND asn_itm_3;
  nand_276_cse <= NOT(asn_itm_2 AND main_stage_0_3 AND (rem_12cyc_st_2_1_0(0)));
  or_88_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1168_nl <= nand_276_cse AND or_tmp_80;
  mux_tmp_32 <= MUX_s_1_2_2(and_1168_nl, or_tmp_80, or_88_cse);
  nor_498_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_32));
  mux_35_nl <= MUX_s_1_2_2(nor_498_nl, mux_tmp_32, or_83_cse);
  and_dcpl_364 <= mux_35_nl AND and_dcpl_362 AND and_dcpl_302;
  and_dcpl_366 <= (rem_12cyc_st_4_1_0(0)) AND main_stage_0_5 AND asn_itm_4;
  nand_274_cse <= NOT(asn_itm_3 AND main_stage_0_4 AND (rem_12cyc_st_3_1_0(0)));
  or_93_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1166_nl <= nand_274_cse AND or_tmp_80;
  mux_tmp_34 <= MUX_s_1_2_2(and_1166_nl, or_tmp_80, or_93_cse);
  and_1167_nl <= nand_276_cse AND mux_tmp_34;
  mux_tmp_35 <= MUX_s_1_2_2(and_1167_nl, mux_tmp_34, or_88_cse);
  nor_497_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_35));
  mux_38_nl <= MUX_s_1_2_2(nor_497_nl, mux_tmp_35, or_83_cse);
  and_dcpl_368 <= mux_38_nl AND and_dcpl_366 AND and_dcpl_308;
  and_dcpl_370 <= (rem_12cyc_st_5_1_0(0)) AND main_stage_0_6 AND asn_itm_5;
  nand_271_cse <= NOT(asn_itm_4 AND main_stage_0_5 AND (rem_12cyc_st_4_1_0(0)));
  or_100_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1163_nl <= nand_271_cse AND or_tmp_80;
  mux_tmp_37 <= MUX_s_1_2_2(and_1163_nl, or_tmp_80, or_100_cse);
  and_1164_nl <= nand_274_cse AND mux_tmp_37;
  mux_tmp_38 <= MUX_s_1_2_2(and_1164_nl, mux_tmp_37, or_93_cse);
  and_1165_nl <= nand_276_cse AND mux_tmp_38;
  mux_tmp_39 <= MUX_s_1_2_2(and_1165_nl, mux_tmp_38, or_88_cse);
  nor_496_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_39));
  mux_42_nl <= MUX_s_1_2_2(nor_496_nl, mux_tmp_39, or_83_cse);
  and_dcpl_372 <= mux_42_nl AND and_dcpl_370 AND and_dcpl_314;
  nand_267_cse <= NOT(asn_itm_5 AND main_stage_0_6 AND (rem_12cyc_st_5_1_0(0)));
  or_109_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1159_nl <= nand_267_cse AND or_tmp_80;
  mux_tmp_41 <= MUX_s_1_2_2(and_1159_nl, or_tmp_80, or_109_cse);
  and_1160_nl <= nand_271_cse AND mux_tmp_41;
  mux_tmp_42 <= MUX_s_1_2_2(and_1160_nl, mux_tmp_41, or_100_cse);
  and_1161_nl <= nand_274_cse AND mux_tmp_42;
  mux_tmp_43 <= MUX_s_1_2_2(and_1161_nl, mux_tmp_42, or_93_cse);
  and_1162_nl <= nand_276_cse AND mux_tmp_43;
  mux_tmp_44 <= MUX_s_1_2_2(and_1162_nl, mux_tmp_43, or_88_cse);
  nor_495_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_44));
  mux_47_nl <= MUX_s_1_2_2(nor_495_nl, mux_tmp_44, or_83_cse);
  and_dcpl_376 <= mux_47_nl AND and_dcpl_112 AND and_dcpl_115;
  or_120_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_493_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_80));
  mux_tmp_46 <= MUX_s_1_2_2(nor_493_nl, or_tmp_80, or_120_cse);
  and_1155_nl <= nand_267_cse AND mux_tmp_46;
  mux_tmp_47 <= MUX_s_1_2_2(and_1155_nl, mux_tmp_46, or_109_cse);
  and_1156_nl <= nand_271_cse AND mux_tmp_47;
  mux_tmp_48 <= MUX_s_1_2_2(and_1156_nl, mux_tmp_47, or_100_cse);
  and_1157_nl <= nand_274_cse AND mux_tmp_48;
  mux_tmp_49 <= MUX_s_1_2_2(and_1157_nl, mux_tmp_48, or_93_cse);
  and_1158_nl <= nand_276_cse AND mux_tmp_49;
  mux_tmp_50 <= MUX_s_1_2_2(and_1158_nl, mux_tmp_49, or_88_cse);
  nor_494_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_50));
  mux_53_nl <= MUX_s_1_2_2(nor_494_nl, mux_tmp_50, or_83_cse);
  and_dcpl_379 <= mux_53_nl AND and_dcpl_85 AND and_dcpl_87;
  or_133_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_490_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_80));
  mux_tmp_52 <= MUX_s_1_2_2(nor_490_nl, or_tmp_80, or_133_cse);
  nor_491_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_52));
  mux_tmp_53 <= MUX_s_1_2_2(nor_491_nl, mux_tmp_52, or_120_cse);
  and_1151_nl <= nand_267_cse AND mux_tmp_53;
  mux_tmp_54 <= MUX_s_1_2_2(and_1151_nl, mux_tmp_53, or_109_cse);
  and_1152_nl <= nand_271_cse AND mux_tmp_54;
  mux_tmp_55 <= MUX_s_1_2_2(and_1152_nl, mux_tmp_54, or_100_cse);
  and_1153_nl <= nand_274_cse AND mux_tmp_55;
  mux_tmp_56 <= MUX_s_1_2_2(and_1153_nl, mux_tmp_55, or_93_cse);
  and_1154_nl <= nand_276_cse AND mux_tmp_56;
  mux_tmp_57 <= MUX_s_1_2_2(and_1154_nl, mux_tmp_56, or_88_cse);
  nor_492_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_57));
  mux_60_nl <= MUX_s_1_2_2(nor_492_nl, mux_tmp_57, or_83_cse);
  and_dcpl_382 <= mux_60_nl AND and_dcpl_58 AND and_dcpl_60;
  or_148_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_486_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_80));
  mux_tmp_59 <= MUX_s_1_2_2(nor_486_nl, or_tmp_80, or_148_cse);
  nor_487_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_59));
  mux_tmp_60 <= MUX_s_1_2_2(nor_487_nl, mux_tmp_59, or_133_cse);
  nor_488_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_60));
  mux_tmp_61 <= MUX_s_1_2_2(nor_488_nl, mux_tmp_60, or_120_cse);
  and_1147_nl <= nand_267_cse AND mux_tmp_61;
  mux_tmp_62 <= MUX_s_1_2_2(and_1147_nl, mux_tmp_61, or_109_cse);
  and_1148_nl <= nand_271_cse AND mux_tmp_62;
  mux_tmp_63 <= MUX_s_1_2_2(and_1148_nl, mux_tmp_62, or_100_cse);
  and_1149_nl <= nand_274_cse AND mux_tmp_63;
  mux_tmp_64 <= MUX_s_1_2_2(and_1149_nl, mux_tmp_63, or_93_cse);
  and_1150_nl <= nand_276_cse AND mux_tmp_64;
  mux_tmp_65 <= MUX_s_1_2_2(and_1150_nl, mux_tmp_64, or_88_cse);
  nor_489_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_65));
  mux_68_nl <= MUX_s_1_2_2(nor_489_nl, mux_tmp_65, or_83_cse);
  and_dcpl_385 <= mux_68_nl AND and_dcpl_31 AND and_dcpl_33;
  nor_481_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_80));
  or_165_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_67 <= MUX_s_1_2_2(nor_481_nl, or_tmp_80, or_165_nl);
  nor_482_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_67));
  mux_tmp_68 <= MUX_s_1_2_2(nor_482_nl, mux_tmp_67, or_148_cse);
  nor_483_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_68));
  mux_tmp_69 <= MUX_s_1_2_2(nor_483_nl, mux_tmp_68, or_133_cse);
  nor_484_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_69));
  mux_tmp_70 <= MUX_s_1_2_2(nor_484_nl, mux_tmp_69, or_120_cse);
  and_1143_nl <= nand_267_cse AND mux_tmp_70;
  mux_tmp_71 <= MUX_s_1_2_2(and_1143_nl, mux_tmp_70, or_109_cse);
  and_1144_nl <= nand_271_cse AND mux_tmp_71;
  mux_tmp_72 <= MUX_s_1_2_2(and_1144_nl, mux_tmp_71, or_100_cse);
  and_1145_nl <= nand_274_cse AND mux_tmp_72;
  mux_tmp_73 <= MUX_s_1_2_2(and_1145_nl, mux_tmp_72, or_93_cse);
  and_1146_nl <= nand_276_cse AND mux_tmp_73;
  mux_tmp_74 <= MUX_s_1_2_2(and_1146_nl, mux_tmp_73, or_88_cse);
  nor_485_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_74));
  mux_77_nl <= MUX_s_1_2_2(nor_485_nl, mux_tmp_74, or_83_cse);
  and_dcpl_388 <= mux_77_nl AND and_dcpl_4 AND and_dcpl_6;
  nand_250_cse <= NOT((acc_1_tmp(0)) AND ccs_ccore_start_rsci_idat);
  and_tmp_44 <= ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_3)
      OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_4)
      OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_5)
      OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_6)
      OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_7)
      OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_11)
      OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR (acc_1_tmp(1)) OR nand_250_cse);
  nor_480_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT and_tmp_44));
  or_175_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_76 <= MUX_s_1_2_2(nor_480_nl, and_tmp_44, or_175_nl);
  and_dcpl_393 <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_394 <= and_dcpl_293 AND and_dcpl_393;
  and_dcpl_395 <= and_dcpl_295 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_185 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_190_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_479_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_185));
  mux_79_nl <= MUX_s_1_2_2(nor_479_nl, or_tmp_185, or_190_cse);
  and_dcpl_397 <= mux_79_nl AND and_dcpl_298 AND and_dcpl_395;
  and_dcpl_398 <= and_dcpl_301 AND (rem_12cyc_st_3_1_0(1));
  or_195_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_45 <= or_195_cse AND or_tmp_185;
  nor_478_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_45));
  mux_80_nl <= MUX_s_1_2_2(nor_478_nl, and_tmp_45, or_190_cse);
  and_dcpl_400 <= mux_80_nl AND and_dcpl_304 AND and_dcpl_398;
  and_dcpl_401 <= and_dcpl_307 AND (rem_12cyc_st_4_1_0(1));
  or_199_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_47 <= or_195_cse AND or_199_cse AND or_tmp_185;
  nor_477_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_47));
  mux_81_nl <= MUX_s_1_2_2(nor_477_nl, and_tmp_47, or_190_cse);
  and_dcpl_403 <= mux_81_nl AND and_dcpl_310 AND and_dcpl_401;
  and_dcpl_404 <= and_dcpl_313 AND (rem_12cyc_st_5_1_0(1));
  or_204_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_50 <= or_195_cse AND or_199_cse AND or_204_cse AND or_tmp_185;
  nor_476_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_50));
  mux_82_nl <= MUX_s_1_2_2(nor_476_nl, and_tmp_50, or_190_cse);
  and_dcpl_406 <= mux_82_nl AND and_dcpl_316 AND and_dcpl_404;
  or_210_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_54 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND or_tmp_185;
  nor_475_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_54));
  mux_83_nl <= MUX_s_1_2_2(nor_475_nl, and_tmp_54, or_190_cse);
  and_dcpl_409 <= mux_83_nl AND and_dcpl_112 AND and_dcpl_117;
  or_217_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_473_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_185));
  mux_84_nl <= MUX_s_1_2_2(nor_473_nl, or_tmp_185, or_217_cse);
  and_tmp_58 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_84_nl;
  nor_474_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_58));
  mux_85_nl <= MUX_s_1_2_2(nor_474_nl, and_tmp_58, or_190_cse);
  and_dcpl_413 <= mux_85_nl AND and_dcpl_85 AND and_dcpl_90;
  or_226_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_470_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_185));
  mux_tmp_84 <= MUX_s_1_2_2(nor_470_nl, or_tmp_185, or_226_cse);
  nor_471_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_84));
  mux_87_nl <= MUX_s_1_2_2(nor_471_nl, mux_tmp_84, or_217_cse);
  and_tmp_62 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_87_nl;
  nor_472_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_62));
  mux_88_nl <= MUX_s_1_2_2(nor_472_nl, and_tmp_62, or_190_cse);
  and_dcpl_417 <= mux_88_nl AND and_dcpl_58 AND and_dcpl_63;
  or_237_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_466_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_185));
  mux_tmp_87 <= MUX_s_1_2_2(nor_466_nl, or_tmp_185, or_237_cse);
  nor_467_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_87));
  mux_tmp_88 <= MUX_s_1_2_2(nor_467_nl, mux_tmp_87, or_226_cse);
  nor_468_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_88));
  mux_91_nl <= MUX_s_1_2_2(nor_468_nl, mux_tmp_88, or_217_cse);
  and_tmp_66 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_91_nl;
  nor_469_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_66));
  mux_92_nl <= MUX_s_1_2_2(nor_469_nl, and_tmp_66, or_190_cse);
  and_dcpl_421 <= mux_92_nl AND and_dcpl_31 AND and_dcpl_36;
  nor_461_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_185));
  or_250_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_91 <= MUX_s_1_2_2(nor_461_nl, or_tmp_185, or_250_nl);
  nor_462_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_91));
  mux_tmp_92 <= MUX_s_1_2_2(nor_462_nl, mux_tmp_91, or_237_cse);
  nor_463_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_92));
  mux_tmp_93 <= MUX_s_1_2_2(nor_463_nl, mux_tmp_92, or_226_cse);
  nor_464_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_93));
  mux_96_nl <= MUX_s_1_2_2(nor_464_nl, mux_tmp_93, or_217_cse);
  and_tmp_70 <= or_195_cse AND or_199_cse AND or_204_cse AND or_210_cse AND mux_96_nl;
  nor_465_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_70));
  mux_97_nl <= MUX_s_1_2_2(nor_465_nl, and_tmp_70, or_190_cse);
  and_dcpl_425 <= mux_97_nl AND and_dcpl_4 AND and_dcpl_9;
  and_tmp_80 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND ((NOT main_stage_0_8)
      OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND or_195_cse
      AND or_199_cse AND or_204_cse AND or_210_cse AND ((NOT main_stage_0_7) OR (NOT
      asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00")))
      AND ((NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_430 <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_431 <= and_dcpl_293 AND and_dcpl_430;
  or_tmp_263 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_54;
  or_270_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"));
  nor_460_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_263));
  mux_98_nl <= MUX_s_1_2_2(nor_460_nl, or_tmp_263, or_270_cse);
  and_dcpl_433 <= mux_98_nl AND and_dcpl_358 AND and_dcpl_395;
  or_275_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1142_nl <= nand_276_cse AND or_tmp_263;
  mux_tmp_97 <= MUX_s_1_2_2(and_1142_nl, or_tmp_263, or_275_cse);
  nor_459_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_97));
  mux_100_nl <= MUX_s_1_2_2(nor_459_nl, mux_tmp_97, or_270_cse);
  and_dcpl_435 <= mux_100_nl AND and_dcpl_362 AND and_dcpl_398;
  or_280_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1140_nl <= nand_274_cse AND or_tmp_263;
  mux_tmp_99 <= MUX_s_1_2_2(and_1140_nl, or_tmp_263, or_280_cse);
  and_1141_nl <= nand_276_cse AND mux_tmp_99;
  mux_tmp_100 <= MUX_s_1_2_2(and_1141_nl, mux_tmp_99, or_275_cse);
  nor_458_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_100));
  mux_103_nl <= MUX_s_1_2_2(nor_458_nl, mux_tmp_100, or_270_cse);
  and_dcpl_437 <= mux_103_nl AND and_dcpl_366 AND and_dcpl_401;
  or_287_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1137_nl <= nand_271_cse AND or_tmp_263;
  mux_tmp_102 <= MUX_s_1_2_2(and_1137_nl, or_tmp_263, or_287_cse);
  and_1138_nl <= nand_274_cse AND mux_tmp_102;
  mux_tmp_103 <= MUX_s_1_2_2(and_1138_nl, mux_tmp_102, or_280_cse);
  and_1139_nl <= nand_276_cse AND mux_tmp_103;
  mux_tmp_104 <= MUX_s_1_2_2(and_1139_nl, mux_tmp_103, or_275_cse);
  nor_457_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_104));
  mux_107_nl <= MUX_s_1_2_2(nor_457_nl, mux_tmp_104, or_270_cse);
  and_dcpl_439 <= mux_107_nl AND and_dcpl_370 AND and_dcpl_404;
  or_296_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"));
  and_1133_nl <= nand_267_cse AND or_tmp_263;
  mux_tmp_106 <= MUX_s_1_2_2(and_1133_nl, or_tmp_263, or_296_cse);
  and_1134_nl <= nand_271_cse AND mux_tmp_106;
  mux_tmp_107 <= MUX_s_1_2_2(and_1134_nl, mux_tmp_106, or_287_cse);
  and_1135_nl <= nand_274_cse AND mux_tmp_107;
  mux_tmp_108 <= MUX_s_1_2_2(and_1135_nl, mux_tmp_107, or_280_cse);
  and_1136_nl <= nand_276_cse AND mux_tmp_108;
  mux_tmp_109 <= MUX_s_1_2_2(and_1136_nl, mux_tmp_108, or_275_cse);
  nor_456_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_109));
  mux_112_nl <= MUX_s_1_2_2(nor_456_nl, mux_tmp_109, or_270_cse);
  and_dcpl_442 <= mux_112_nl AND and_dcpl_112 AND and_dcpl_119;
  or_307_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_454_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_263));
  mux_tmp_111 <= MUX_s_1_2_2(nor_454_nl, or_tmp_263, or_307_cse);
  and_1129_nl <= nand_267_cse AND mux_tmp_111;
  mux_tmp_112 <= MUX_s_1_2_2(and_1129_nl, mux_tmp_111, or_296_cse);
  and_1130_nl <= nand_271_cse AND mux_tmp_112;
  mux_tmp_113 <= MUX_s_1_2_2(and_1130_nl, mux_tmp_112, or_287_cse);
  and_1131_nl <= nand_274_cse AND mux_tmp_113;
  mux_tmp_114 <= MUX_s_1_2_2(and_1131_nl, mux_tmp_113, or_280_cse);
  and_1132_nl <= nand_276_cse AND mux_tmp_114;
  mux_tmp_115 <= MUX_s_1_2_2(and_1132_nl, mux_tmp_114, or_275_cse);
  nor_455_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_115));
  mux_118_nl <= MUX_s_1_2_2(nor_455_nl, mux_tmp_115, or_270_cse);
  and_dcpl_445 <= mux_118_nl AND and_dcpl_85 AND and_dcpl_92;
  or_320_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_451_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_263));
  mux_tmp_117 <= MUX_s_1_2_2(nor_451_nl, or_tmp_263, or_320_cse);
  nor_452_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_117));
  mux_tmp_118 <= MUX_s_1_2_2(nor_452_nl, mux_tmp_117, or_307_cse);
  and_1125_nl <= nand_267_cse AND mux_tmp_118;
  mux_tmp_119 <= MUX_s_1_2_2(and_1125_nl, mux_tmp_118, or_296_cse);
  and_1126_nl <= nand_271_cse AND mux_tmp_119;
  mux_tmp_120 <= MUX_s_1_2_2(and_1126_nl, mux_tmp_119, or_287_cse);
  and_1127_nl <= nand_274_cse AND mux_tmp_120;
  mux_tmp_121 <= MUX_s_1_2_2(and_1127_nl, mux_tmp_120, or_280_cse);
  and_1128_nl <= nand_276_cse AND mux_tmp_121;
  mux_tmp_122 <= MUX_s_1_2_2(and_1128_nl, mux_tmp_121, or_275_cse);
  nor_453_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_122));
  mux_125_nl <= MUX_s_1_2_2(nor_453_nl, mux_tmp_122, or_270_cse);
  and_dcpl_448 <= mux_125_nl AND and_dcpl_58 AND and_dcpl_65;
  or_335_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"));
  nor_447_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_263));
  mux_tmp_124 <= MUX_s_1_2_2(nor_447_nl, or_tmp_263, or_335_cse);
  nor_448_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_124));
  mux_tmp_125 <= MUX_s_1_2_2(nor_448_nl, mux_tmp_124, or_320_cse);
  nor_449_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_125));
  mux_tmp_126 <= MUX_s_1_2_2(nor_449_nl, mux_tmp_125, or_307_cse);
  and_1121_nl <= nand_267_cse AND mux_tmp_126;
  mux_tmp_127 <= MUX_s_1_2_2(and_1121_nl, mux_tmp_126, or_296_cse);
  and_1122_nl <= nand_271_cse AND mux_tmp_127;
  mux_tmp_128 <= MUX_s_1_2_2(and_1122_nl, mux_tmp_127, or_287_cse);
  and_1123_nl <= nand_274_cse AND mux_tmp_128;
  mux_tmp_129 <= MUX_s_1_2_2(and_1123_nl, mux_tmp_128, or_280_cse);
  and_1124_nl <= nand_276_cse AND mux_tmp_129;
  mux_tmp_130 <= MUX_s_1_2_2(and_1124_nl, mux_tmp_129, or_275_cse);
  nor_450_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_130));
  mux_133_nl <= MUX_s_1_2_2(nor_450_nl, mux_tmp_130, or_270_cse);
  and_dcpl_451 <= mux_133_nl AND and_dcpl_31 AND and_dcpl_38;
  nor_442_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_263));
  or_352_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_132 <= MUX_s_1_2_2(nor_442_nl, or_tmp_263, or_352_nl);
  nor_443_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_132));
  mux_tmp_133 <= MUX_s_1_2_2(nor_443_nl, mux_tmp_132, or_335_cse);
  nor_444_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_133));
  mux_tmp_134 <= MUX_s_1_2_2(nor_444_nl, mux_tmp_133, or_320_cse);
  nor_445_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_134));
  mux_tmp_135 <= MUX_s_1_2_2(nor_445_nl, mux_tmp_134, or_307_cse);
  and_1117_nl <= nand_267_cse AND mux_tmp_135;
  mux_tmp_136 <= MUX_s_1_2_2(and_1117_nl, mux_tmp_135, or_296_cse);
  and_1118_nl <= nand_271_cse AND mux_tmp_136;
  mux_tmp_137 <= MUX_s_1_2_2(and_1118_nl, mux_tmp_136, or_287_cse);
  and_1119_nl <= nand_274_cse AND mux_tmp_137;
  mux_tmp_138 <= MUX_s_1_2_2(and_1119_nl, mux_tmp_137, or_280_cse);
  and_1120_nl <= nand_276_cse AND mux_tmp_138;
  mux_tmp_139 <= MUX_s_1_2_2(and_1120_nl, mux_tmp_138, or_275_cse);
  nor_446_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_139));
  mux_142_nl <= MUX_s_1_2_2(nor_446_nl, mux_tmp_139, or_270_cse);
  and_dcpl_454 <= mux_142_nl AND and_dcpl_4 AND and_dcpl_11;
  nand_222_cse <= NOT(CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND ccs_ccore_start_rsci_idat);
  and_tmp_89 <= ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_3)
      OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_4)
      OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_5)
      OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_6)
      OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_7)
      OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_11)
      OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("00"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("00"))
      OR nand_222_cse);
  nand_223_cse <= NOT(CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11")));
  and_1116_nl <= nand_223_cse AND and_tmp_89;
  or_362_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_141 <= MUX_s_1_2_2(and_1116_nl, and_tmp_89, or_362_nl);
  and_dcpl_460 <= ccs_ccore_start_rsci_idat AND CONV_SL_1_1(acc_tmp=STD_LOGIC_VECTOR'("01"));
  and_dcpl_461 <= and_dcpl_460 AND and_dcpl_291;
  and_dcpl_462 <= CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_463 <= and_dcpl_462 AND (NOT (rem_12cyc_st_2_1_0(1)));
  not_tmp_332 <= NOT((rem_12cyc_3_2(0)) AND asn_itm_1 AND main_stage_0_2);
  or_tmp_368 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  nand_281_cse <= NOT((acc_tmp(0)) AND ccs_ccore_start_rsci_idat);
  or_377_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (acc_tmp(1));
  and_1172_nl <= nand_281_cse AND or_tmp_368;
  mux_144_nl <= MUX_s_1_2_2(and_1172_nl, or_tmp_368, or_377_cse);
  and_dcpl_465 <= mux_144_nl AND and_dcpl_298 AND and_dcpl_463;
  and_dcpl_466 <= CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_467 <= and_dcpl_466 AND (NOT (rem_12cyc_st_3_1_0(1)));
  or_382_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_90 <= or_382_cse AND or_tmp_368;
  and_1114_nl <= nand_281_cse AND and_tmp_90;
  mux_145_nl <= MUX_s_1_2_2(and_1114_nl, and_tmp_90, or_377_cse);
  and_dcpl_469 <= mux_145_nl AND and_dcpl_304 AND and_dcpl_467;
  and_dcpl_470 <= CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_471 <= and_dcpl_470 AND (NOT (rem_12cyc_st_4_1_0(1)));
  or_386_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_92 <= or_382_cse AND or_386_cse AND or_tmp_368;
  and_1113_nl <= nand_281_cse AND and_tmp_92;
  mux_146_nl <= MUX_s_1_2_2(and_1113_nl, and_tmp_92, or_377_cse);
  and_dcpl_473 <= mux_146_nl AND and_dcpl_310 AND and_dcpl_471;
  and_dcpl_474 <= CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("01"));
  and_dcpl_475 <= and_dcpl_474 AND (NOT (rem_12cyc_st_5_1_0(1)));
  or_391_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_95 <= or_382_cse AND or_386_cse AND or_391_cse AND or_tmp_368;
  and_1112_nl <= nand_281_cse AND and_tmp_95;
  mux_147_nl <= MUX_s_1_2_2(and_1112_nl, and_tmp_95, or_377_cse);
  and_dcpl_477 <= mux_147_nl AND and_dcpl_316 AND and_dcpl_475;
  or_397_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_99 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND or_tmp_368;
  and_1111_nl <= nand_281_cse AND and_tmp_99;
  mux_148_nl <= MUX_s_1_2_2(and_1111_nl, and_tmp_99, or_377_cse);
  and_dcpl_480 <= mux_148_nl AND and_dcpl_121 AND and_dcpl_110;
  nand_215_cse <= NOT((rem_12cyc_st_6_3_2(0)) AND asn_itm_6 AND main_stage_0_7);
  or_404_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_6_3_2(1));
  and_1109_nl <= nand_215_cse AND or_tmp_368;
  mux_149_nl <= MUX_s_1_2_2(and_1109_nl, or_tmp_368, or_404_cse);
  and_tmp_103 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_149_nl;
  and_1110_nl <= nand_281_cse AND and_tmp_103;
  mux_150_nl <= MUX_s_1_2_2(and_1110_nl, and_tmp_103, or_377_cse);
  and_dcpl_483 <= mux_150_nl AND and_dcpl_94 AND and_dcpl_83;
  nand_212_cse <= NOT((rem_12cyc_st_7_3_2(0)) AND asn_itm_7 AND main_stage_0_8);
  or_413_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_7_3_2(1));
  and_1106_nl <= nand_212_cse AND or_tmp_368;
  mux_tmp_149 <= MUX_s_1_2_2(and_1106_nl, or_tmp_368, or_413_cse);
  and_1107_nl <= nand_215_cse AND mux_tmp_149;
  mux_152_nl <= MUX_s_1_2_2(and_1107_nl, mux_tmp_149, or_404_cse);
  and_tmp_107 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_152_nl;
  and_1108_nl <= nand_281_cse AND and_tmp_107;
  mux_153_nl <= MUX_s_1_2_2(and_1108_nl, and_tmp_107, or_377_cse);
  and_dcpl_486 <= mux_153_nl AND and_dcpl_67 AND and_dcpl_56;
  nand_208_cse <= NOT((rem_12cyc_st_8_3_2(0)) AND asn_itm_8 AND main_stage_0_9);
  or_424_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_8_3_2(1));
  and_1102_nl <= nand_208_cse AND or_tmp_368;
  mux_tmp_152 <= MUX_s_1_2_2(and_1102_nl, or_tmp_368, or_424_cse);
  and_1103_nl <= nand_212_cse AND mux_tmp_152;
  mux_tmp_153 <= MUX_s_1_2_2(and_1103_nl, mux_tmp_152, or_413_cse);
  and_1104_nl <= nand_215_cse AND mux_tmp_153;
  mux_156_nl <= MUX_s_1_2_2(and_1104_nl, mux_tmp_153, or_404_cse);
  and_tmp_111 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_156_nl;
  and_1105_nl <= nand_281_cse AND and_tmp_111;
  mux_157_nl <= MUX_s_1_2_2(and_1105_nl, and_tmp_111, or_377_cse);
  and_dcpl_489 <= mux_157_nl AND and_dcpl_40 AND and_dcpl_29;
  nand_203_cse <= NOT((rem_12cyc_st_9_3_2(0)) AND asn_itm_9 AND main_stage_0_10);
  and_1097_nl <= nand_203_cse AND or_tmp_368;
  or_437_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_156 <= MUX_s_1_2_2(and_1097_nl, or_tmp_368, or_437_nl);
  and_1098_nl <= nand_208_cse AND mux_tmp_156;
  mux_tmp_157 <= MUX_s_1_2_2(and_1098_nl, mux_tmp_156, or_424_cse);
  and_1099_nl <= nand_212_cse AND mux_tmp_157;
  mux_tmp_158 <= MUX_s_1_2_2(and_1099_nl, mux_tmp_157, or_413_cse);
  and_1100_nl <= nand_215_cse AND mux_tmp_158;
  mux_161_nl <= MUX_s_1_2_2(and_1100_nl, mux_tmp_158, or_404_cse);
  and_tmp_115 <= or_382_cse AND or_386_cse AND or_391_cse AND or_397_cse AND mux_161_nl;
  and_1101_nl <= nand_281_cse AND and_tmp_115;
  mux_162_nl <= MUX_s_1_2_2(and_1101_nl, and_tmp_115, or_377_cse);
  and_dcpl_492 <= mux_162_nl AND and_dcpl_13 AND and_dcpl_2;
  and_tmp_125 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND ((NOT main_stage_0_8)
      OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND or_382_cse
      AND or_386_cse AND or_391_cse AND or_397_cse AND ((NOT main_stage_0_7) OR (NOT
      asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01")))
      AND ((NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_498 <= and_dcpl_460 AND and_dcpl_355;
  or_tmp_446 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_458_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR (acc_tmp(1));
  and_1171_nl <= nand_281_cse AND or_tmp_446;
  mux_163_nl <= MUX_s_1_2_2(and_1171_nl, or_tmp_446, or_458_cse);
  and_dcpl_500 <= mux_163_nl AND and_dcpl_358 AND and_dcpl_463;
  or_463_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1094_nl <= nand_276_cse AND or_tmp_446;
  mux_tmp_162 <= MUX_s_1_2_2(and_1094_nl, or_tmp_446, or_463_cse);
  and_1095_nl <= nand_281_cse AND mux_tmp_162;
  mux_165_nl <= MUX_s_1_2_2(and_1095_nl, mux_tmp_162, or_458_cse);
  and_dcpl_502 <= mux_165_nl AND and_dcpl_362 AND and_dcpl_467;
  nand_198_cse <= NOT((rem_12cyc_st_3_3_2(0)) AND asn_itm_3 AND main_stage_0_4 AND
      (rem_12cyc_st_3_1_0(0)));
  or_468_cse <= (rem_12cyc_st_3_1_0(1)) OR (rem_12cyc_st_3_3_2(1));
  and_1091_nl <= nand_198_cse AND or_tmp_446;
  mux_tmp_164 <= MUX_s_1_2_2(and_1091_nl, or_tmp_446, or_468_cse);
  and_1092_nl <= nand_276_cse AND mux_tmp_164;
  mux_tmp_165 <= MUX_s_1_2_2(and_1092_nl, mux_tmp_164, or_463_cse);
  and_1093_nl <= nand_281_cse AND mux_tmp_165;
  mux_168_nl <= MUX_s_1_2_2(and_1093_nl, mux_tmp_165, or_458_cse);
  and_dcpl_504 <= mux_168_nl AND and_dcpl_366 AND and_dcpl_471;
  or_475_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1087_nl <= nand_271_cse AND or_tmp_446;
  mux_tmp_167 <= MUX_s_1_2_2(and_1087_nl, or_tmp_446, or_475_cse);
  and_1088_nl <= nand_198_cse AND mux_tmp_167;
  mux_tmp_168 <= MUX_s_1_2_2(and_1088_nl, mux_tmp_167, or_468_cse);
  and_1089_nl <= nand_276_cse AND mux_tmp_168;
  mux_tmp_169 <= MUX_s_1_2_2(and_1089_nl, mux_tmp_168, or_463_cse);
  and_1090_nl <= nand_281_cse AND mux_tmp_169;
  mux_172_nl <= MUX_s_1_2_2(and_1090_nl, mux_tmp_169, or_458_cse);
  and_dcpl_506 <= mux_172_nl AND and_dcpl_370 AND and_dcpl_475;
  nand_189_cse <= NOT((rem_12cyc_st_5_3_2(0)) AND asn_itm_5 AND main_stage_0_6 AND
      (rem_12cyc_st_5_1_0(0)));
  or_484_cse <= (rem_12cyc_st_5_1_0(1)) OR (rem_12cyc_st_5_3_2(1));
  and_1082_nl <= nand_189_cse AND or_tmp_446;
  mux_tmp_171 <= MUX_s_1_2_2(and_1082_nl, or_tmp_446, or_484_cse);
  and_1083_nl <= nand_271_cse AND mux_tmp_171;
  mux_tmp_172 <= MUX_s_1_2_2(and_1083_nl, mux_tmp_171, or_475_cse);
  and_1084_nl <= nand_198_cse AND mux_tmp_172;
  mux_tmp_173 <= MUX_s_1_2_2(and_1084_nl, mux_tmp_172, or_468_cse);
  and_1085_nl <= nand_276_cse AND mux_tmp_173;
  mux_tmp_174 <= MUX_s_1_2_2(and_1085_nl, mux_tmp_173, or_463_cse);
  and_1086_nl <= nand_281_cse AND mux_tmp_174;
  mux_177_nl <= MUX_s_1_2_2(and_1086_nl, mux_tmp_174, or_458_cse);
  and_dcpl_508 <= mux_177_nl AND and_dcpl_121 AND and_dcpl_115;
  or_495_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_6_3_2(1));
  and_1076_nl <= nand_215_cse AND or_tmp_446;
  mux_tmp_176 <= MUX_s_1_2_2(and_1076_nl, or_tmp_446, or_495_cse);
  and_1077_nl <= nand_189_cse AND mux_tmp_176;
  mux_tmp_177 <= MUX_s_1_2_2(and_1077_nl, mux_tmp_176, or_484_cse);
  and_1078_nl <= nand_271_cse AND mux_tmp_177;
  mux_tmp_178 <= MUX_s_1_2_2(and_1078_nl, mux_tmp_177, or_475_cse);
  and_1079_nl <= nand_198_cse AND mux_tmp_178;
  mux_tmp_179 <= MUX_s_1_2_2(and_1079_nl, mux_tmp_178, or_468_cse);
  and_1080_nl <= nand_276_cse AND mux_tmp_179;
  mux_tmp_180 <= MUX_s_1_2_2(and_1080_nl, mux_tmp_179, or_463_cse);
  and_1081_nl <= nand_281_cse AND mux_tmp_180;
  mux_183_nl <= MUX_s_1_2_2(and_1081_nl, mux_tmp_180, or_458_cse);
  and_dcpl_510 <= mux_183_nl AND and_dcpl_94 AND and_dcpl_87;
  or_508_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_7_3_2(1));
  and_1069_nl <= nand_212_cse AND or_tmp_446;
  mux_tmp_182 <= MUX_s_1_2_2(and_1069_nl, or_tmp_446, or_508_cse);
  and_1070_nl <= nand_215_cse AND mux_tmp_182;
  mux_tmp_183 <= MUX_s_1_2_2(and_1070_nl, mux_tmp_182, or_495_cse);
  and_1071_nl <= nand_189_cse AND mux_tmp_183;
  mux_tmp_184 <= MUX_s_1_2_2(and_1071_nl, mux_tmp_183, or_484_cse);
  and_1072_nl <= nand_271_cse AND mux_tmp_184;
  mux_tmp_185 <= MUX_s_1_2_2(and_1072_nl, mux_tmp_184, or_475_cse);
  and_1073_nl <= nand_198_cse AND mux_tmp_185;
  mux_tmp_186 <= MUX_s_1_2_2(and_1073_nl, mux_tmp_185, or_468_cse);
  and_1074_nl <= nand_276_cse AND mux_tmp_186;
  mux_tmp_187 <= MUX_s_1_2_2(and_1074_nl, mux_tmp_186, or_463_cse);
  and_1075_nl <= nand_281_cse AND mux_tmp_187;
  mux_190_nl <= MUX_s_1_2_2(and_1075_nl, mux_tmp_187, or_458_cse);
  and_dcpl_512 <= mux_190_nl AND and_dcpl_67 AND and_dcpl_60;
  or_523_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_8_3_2(1));
  and_1061_nl <= nand_208_cse AND or_tmp_446;
  mux_tmp_189 <= MUX_s_1_2_2(and_1061_nl, or_tmp_446, or_523_cse);
  and_1062_nl <= nand_212_cse AND mux_tmp_189;
  mux_tmp_190 <= MUX_s_1_2_2(and_1062_nl, mux_tmp_189, or_508_cse);
  and_1063_nl <= nand_215_cse AND mux_tmp_190;
  mux_tmp_191 <= MUX_s_1_2_2(and_1063_nl, mux_tmp_190, or_495_cse);
  and_1064_nl <= nand_189_cse AND mux_tmp_191;
  mux_tmp_192 <= MUX_s_1_2_2(and_1064_nl, mux_tmp_191, or_484_cse);
  and_1065_nl <= nand_271_cse AND mux_tmp_192;
  mux_tmp_193 <= MUX_s_1_2_2(and_1065_nl, mux_tmp_192, or_475_cse);
  and_1066_nl <= nand_198_cse AND mux_tmp_193;
  mux_tmp_194 <= MUX_s_1_2_2(and_1066_nl, mux_tmp_193, or_468_cse);
  and_1067_nl <= nand_276_cse AND mux_tmp_194;
  mux_tmp_195 <= MUX_s_1_2_2(and_1067_nl, mux_tmp_194, or_463_cse);
  and_1068_nl <= nand_281_cse AND mux_tmp_195;
  mux_198_nl <= MUX_s_1_2_2(and_1068_nl, mux_tmp_195, or_458_cse);
  and_dcpl_514 <= mux_198_nl AND and_dcpl_40 AND and_dcpl_33;
  and_1052_nl <= nand_203_cse AND or_tmp_446;
  or_540_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_197 <= MUX_s_1_2_2(and_1052_nl, or_tmp_446, or_540_nl);
  and_1053_nl <= nand_208_cse AND mux_tmp_197;
  mux_tmp_198 <= MUX_s_1_2_2(and_1053_nl, mux_tmp_197, or_523_cse);
  and_1054_nl <= nand_212_cse AND mux_tmp_198;
  mux_tmp_199 <= MUX_s_1_2_2(and_1054_nl, mux_tmp_198, or_508_cse);
  and_1055_nl <= nand_215_cse AND mux_tmp_199;
  mux_tmp_200 <= MUX_s_1_2_2(and_1055_nl, mux_tmp_199, or_495_cse);
  and_1056_nl <= nand_189_cse AND mux_tmp_200;
  mux_tmp_201 <= MUX_s_1_2_2(and_1056_nl, mux_tmp_200, or_484_cse);
  and_1057_nl <= nand_271_cse AND mux_tmp_201;
  mux_tmp_202 <= MUX_s_1_2_2(and_1057_nl, mux_tmp_201, or_475_cse);
  and_1058_nl <= nand_198_cse AND mux_tmp_202;
  mux_tmp_203 <= MUX_s_1_2_2(and_1058_nl, mux_tmp_202, or_468_cse);
  and_1059_nl <= nand_276_cse AND mux_tmp_203;
  mux_tmp_204 <= MUX_s_1_2_2(and_1059_nl, mux_tmp_203, or_463_cse);
  and_1060_nl <= nand_281_cse AND mux_tmp_204;
  mux_207_nl <= MUX_s_1_2_2(and_1060_nl, mux_tmp_204, or_458_cse);
  and_dcpl_516 <= mux_207_nl AND and_dcpl_13 AND and_dcpl_6;
  and_tmp_134 <= ((NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_3)
      OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_4)
      OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_5)
      OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_6)
      OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_7)
      OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_11)
      OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR (acc_1_tmp(1)) OR nand_250_cse);
  nor_439_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT and_tmp_134));
  or_550_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_206 <= MUX_s_1_2_2(nor_439_nl, and_tmp_134, or_550_nl);
  and_dcpl_520 <= and_dcpl_460 AND and_dcpl_393;
  and_dcpl_521 <= and_dcpl_462 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_551 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_564_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (acc_tmp(1));
  and_1170_nl <= nand_281_cse AND or_tmp_551;
  mux_209_nl <= MUX_s_1_2_2(and_1170_nl, or_tmp_551, or_564_cse);
  and_dcpl_523 <= mux_209_nl AND and_dcpl_298 AND and_dcpl_521;
  and_dcpl_524 <= and_dcpl_466 AND (rem_12cyc_st_3_1_0(1));
  or_569_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_135 <= or_569_cse AND or_tmp_551;
  and_1050_nl <= nand_281_cse AND and_tmp_135;
  mux_210_nl <= MUX_s_1_2_2(and_1050_nl, and_tmp_135, or_564_cse);
  and_dcpl_526 <= mux_210_nl AND and_dcpl_304 AND and_dcpl_524;
  and_dcpl_527 <= and_dcpl_470 AND (rem_12cyc_st_4_1_0(1));
  or_573_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_137 <= or_569_cse AND or_573_cse AND or_tmp_551;
  and_1049_nl <= nand_281_cse AND and_tmp_137;
  mux_211_nl <= MUX_s_1_2_2(and_1049_nl, and_tmp_137, or_564_cse);
  and_dcpl_529 <= mux_211_nl AND and_dcpl_310 AND and_dcpl_527;
  and_dcpl_530 <= and_dcpl_474 AND (rem_12cyc_st_5_1_0(1));
  or_578_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_140 <= or_569_cse AND or_573_cse AND or_578_cse AND or_tmp_551;
  and_1048_nl <= nand_281_cse AND and_tmp_140;
  mux_212_nl <= MUX_s_1_2_2(and_1048_nl, and_tmp_140, or_564_cse);
  and_dcpl_532 <= mux_212_nl AND and_dcpl_316 AND and_dcpl_530;
  or_584_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("01"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_144 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND or_tmp_551;
  and_1047_nl <= nand_281_cse AND and_tmp_144;
  mux_213_nl <= MUX_s_1_2_2(and_1047_nl, and_tmp_144, or_564_cse);
  and_dcpl_534 <= mux_213_nl AND and_dcpl_121 AND and_dcpl_117;
  or_591_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_6_3_2(1));
  and_1045_nl <= nand_215_cse AND or_tmp_551;
  mux_214_nl <= MUX_s_1_2_2(and_1045_nl, or_tmp_551, or_591_cse);
  and_tmp_148 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_214_nl;
  and_1046_nl <= nand_281_cse AND and_tmp_148;
  mux_215_nl <= MUX_s_1_2_2(and_1046_nl, and_tmp_148, or_564_cse);
  and_dcpl_536 <= mux_215_nl AND and_dcpl_94 AND and_dcpl_90;
  or_600_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_7_3_2(1));
  and_1042_nl <= nand_212_cse AND or_tmp_551;
  mux_tmp_214 <= MUX_s_1_2_2(and_1042_nl, or_tmp_551, or_600_cse);
  and_1043_nl <= nand_215_cse AND mux_tmp_214;
  mux_217_nl <= MUX_s_1_2_2(and_1043_nl, mux_tmp_214, or_591_cse);
  and_tmp_152 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_217_nl;
  and_1044_nl <= nand_281_cse AND and_tmp_152;
  mux_218_nl <= MUX_s_1_2_2(and_1044_nl, and_tmp_152, or_564_cse);
  and_dcpl_538 <= mux_218_nl AND and_dcpl_67 AND and_dcpl_63;
  or_611_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_8_3_2(1));
  and_1038_nl <= nand_208_cse AND or_tmp_551;
  mux_tmp_217 <= MUX_s_1_2_2(and_1038_nl, or_tmp_551, or_611_cse);
  and_1039_nl <= nand_212_cse AND mux_tmp_217;
  mux_tmp_218 <= MUX_s_1_2_2(and_1039_nl, mux_tmp_217, or_600_cse);
  and_1040_nl <= nand_215_cse AND mux_tmp_218;
  mux_221_nl <= MUX_s_1_2_2(and_1040_nl, mux_tmp_218, or_591_cse);
  and_tmp_156 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_221_nl;
  and_1041_nl <= nand_281_cse AND and_tmp_156;
  mux_222_nl <= MUX_s_1_2_2(and_1041_nl, and_tmp_156, or_564_cse);
  and_dcpl_540 <= mux_222_nl AND and_dcpl_40 AND and_dcpl_36;
  and_1033_nl <= nand_203_cse AND or_tmp_551;
  or_624_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_221 <= MUX_s_1_2_2(and_1033_nl, or_tmp_551, or_624_nl);
  and_1034_nl <= nand_208_cse AND mux_tmp_221;
  mux_tmp_222 <= MUX_s_1_2_2(and_1034_nl, mux_tmp_221, or_611_cse);
  and_1035_nl <= nand_212_cse AND mux_tmp_222;
  mux_tmp_223 <= MUX_s_1_2_2(and_1035_nl, mux_tmp_222, or_600_cse);
  and_1036_nl <= nand_215_cse AND mux_tmp_223;
  mux_226_nl <= MUX_s_1_2_2(and_1036_nl, mux_tmp_223, or_591_cse);
  and_tmp_160 <= or_569_cse AND or_573_cse AND or_578_cse AND or_584_cse AND mux_226_nl;
  and_1037_nl <= nand_281_cse AND and_tmp_160;
  mux_227_nl <= MUX_s_1_2_2(and_1037_nl, and_tmp_160, or_564_cse);
  and_dcpl_542 <= mux_227_nl AND and_dcpl_13 AND and_dcpl_9;
  and_tmp_170 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND ((NOT main_stage_0_8)
      OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_9)
      OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("01"))) AND ((NOT main_stage_0_10)
      OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("01"))) AND or_569_cse
      AND or_573_cse AND or_578_cse AND or_584_cse AND ((NOT main_stage_0_7) OR (NOT
      asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("01")))
      AND ((NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_st_10_3_2/=STD_LOGIC_VECTOR'("01"))) AND (CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT ccs_ccore_start_rsci_idat));
  and_dcpl_546 <= and_dcpl_460 AND and_dcpl_430;
  or_tmp_629 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_3_2(1))
      OR not_tmp_332;
  or_643_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (acc_tmp(1));
  and_1169_nl <= nand_281_cse AND or_tmp_629;
  mux_228_nl <= MUX_s_1_2_2(and_1169_nl, or_tmp_629, or_643_cse);
  and_dcpl_548 <= mux_228_nl AND and_dcpl_358 AND and_dcpl_521;
  or_648_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1030_nl <= nand_276_cse AND or_tmp_629;
  mux_tmp_227 <= MUX_s_1_2_2(and_1030_nl, or_tmp_629, or_648_cse);
  and_1031_nl <= nand_281_cse AND mux_tmp_227;
  mux_230_nl <= MUX_s_1_2_2(and_1031_nl, mux_tmp_227, or_643_cse);
  and_dcpl_550 <= mux_230_nl AND and_dcpl_362 AND and_dcpl_524;
  or_653_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR (rem_12cyc_st_3_3_2(1));
  and_1027_nl <= nand_198_cse AND or_tmp_629;
  mux_tmp_229 <= MUX_s_1_2_2(and_1027_nl, or_tmp_629, or_653_cse);
  and_1028_nl <= nand_276_cse AND mux_tmp_229;
  mux_tmp_230 <= MUX_s_1_2_2(and_1028_nl, mux_tmp_229, or_648_cse);
  and_1029_nl <= nand_281_cse AND mux_tmp_230;
  mux_233_nl <= MUX_s_1_2_2(and_1029_nl, mux_tmp_230, or_643_cse);
  and_dcpl_552 <= mux_233_nl AND and_dcpl_366 AND and_dcpl_527;
  or_660_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("01"));
  and_1023_nl <= nand_271_cse AND or_tmp_629;
  mux_tmp_232 <= MUX_s_1_2_2(and_1023_nl, or_tmp_629, or_660_cse);
  and_1024_nl <= nand_198_cse AND mux_tmp_232;
  mux_tmp_233 <= MUX_s_1_2_2(and_1024_nl, mux_tmp_232, or_653_cse);
  and_1025_nl <= nand_276_cse AND mux_tmp_233;
  mux_tmp_234 <= MUX_s_1_2_2(and_1025_nl, mux_tmp_233, or_648_cse);
  and_1026_nl <= nand_281_cse AND mux_tmp_234;
  mux_237_nl <= MUX_s_1_2_2(and_1026_nl, mux_tmp_234, or_643_cse);
  and_dcpl_554 <= mux_237_nl AND and_dcpl_370 AND and_dcpl_530;
  or_669_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR (rem_12cyc_st_5_3_2(1));
  and_1018_nl <= nand_189_cse AND or_tmp_629;
  mux_tmp_236 <= MUX_s_1_2_2(and_1018_nl, or_tmp_629, or_669_cse);
  and_1019_nl <= nand_271_cse AND mux_tmp_236;
  mux_tmp_237 <= MUX_s_1_2_2(and_1019_nl, mux_tmp_236, or_660_cse);
  and_1020_nl <= nand_198_cse AND mux_tmp_237;
  mux_tmp_238 <= MUX_s_1_2_2(and_1020_nl, mux_tmp_237, or_653_cse);
  and_1021_nl <= nand_276_cse AND mux_tmp_238;
  mux_tmp_239 <= MUX_s_1_2_2(and_1021_nl, mux_tmp_238, or_648_cse);
  and_1022_nl <= nand_281_cse AND mux_tmp_239;
  mux_242_nl <= MUX_s_1_2_2(and_1022_nl, mux_tmp_239, or_643_cse);
  and_dcpl_556 <= mux_242_nl AND and_dcpl_121 AND and_dcpl_119;
  or_680_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_6_3_2(1));
  and_1012_nl <= nand_215_cse AND or_tmp_629;
  mux_tmp_241 <= MUX_s_1_2_2(and_1012_nl, or_tmp_629, or_680_cse);
  and_1013_nl <= nand_189_cse AND mux_tmp_241;
  mux_tmp_242 <= MUX_s_1_2_2(and_1013_nl, mux_tmp_241, or_669_cse);
  and_1014_nl <= nand_271_cse AND mux_tmp_242;
  mux_tmp_243 <= MUX_s_1_2_2(and_1014_nl, mux_tmp_242, or_660_cse);
  and_1015_nl <= nand_198_cse AND mux_tmp_243;
  mux_tmp_244 <= MUX_s_1_2_2(and_1015_nl, mux_tmp_243, or_653_cse);
  and_1016_nl <= nand_276_cse AND mux_tmp_244;
  mux_tmp_245 <= MUX_s_1_2_2(and_1016_nl, mux_tmp_244, or_648_cse);
  and_1017_nl <= nand_281_cse AND mux_tmp_245;
  mux_248_nl <= MUX_s_1_2_2(and_1017_nl, mux_tmp_245, or_643_cse);
  and_dcpl_558 <= mux_248_nl AND and_dcpl_94 AND and_dcpl_92;
  or_693_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_7_3_2(1));
  and_1005_nl <= nand_212_cse AND or_tmp_629;
  mux_tmp_247 <= MUX_s_1_2_2(and_1005_nl, or_tmp_629, or_693_cse);
  and_1006_nl <= nand_215_cse AND mux_tmp_247;
  mux_tmp_248 <= MUX_s_1_2_2(and_1006_nl, mux_tmp_247, or_680_cse);
  and_1007_nl <= nand_189_cse AND mux_tmp_248;
  mux_tmp_249 <= MUX_s_1_2_2(and_1007_nl, mux_tmp_248, or_669_cse);
  and_1008_nl <= nand_271_cse AND mux_tmp_249;
  mux_tmp_250 <= MUX_s_1_2_2(and_1008_nl, mux_tmp_249, or_660_cse);
  and_1009_nl <= nand_198_cse AND mux_tmp_250;
  mux_tmp_251 <= MUX_s_1_2_2(and_1009_nl, mux_tmp_250, or_653_cse);
  and_1010_nl <= nand_276_cse AND mux_tmp_251;
  mux_tmp_252 <= MUX_s_1_2_2(and_1010_nl, mux_tmp_251, or_648_cse);
  and_1011_nl <= nand_281_cse AND mux_tmp_252;
  mux_255_nl <= MUX_s_1_2_2(and_1011_nl, mux_tmp_252, or_643_cse);
  and_dcpl_560 <= mux_255_nl AND and_dcpl_67 AND and_dcpl_65;
  or_708_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_8_3_2(1));
  and_997_nl <= nand_208_cse AND or_tmp_629;
  mux_tmp_254 <= MUX_s_1_2_2(and_997_nl, or_tmp_629, or_708_cse);
  and_998_nl <= nand_212_cse AND mux_tmp_254;
  mux_tmp_255 <= MUX_s_1_2_2(and_998_nl, mux_tmp_254, or_693_cse);
  and_999_nl <= nand_215_cse AND mux_tmp_255;
  mux_tmp_256 <= MUX_s_1_2_2(and_999_nl, mux_tmp_255, or_680_cse);
  and_1000_nl <= nand_189_cse AND mux_tmp_256;
  mux_tmp_257 <= MUX_s_1_2_2(and_1000_nl, mux_tmp_256, or_669_cse);
  and_1001_nl <= nand_271_cse AND mux_tmp_257;
  mux_tmp_258 <= MUX_s_1_2_2(and_1001_nl, mux_tmp_257, or_660_cse);
  and_1002_nl <= nand_198_cse AND mux_tmp_258;
  mux_tmp_259 <= MUX_s_1_2_2(and_1002_nl, mux_tmp_258, or_653_cse);
  and_1003_nl <= nand_276_cse AND mux_tmp_259;
  mux_tmp_260 <= MUX_s_1_2_2(and_1003_nl, mux_tmp_259, or_648_cse);
  and_1004_nl <= nand_281_cse AND mux_tmp_260;
  mux_263_nl <= MUX_s_1_2_2(and_1004_nl, mux_tmp_260, or_643_cse);
  and_dcpl_562 <= mux_263_nl AND and_dcpl_40 AND and_dcpl_38;
  and_988_nl <= nand_203_cse AND or_tmp_629;
  or_725_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("11")) OR (rem_12cyc_st_9_3_2(1));
  mux_tmp_262 <= MUX_s_1_2_2(and_988_nl, or_tmp_629, or_725_nl);
  and_989_nl <= nand_208_cse AND mux_tmp_262;
  mux_tmp_263 <= MUX_s_1_2_2(and_989_nl, mux_tmp_262, or_708_cse);
  and_990_nl <= nand_212_cse AND mux_tmp_263;
  mux_tmp_264 <= MUX_s_1_2_2(and_990_nl, mux_tmp_263, or_693_cse);
  and_991_nl <= nand_215_cse AND mux_tmp_264;
  mux_tmp_265 <= MUX_s_1_2_2(and_991_nl, mux_tmp_264, or_680_cse);
  and_992_nl <= nand_189_cse AND mux_tmp_265;
  mux_tmp_266 <= MUX_s_1_2_2(and_992_nl, mux_tmp_265, or_669_cse);
  and_993_nl <= nand_271_cse AND mux_tmp_266;
  mux_tmp_267 <= MUX_s_1_2_2(and_993_nl, mux_tmp_266, or_660_cse);
  and_994_nl <= nand_198_cse AND mux_tmp_267;
  mux_tmp_268 <= MUX_s_1_2_2(and_994_nl, mux_tmp_267, or_653_cse);
  and_995_nl <= nand_276_cse AND mux_tmp_268;
  mux_tmp_269 <= MUX_s_1_2_2(and_995_nl, mux_tmp_268, or_648_cse);
  and_996_nl <= nand_281_cse AND mux_tmp_269;
  mux_272_nl <= MUX_s_1_2_2(and_996_nl, mux_tmp_269, or_643_cse);
  and_dcpl_564 <= mux_272_nl AND and_dcpl_13 AND and_dcpl_11;
  and_tmp_179 <= (NOT(main_stage_0_8 AND asn_itm_7 AND CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_7_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_9
      AND asn_itm_8 AND CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_8_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_10
      AND asn_itm_9 AND CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_9_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_3
      AND asn_itm_2 AND CONV_SL_1_1(rem_12cyc_st_2_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_4
      AND asn_itm_3 AND CONV_SL_1_1(rem_12cyc_st_3_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_5
      AND asn_itm_4 AND CONV_SL_1_1(rem_12cyc_st_4_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_6
      AND asn_itm_5 AND CONV_SL_1_1(rem_12cyc_st_5_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_7
      AND asn_itm_6 AND CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_6_3_2=STD_LOGIC_VECTOR'("01")))) AND (NOT(main_stage_0_11
      AND asn_itm_10 AND CONV_SL_1_1(rem_12cyc_st_10_1_0=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(rem_12cyc_st_10_3_2=STD_LOGIC_VECTOR'("01")))) AND ((acc_tmp(1))
      OR (NOT((acc_tmp(0)) AND CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND ccs_ccore_start_rsci_idat)));
  and_987_nl <= (NOT((rem_12cyc_3_2(0)) AND CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11"))))
      AND and_tmp_179;
  or_735_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR (rem_12cyc_3_2(1));
  mux_tmp_271 <= MUX_s_1_2_2(and_987_nl, and_tmp_179, or_735_nl);
  and_dcpl_568 <= and_dcpl_292 AND (acc_tmp(1));
  and_dcpl_569 <= and_dcpl_568 AND and_dcpl_291;
  and_dcpl_570 <= CONV_SL_1_1(rem_12cyc_st_2_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_571 <= and_dcpl_570 AND (NOT (rem_12cyc_st_2_1_0(1)));
  or_tmp_733 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_748_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_436_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_733));
  mux_274_nl <= MUX_s_1_2_2(nor_436_nl, or_tmp_733, or_748_cse);
  and_dcpl_573 <= mux_274_nl AND and_dcpl_298 AND and_dcpl_571;
  and_dcpl_574 <= CONV_SL_1_1(rem_12cyc_st_3_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_575 <= and_dcpl_574 AND (NOT (rem_12cyc_st_3_1_0(1)));
  or_753_cse <= (rem_12cyc_st_2_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_180 <= or_753_cse AND or_tmp_733;
  nor_435_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_180));
  mux_275_nl <= MUX_s_1_2_2(nor_435_nl, and_tmp_180, or_748_cse);
  and_dcpl_577 <= mux_275_nl AND and_dcpl_304 AND and_dcpl_575;
  and_dcpl_578 <= CONV_SL_1_1(rem_12cyc_st_4_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_579 <= and_dcpl_578 AND (NOT (rem_12cyc_st_4_1_0(1)));
  or_757_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_182 <= or_753_cse AND or_757_cse AND or_tmp_733;
  nor_434_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_182));
  mux_276_nl <= MUX_s_1_2_2(nor_434_nl, and_tmp_182, or_748_cse);
  and_dcpl_581 <= mux_276_nl AND and_dcpl_310 AND and_dcpl_579;
  and_dcpl_582 <= CONV_SL_1_1(rem_12cyc_st_5_3_2=STD_LOGIC_VECTOR'("10"));
  and_dcpl_583 <= and_dcpl_582 AND (NOT (rem_12cyc_st_5_1_0(1)));
  or_762_cse <= (rem_12cyc_st_4_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_185 <= or_753_cse AND or_757_cse AND or_762_cse AND or_tmp_733;
  nor_433_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_185));
  mux_277_nl <= MUX_s_1_2_2(nor_433_nl, and_tmp_185, or_748_cse);
  and_dcpl_585 <= mux_277_nl AND and_dcpl_316 AND and_dcpl_583;
  or_768_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_189 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND or_tmp_733;
  nor_432_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_189));
  mux_278_nl <= MUX_s_1_2_2(nor_432_nl, and_tmp_189, or_748_cse);
  and_dcpl_589 <= mux_278_nl AND and_dcpl_112 AND and_dcpl_126 AND (NOT (rem_12cyc_st_6_1_0(1)));
  or_775_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_430_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_733));
  mux_279_nl <= MUX_s_1_2_2(nor_430_nl, or_tmp_733, or_775_cse);
  and_tmp_193 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_279_nl;
  nor_431_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_193));
  mux_280_nl <= MUX_s_1_2_2(nor_431_nl, and_tmp_193, or_748_cse);
  and_dcpl_593 <= mux_280_nl AND and_dcpl_85 AND and_dcpl_99 AND (NOT (rem_12cyc_st_7_1_0(0)));
  or_784_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_427_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_733));
  mux_tmp_279 <= MUX_s_1_2_2(nor_427_nl, or_tmp_733, or_784_cse);
  nor_428_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_279));
  mux_282_nl <= MUX_s_1_2_2(nor_428_nl, mux_tmp_279, or_775_cse);
  and_tmp_197 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_282_nl;
  nor_429_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_197));
  mux_283_nl <= MUX_s_1_2_2(nor_429_nl, and_tmp_197, or_748_cse);
  and_dcpl_597 <= mux_283_nl AND and_dcpl_58 AND and_dcpl_72 AND (NOT (rem_12cyc_st_8_1_0(0)));
  or_795_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_423_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_733));
  mux_tmp_282 <= MUX_s_1_2_2(nor_423_nl, or_tmp_733, or_795_cse);
  nor_424_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_282));
  mux_tmp_283 <= MUX_s_1_2_2(nor_424_nl, mux_tmp_282, or_784_cse);
  nor_425_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_283));
  mux_286_nl <= MUX_s_1_2_2(nor_425_nl, mux_tmp_283, or_775_cse);
  and_tmp_201 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_286_nl;
  nor_426_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_201));
  mux_287_nl <= MUX_s_1_2_2(nor_426_nl, and_tmp_201, or_748_cse);
  and_dcpl_601 <= mux_287_nl AND and_dcpl_31 AND and_dcpl_45 AND (NOT (rem_12cyc_st_9_1_0(0)));
  nor_418_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_733));
  or_808_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_286 <= MUX_s_1_2_2(nor_418_nl, or_tmp_733, or_808_nl);
  nor_419_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_286));
  mux_tmp_287 <= MUX_s_1_2_2(nor_419_nl, mux_tmp_286, or_795_cse);
  nor_420_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_287));
  mux_tmp_288 <= MUX_s_1_2_2(nor_420_nl, mux_tmp_287, or_784_cse);
  nor_421_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_288));
  mux_291_nl <= MUX_s_1_2_2(nor_421_nl, mux_tmp_288, or_775_cse);
  and_tmp_205 <= or_753_cse AND or_757_cse AND or_762_cse AND or_768_cse AND mux_291_nl;
  nor_422_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_205));
  mux_292_nl <= MUX_s_1_2_2(nor_422_nl, and_tmp_205, or_748_cse);
  and_dcpl_605 <= mux_292_nl AND and_dcpl_4 AND and_dcpl_18 AND (NOT (rem_12cyc_st_10_1_0(0)));
  or_tmp_808 <= CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(acc_1_tmp(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR (NOT ccs_ccore_start_rsci_idat);
  nor_409_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_808));
  or_823_nl <= (NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_291 <= MUX_s_1_2_2(nor_409_nl, or_tmp_808, or_823_nl);
  nor_410_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_291));
  or_822_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_292 <= MUX_s_1_2_2(nor_410_nl, mux_tmp_291, or_822_nl);
  nor_411_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_292));
  or_821_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_293 <= MUX_s_1_2_2(nor_411_nl, mux_tmp_292, or_821_nl);
  nor_412_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_293));
  or_820_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_294 <= MUX_s_1_2_2(nor_412_nl, mux_tmp_293, or_820_nl);
  nor_413_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_294));
  or_819_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_295 <= MUX_s_1_2_2(nor_413_nl, mux_tmp_294, or_819_nl);
  nor_414_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_295));
  or_818_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_296 <= MUX_s_1_2_2(nor_414_nl, mux_tmp_295, or_818_nl);
  nor_415_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_296));
  or_817_nl <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_297 <= MUX_s_1_2_2(nor_415_nl, mux_tmp_296, or_817_nl);
  nor_416_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_297));
  or_816_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_298 <= MUX_s_1_2_2(nor_416_nl, mux_tmp_297, or_816_nl);
  nor_417_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_298));
  or_815_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("00"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_301_nl <= MUX_s_1_2_2(nor_417_nl, mux_tmp_298, or_815_nl);
  and_tmp_206 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("00"))) AND mux_301_nl;
  and_dcpl_610 <= and_dcpl_568 AND and_dcpl_355;
  or_tmp_820 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_837_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_408_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_820));
  mux_302_nl <= MUX_s_1_2_2(nor_408_nl, or_tmp_820, or_837_cse);
  and_dcpl_612 <= mux_302_nl AND and_dcpl_358 AND and_dcpl_571;
  nand_84_cse <= NOT((rem_12cyc_st_2_3_2(1)) AND asn_itm_2 AND main_stage_0_3 AND
      (rem_12cyc_st_2_1_0(0)));
  or_842_cse <= (rem_12cyc_st_2_1_0(1)) OR (rem_12cyc_st_2_3_2(0));
  and_986_nl <= nand_84_cse AND or_tmp_820;
  mux_tmp_301 <= MUX_s_1_2_2(and_986_nl, or_tmp_820, or_842_cse);
  nor_407_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_301));
  mux_304_nl <= MUX_s_1_2_2(nor_407_nl, mux_tmp_301, or_837_cse);
  and_dcpl_614 <= mux_304_nl AND and_dcpl_362 AND and_dcpl_575;
  or_847_cse <= (rem_12cyc_st_3_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"));
  and_984_nl <= nand_274_cse AND or_tmp_820;
  mux_tmp_303 <= MUX_s_1_2_2(and_984_nl, or_tmp_820, or_847_cse);
  and_985_nl <= nand_84_cse AND mux_tmp_303;
  mux_tmp_304 <= MUX_s_1_2_2(and_985_nl, mux_tmp_303, or_842_cse);
  nor_406_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_304));
  mux_307_nl <= MUX_s_1_2_2(nor_406_nl, mux_tmp_304, or_837_cse);
  and_dcpl_616 <= mux_307_nl AND and_dcpl_366 AND and_dcpl_579;
  nand_79_cse <= NOT((rem_12cyc_st_4_3_2(1)) AND asn_itm_4 AND main_stage_0_5 AND
      (rem_12cyc_st_4_1_0(0)));
  or_854_cse <= (rem_12cyc_st_4_1_0(1)) OR (rem_12cyc_st_4_3_2(0));
  and_981_nl <= nand_79_cse AND or_tmp_820;
  mux_tmp_306 <= MUX_s_1_2_2(and_981_nl, or_tmp_820, or_854_cse);
  and_982_nl <= nand_274_cse AND mux_tmp_306;
  mux_tmp_307 <= MUX_s_1_2_2(and_982_nl, mux_tmp_306, or_847_cse);
  and_983_nl <= nand_84_cse AND mux_tmp_307;
  mux_tmp_308 <= MUX_s_1_2_2(and_983_nl, mux_tmp_307, or_842_cse);
  nor_405_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_308));
  mux_311_nl <= MUX_s_1_2_2(nor_405_nl, mux_tmp_308, or_837_cse);
  and_dcpl_618 <= mux_311_nl AND and_dcpl_370 AND and_dcpl_583;
  or_863_cse <= (rem_12cyc_st_5_1_0(1)) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"));
  and_977_nl <= nand_267_cse AND or_tmp_820;
  mux_tmp_310 <= MUX_s_1_2_2(and_977_nl, or_tmp_820, or_863_cse);
  and_978_nl <= nand_79_cse AND mux_tmp_310;
  mux_tmp_311 <= MUX_s_1_2_2(and_978_nl, mux_tmp_310, or_854_cse);
  and_979_nl <= nand_274_cse AND mux_tmp_311;
  mux_tmp_312 <= MUX_s_1_2_2(and_979_nl, mux_tmp_311, or_847_cse);
  and_980_nl <= nand_84_cse AND mux_tmp_312;
  mux_tmp_313 <= MUX_s_1_2_2(and_980_nl, mux_tmp_312, or_842_cse);
  nor_404_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_313));
  mux_316_nl <= MUX_s_1_2_2(nor_404_nl, mux_tmp_313, or_837_cse);
  and_dcpl_622 <= mux_316_nl AND and_dcpl_112 AND and_dcpl_129 AND (NOT (rem_12cyc_st_6_1_0(1)));
  or_874_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_402_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_820));
  mux_tmp_315 <= MUX_s_1_2_2(nor_402_nl, or_tmp_820, or_874_cse);
  and_973_nl <= nand_267_cse AND mux_tmp_315;
  mux_tmp_316 <= MUX_s_1_2_2(and_973_nl, mux_tmp_315, or_863_cse);
  and_974_nl <= nand_79_cse AND mux_tmp_316;
  mux_tmp_317 <= MUX_s_1_2_2(and_974_nl, mux_tmp_316, or_854_cse);
  and_975_nl <= nand_274_cse AND mux_tmp_317;
  mux_tmp_318 <= MUX_s_1_2_2(and_975_nl, mux_tmp_317, or_847_cse);
  and_976_nl <= nand_84_cse AND mux_tmp_318;
  mux_tmp_319 <= MUX_s_1_2_2(and_976_nl, mux_tmp_318, or_842_cse);
  nor_403_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_319));
  mux_322_nl <= MUX_s_1_2_2(nor_403_nl, mux_tmp_319, or_837_cse);
  and_dcpl_625 <= mux_322_nl AND and_dcpl_85 AND and_dcpl_99 AND (rem_12cyc_st_7_1_0(0));
  or_887_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_399_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_820));
  mux_tmp_321 <= MUX_s_1_2_2(nor_399_nl, or_tmp_820, or_887_cse);
  nor_400_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_321));
  mux_tmp_322 <= MUX_s_1_2_2(nor_400_nl, mux_tmp_321, or_874_cse);
  and_969_nl <= nand_267_cse AND mux_tmp_322;
  mux_tmp_323 <= MUX_s_1_2_2(and_969_nl, mux_tmp_322, or_863_cse);
  and_970_nl <= nand_79_cse AND mux_tmp_323;
  mux_tmp_324 <= MUX_s_1_2_2(and_970_nl, mux_tmp_323, or_854_cse);
  and_971_nl <= nand_274_cse AND mux_tmp_324;
  mux_tmp_325 <= MUX_s_1_2_2(and_971_nl, mux_tmp_324, or_847_cse);
  and_972_nl <= nand_84_cse AND mux_tmp_325;
  mux_tmp_326 <= MUX_s_1_2_2(and_972_nl, mux_tmp_325, or_842_cse);
  nor_401_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_326));
  mux_329_nl <= MUX_s_1_2_2(nor_401_nl, mux_tmp_326, or_837_cse);
  and_dcpl_628 <= mux_329_nl AND and_dcpl_58 AND and_dcpl_72 AND (rem_12cyc_st_8_1_0(0));
  or_902_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_395_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_820));
  mux_tmp_328 <= MUX_s_1_2_2(nor_395_nl, or_tmp_820, or_902_cse);
  nor_396_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_328));
  mux_tmp_329 <= MUX_s_1_2_2(nor_396_nl, mux_tmp_328, or_887_cse);
  nor_397_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_329));
  mux_tmp_330 <= MUX_s_1_2_2(nor_397_nl, mux_tmp_329, or_874_cse);
  and_965_nl <= nand_267_cse AND mux_tmp_330;
  mux_tmp_331 <= MUX_s_1_2_2(and_965_nl, mux_tmp_330, or_863_cse);
  and_966_nl <= nand_79_cse AND mux_tmp_331;
  mux_tmp_332 <= MUX_s_1_2_2(and_966_nl, mux_tmp_331, or_854_cse);
  and_967_nl <= nand_274_cse AND mux_tmp_332;
  mux_tmp_333 <= MUX_s_1_2_2(and_967_nl, mux_tmp_332, or_847_cse);
  and_968_nl <= nand_84_cse AND mux_tmp_333;
  mux_tmp_334 <= MUX_s_1_2_2(and_968_nl, mux_tmp_333, or_842_cse);
  nor_398_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_334));
  mux_337_nl <= MUX_s_1_2_2(nor_398_nl, mux_tmp_334, or_837_cse);
  and_dcpl_631 <= mux_337_nl AND and_dcpl_31 AND and_dcpl_45 AND (rem_12cyc_st_9_1_0(0));
  nor_390_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_820));
  or_919_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_336 <= MUX_s_1_2_2(nor_390_nl, or_tmp_820, or_919_nl);
  nor_391_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_336));
  mux_tmp_337 <= MUX_s_1_2_2(nor_391_nl, mux_tmp_336, or_902_cse);
  nor_392_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_337));
  mux_tmp_338 <= MUX_s_1_2_2(nor_392_nl, mux_tmp_337, or_887_cse);
  nor_393_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_338));
  mux_tmp_339 <= MUX_s_1_2_2(nor_393_nl, mux_tmp_338, or_874_cse);
  and_961_nl <= nand_267_cse AND mux_tmp_339;
  mux_tmp_340 <= MUX_s_1_2_2(and_961_nl, mux_tmp_339, or_863_cse);
  and_962_nl <= nand_79_cse AND mux_tmp_340;
  mux_tmp_341 <= MUX_s_1_2_2(and_962_nl, mux_tmp_340, or_854_cse);
  and_963_nl <= nand_274_cse AND mux_tmp_341;
  mux_tmp_342 <= MUX_s_1_2_2(and_963_nl, mux_tmp_341, or_847_cse);
  and_964_nl <= nand_84_cse AND mux_tmp_342;
  mux_tmp_343 <= MUX_s_1_2_2(and_964_nl, mux_tmp_342, or_842_cse);
  nor_394_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_343));
  mux_346_nl <= MUX_s_1_2_2(nor_394_nl, mux_tmp_343, or_837_cse);
  and_dcpl_634 <= mux_346_nl AND and_dcpl_4 AND and_dcpl_18 AND (rem_12cyc_st_10_1_0(0));
  or_tmp_921 <= CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10")) OR (acc_1_tmp(1)) OR
      nand_250_cse;
  nor_380_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_921));
  or_938_nl <= (NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_345 <= MUX_s_1_2_2(nor_380_nl, or_tmp_921, or_938_nl);
  nor_381_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_345));
  or_937_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_346 <= MUX_s_1_2_2(nor_381_nl, mux_tmp_345, or_937_nl);
  nor_382_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_346));
  or_936_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_347 <= MUX_s_1_2_2(nor_382_nl, mux_tmp_346, or_936_nl);
  nor_383_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_347));
  or_935_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_348 <= MUX_s_1_2_2(nor_383_nl, mux_tmp_347, or_935_nl);
  nor_384_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_348));
  or_934_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_349 <= MUX_s_1_2_2(nor_384_nl, mux_tmp_348, or_934_nl);
  nor_385_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_349));
  or_933_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_350 <= MUX_s_1_2_2(nor_385_nl, mux_tmp_349, or_933_nl);
  nor_386_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_350));
  or_932_nl <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_351 <= MUX_s_1_2_2(nor_386_nl, mux_tmp_350, or_932_nl);
  nor_387_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_351));
  or_931_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_352 <= MUX_s_1_2_2(nor_387_nl, mux_tmp_351, or_931_nl);
  nor_388_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_352));
  or_930_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("01"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_tmp_353 <= MUX_s_1_2_2(nor_388_nl, mux_tmp_352, or_930_nl);
  nor_389_nl <= NOT((rem_12cyc_1_0(0)) OR (NOT mux_tmp_353));
  or_929_nl <= (NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_1_0(1));
  mux_tmp_354 <= MUX_s_1_2_2(nor_389_nl, mux_tmp_353, or_929_nl);
  and_dcpl_638 <= and_dcpl_568 AND and_dcpl_393;
  and_dcpl_639 <= and_dcpl_570 AND (rem_12cyc_st_2_1_0(1));
  or_tmp_934 <= CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_54;
  or_952_cse <= CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10"));
  nor_379_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_934));
  mux_357_nl <= MUX_s_1_2_2(nor_379_nl, or_tmp_934, or_952_cse);
  and_dcpl_641 <= mux_357_nl AND and_dcpl_298 AND and_dcpl_639;
  and_dcpl_642 <= and_dcpl_574 AND (rem_12cyc_st_3_1_0(1));
  or_957_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_2_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_2) OR (NOT main_stage_0_3) OR (rem_12cyc_st_2_1_0(0));
  and_tmp_207 <= or_957_cse AND or_tmp_934;
  nor_378_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_207));
  mux_358_nl <= MUX_s_1_2_2(nor_378_nl, and_tmp_207, or_952_cse);
  and_dcpl_644 <= mux_358_nl AND and_dcpl_304 AND and_dcpl_642;
  and_dcpl_645 <= and_dcpl_578 AND (rem_12cyc_st_4_1_0(1));
  or_961_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_3) OR (NOT main_stage_0_4) OR (rem_12cyc_st_3_1_0(0));
  and_tmp_209 <= or_957_cse AND or_961_cse AND or_tmp_934;
  nor_377_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_209));
  mux_359_nl <= MUX_s_1_2_2(nor_377_nl, and_tmp_209, or_952_cse);
  and_dcpl_647 <= mux_359_nl AND and_dcpl_310 AND and_dcpl_645;
  and_dcpl_648 <= and_dcpl_582 AND (rem_12cyc_st_5_1_0(1));
  or_966_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_4_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_4) OR (NOT main_stage_0_5) OR (rem_12cyc_st_4_1_0(0));
  and_tmp_212 <= or_957_cse AND or_961_cse AND or_966_cse AND or_tmp_934;
  nor_376_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_212));
  mux_360_nl <= MUX_s_1_2_2(nor_376_nl, and_tmp_212, or_952_cse);
  and_dcpl_650 <= mux_360_nl AND and_dcpl_316 AND and_dcpl_648;
  or_972_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"))
      OR (NOT asn_itm_5) OR (NOT main_stage_0_6) OR (rem_12cyc_st_5_1_0(0));
  and_tmp_216 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND or_tmp_934;
  nor_375_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_216));
  mux_361_nl <= MUX_s_1_2_2(nor_375_nl, and_tmp_216, or_952_cse);
  and_dcpl_653 <= mux_361_nl AND and_dcpl_112 AND and_dcpl_126 AND (rem_12cyc_st_6_1_0(1));
  or_979_cse <= CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_6_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_373_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_934));
  mux_362_nl <= MUX_s_1_2_2(nor_373_nl, or_tmp_934, or_979_cse);
  and_tmp_220 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_362_nl;
  nor_374_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_220));
  mux_363_nl <= MUX_s_1_2_2(nor_374_nl, and_tmp_220, or_952_cse);
  and_dcpl_657 <= mux_363_nl AND and_dcpl_85 AND and_dcpl_104 AND (NOT (rem_12cyc_st_7_1_0(0)));
  or_988_cse <= CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_7_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_370_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_934));
  mux_tmp_362 <= MUX_s_1_2_2(nor_370_nl, or_tmp_934, or_988_cse);
  nor_371_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_362));
  mux_365_nl <= MUX_s_1_2_2(nor_371_nl, mux_tmp_362, or_979_cse);
  and_tmp_224 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_365_nl;
  nor_372_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_224));
  mux_366_nl <= MUX_s_1_2_2(nor_372_nl, and_tmp_224, or_952_cse);
  and_dcpl_661 <= mux_366_nl AND and_dcpl_58 AND and_dcpl_77 AND (NOT (rem_12cyc_st_8_1_0(0)));
  or_999_cse <= CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_8_3_2/=STD_LOGIC_VECTOR'("10"));
  nor_366_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_934));
  mux_tmp_365 <= MUX_s_1_2_2(nor_366_nl, or_tmp_934, or_999_cse);
  nor_367_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_365));
  mux_tmp_366 <= MUX_s_1_2_2(nor_367_nl, mux_tmp_365, or_988_cse);
  nor_368_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_366));
  mux_369_nl <= MUX_s_1_2_2(nor_368_nl, mux_tmp_366, or_979_cse);
  and_tmp_228 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_369_nl;
  nor_369_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_228));
  mux_370_nl <= MUX_s_1_2_2(nor_369_nl, and_tmp_228, or_952_cse);
  and_dcpl_665 <= mux_370_nl AND and_dcpl_31 AND and_dcpl_50 AND (NOT (rem_12cyc_st_9_1_0(0)));
  nor_361_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_934));
  or_1012_nl <= CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(rem_12cyc_st_9_3_2/=STD_LOGIC_VECTOR'("10"));
  mux_tmp_369 <= MUX_s_1_2_2(nor_361_nl, or_tmp_934, or_1012_nl);
  nor_362_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_369));
  mux_tmp_370 <= MUX_s_1_2_2(nor_362_nl, mux_tmp_369, or_999_cse);
  nor_363_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_370));
  mux_tmp_371 <= MUX_s_1_2_2(nor_363_nl, mux_tmp_370, or_988_cse);
  nor_364_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_371));
  mux_374_nl <= MUX_s_1_2_2(nor_364_nl, mux_tmp_371, or_979_cse);
  and_tmp_232 <= or_957_cse AND or_961_cse AND or_966_cse AND or_972_cse AND mux_374_nl;
  nor_365_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT and_tmp_232));
  mux_375_nl <= MUX_s_1_2_2(nor_365_nl, and_tmp_232, or_952_cse);
  and_dcpl_669 <= mux_375_nl AND and_dcpl_4 AND and_dcpl_23 AND (NOT (rem_12cyc_st_10_1_0(0)));
  or_tmp_1009 <= CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(acc_1_tmp(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR (NOT ccs_ccore_start_rsci_idat);
  nor_352_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_1009));
  or_1027_nl <= (NOT main_stage_0_11) OR (NOT asn_itm_10) OR CONV_SL_1_1(rem_12cyc_st_10_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_10_3_2(0));
  mux_tmp_374 <= MUX_s_1_2_2(nor_352_nl, or_tmp_1009, or_1027_nl);
  nor_353_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_374));
  or_1026_nl <= (NOT main_stage_0_7) OR (NOT asn_itm_6) OR CONV_SL_1_1(rem_12cyc_st_6_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_6_3_2(0));
  mux_tmp_375 <= MUX_s_1_2_2(nor_353_nl, mux_tmp_374, or_1026_nl);
  nor_354_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_375));
  or_1025_nl <= (NOT main_stage_0_6) OR (NOT asn_itm_5) OR CONV_SL_1_1(rem_12cyc_st_5_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_5_3_2(0));
  mux_tmp_376 <= MUX_s_1_2_2(nor_354_nl, mux_tmp_375, or_1025_nl);
  nor_355_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_376));
  or_1024_nl <= (NOT main_stage_0_5) OR (NOT asn_itm_4) OR CONV_SL_1_1(rem_12cyc_st_4_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_4_3_2(0));
  mux_tmp_377 <= MUX_s_1_2_2(nor_355_nl, mux_tmp_376, or_1024_nl);
  nor_356_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_377));
  or_1023_nl <= (NOT main_stage_0_4) OR (NOT asn_itm_3) OR CONV_SL_1_1(rem_12cyc_st_3_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_3_3_2(0));
  mux_tmp_378 <= MUX_s_1_2_2(nor_356_nl, mux_tmp_377, or_1023_nl);
  nor_357_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_378));
  or_1022_nl <= (NOT main_stage_0_3) OR (NOT asn_itm_2) OR CONV_SL_1_1(rem_12cyc_st_2_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_2_3_2(0));
  mux_tmp_379 <= MUX_s_1_2_2(nor_357_nl, mux_tmp_378, or_1022_nl);
  nor_358_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_379));
  or_1021_nl <= (NOT main_stage_0_10) OR (NOT asn_itm_9) OR CONV_SL_1_1(rem_12cyc_st_9_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_9_3_2(0));
  mux_tmp_380 <= MUX_s_1_2_2(nor_358_nl, mux_tmp_379, or_1021_nl);
  nor_359_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_380));
  or_1020_nl <= (NOT main_stage_0_9) OR (NOT asn_itm_8) OR CONV_SL_1_1(rem_12cyc_st_8_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_8_3_2(0));
  mux_tmp_381 <= MUX_s_1_2_2(nor_359_nl, mux_tmp_380, or_1020_nl);
  nor_360_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_381));
  or_1019_nl <= (NOT main_stage_0_8) OR (NOT asn_itm_7) OR CONV_SL_1_1(rem_12cyc_st_7_1_0/=STD_LOGIC_VECTOR'("10"))
      OR (rem_12cyc_st_7_3_2(0));
  mux_384_nl <= MUX_s_1_2_2(nor_360_nl, mux_tmp_381, or_1019_nl);
  and_tmp_233 <= ((NOT main_stage_0_2) OR (NOT asn_itm_1) OR CONV_SL_1_1(rem_12cyc_3_2/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(rem_12cyc_1_0/=STD_LOGIC_VECTOR'("10"))) AND mux_384_nl;
  and_dcpl_673 <= and_dcpl_568 AND and_dcpl_430;
  or_tmp_1021 <= (NOT(CONV_SL_1_1(rem_12cyc_1_0=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(rem_12cyc_3_2=STD_LOGIC_VECTOR'("10"))))
      OR not_tmp_54;
  nand_57_cse <= NOT(CONV_SL_1_1(acc_1_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(acc_tmp=STD_LOGIC_VECTOR'("10")));
  nor_351_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT or_tmp_1021));
  mux_385_nl <= MUX_s_1_2_2(nor_351_nl, or_tmp_1021, nand_57_cse);
  and_dcpl_675 <= mux_385_nl AND and_dcpl_358 AND and_dcpl_639;
  or_1045_cse <= (NOT (rem_12cyc_st_2_1_0(1))) OR (rem_12cyc_st_2_3_2(0));
  and_960_nl <= nand_84_cse AND or_tmp_1021;
  mux_tmp_384 <= MUX_s_1_2_2(and_960_nl, or_tmp_1021, or_1045_cse);
  nor_350_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_384));
  mux_387_nl <= MUX_s_1_2_2(nor_350_nl, mux_tmp_384, nand_57_cse);
  and_dcpl_677 <= mux_387_nl AND and_dcpl_362 AND and_dcpl_642;
  or_1050_cse <= (NOT (rem_12cyc_st_3_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_3_3_2/=STD_LOGIC_VECTOR'("10"));
  and_958_nl <= nand_274_cse AND or_tmp_1021;
  mux_tmp_386 <= MUX_s_1_2_2(and_958_nl, or_tmp_1021, or_1050_cse);
  and_959_nl <= nand_84_cse AND mux_tmp_386;
  mux_tmp_387 <= MUX_s_1_2_2(and_959_nl, mux_tmp_386, or_1045_cse);
  nor_349_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_387));
  mux_390_nl <= MUX_s_1_2_2(nor_349_nl, mux_tmp_387, nand_57_cse);
  and_dcpl_679 <= mux_390_nl AND and_dcpl_366 AND and_dcpl_645;
  or_1057_cse <= (NOT (rem_12cyc_st_4_1_0(1))) OR (rem_12cyc_st_4_3_2(0));
  and_955_nl <= nand_79_cse AND or_tmp_1021;
  mux_tmp_389 <= MUX_s_1_2_2(and_955_nl, or_tmp_1021, or_1057_cse);
  and_956_nl <= nand_274_cse AND mux_tmp_389;
  mux_tmp_390 <= MUX_s_1_2_2(and_956_nl, mux_tmp_389, or_1050_cse);
  and_957_nl <= nand_84_cse AND mux_tmp_390;
  mux_tmp_391 <= MUX_s_1_2_2(and_957_nl, mux_tmp_390, or_1045_cse);
  nor_348_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_391));
  mux_394_nl <= MUX_s_1_2_2(nor_348_nl, mux_tmp_391, nand_57_cse);
  and_dcpl_681 <= mux_394_nl AND and_dcpl_370 AND and_dcpl_648;
  or_1066_cse <= (NOT (rem_12cyc_st_5_1_0(1))) OR CONV_SL_1_1(rem_12cyc_st_5_3_2/=STD_LOGIC_VECTOR'("10"));
  and_951_nl <= nand_267_cse AND or_tmp_1021;
  mux_tmp_393 <= MUX_s_1_2_2(and_951_nl, or_tmp_1021, or_1066_cse);
  and_952_nl <= nand_79_cse AND mux_tmp_393;
  mux_tmp_394 <= MUX_s_1_2_2(and_952_nl, mux_tmp_393, or_1057_cse);
  and_953_nl <= nand_274_cse AND mux_tmp_394;
  mux_tmp_395 <= MUX_s_1_2_2(and_953_nl, mux_tmp_394, or_1050_cse);
  and_954_nl <= nand_84_cse AND mux_tmp_395;
  mux_tmp_396 <= MUX_s_1_2_2(and_954_nl, mux_tmp_395, or_1045_cse);
  nor_347_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_396));
  mux_399_nl <= MUX_s_1_2_2(nor_347_nl, mux_tmp_396, nand_57_cse);
  and_dcpl_684 <= mux_399_nl AND and_dcpl_112 AND and_dcpl_129 AND (rem_12cyc_st_6_1_0(1));
  nand_36_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_6_3_2=STD_LOGIC_VECTOR'("10")));
  nor_345_nl <= NOT(and_dcpl_111 OR (NOT or_tmp_1021));
  mux_tmp_398 <= MUX_s_1_2_2(nor_345_nl, or_tmp_1021, nand_36_cse);
  and_947_nl <= nand_267_cse AND mux_tmp_398;
  mux_tmp_399 <= MUX_s_1_2_2(and_947_nl, mux_tmp_398, or_1066_cse);
  and_948_nl <= nand_79_cse AND mux_tmp_399;
  mux_tmp_400 <= MUX_s_1_2_2(and_948_nl, mux_tmp_399, or_1057_cse);
  and_949_nl <= nand_274_cse AND mux_tmp_400;
  mux_tmp_401 <= MUX_s_1_2_2(and_949_nl, mux_tmp_400, or_1050_cse);
  and_950_nl <= nand_84_cse AND mux_tmp_401;
  mux_tmp_402 <= MUX_s_1_2_2(and_950_nl, mux_tmp_401, or_1045_cse);
  nor_346_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_402));
  mux_405_nl <= MUX_s_1_2_2(nor_346_nl, mux_tmp_402, nand_57_cse);
  and_dcpl_687 <= mux_405_nl AND and_dcpl_85 AND and_dcpl_104 AND (rem_12cyc_st_7_1_0(0));
  nand_29_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_7_3_2=STD_LOGIC_VECTOR'("10")));
  nor_342_nl <= NOT(and_dcpl_84 OR (NOT or_tmp_1021));
  mux_tmp_404 <= MUX_s_1_2_2(nor_342_nl, or_tmp_1021, nand_29_cse);
  nor_343_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_404));
  mux_tmp_405 <= MUX_s_1_2_2(nor_343_nl, mux_tmp_404, nand_36_cse);
  and_943_nl <= nand_267_cse AND mux_tmp_405;
  mux_tmp_406 <= MUX_s_1_2_2(and_943_nl, mux_tmp_405, or_1066_cse);
  and_944_nl <= nand_79_cse AND mux_tmp_406;
  mux_tmp_407 <= MUX_s_1_2_2(and_944_nl, mux_tmp_406, or_1057_cse);
  and_945_nl <= nand_274_cse AND mux_tmp_407;
  mux_tmp_408 <= MUX_s_1_2_2(and_945_nl, mux_tmp_407, or_1050_cse);
  and_946_nl <= nand_84_cse AND mux_tmp_408;
  mux_tmp_409 <= MUX_s_1_2_2(and_946_nl, mux_tmp_408, or_1045_cse);
  nor_344_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_409));
  mux_412_nl <= MUX_s_1_2_2(nor_344_nl, mux_tmp_409, nand_57_cse);
  and_dcpl_690 <= mux_412_nl AND and_dcpl_58 AND and_dcpl_77 AND (rem_12cyc_st_8_1_0(0));
  nand_21_cse <= NOT(CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(rem_12cyc_st_8_3_2=STD_LOGIC_VECTOR'("10")));
  nor_338_nl <= NOT(and_dcpl_57 OR (NOT or_tmp_1021));
  mux_tmp_411 <= MUX_s_1_2_2(nor_338_nl, or_tmp_1021, nand_21_cse);
  nor_339_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_411));
  mux_tmp_412 <= MUX_s_1_2_2(nor_339_nl, mux_tmp_411, nand_29_cse);
  nor_340_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_412));
  mux_tmp_413 <= MUX_s_1_2_2(nor_340_nl, mux_tmp_412, nand_36_cse);
  and_939_nl <= nand_267_cse AND mux_tmp_413;
  mux_tmp_414 <= MUX_s_1_2_2(and_939_nl, mux_tmp_413, or_1066_cse);
  and_940_nl <= nand_79_cse AND mux_tmp_414;
  mux_tmp_415 <= MUX_s_1_2_2(and_940_nl, mux_tmp_414, or_1057_cse);
  and_941_nl <= nand_274_cse AND mux_tmp_415;
  mux_tmp_416 <= MUX_s_1_2_2(and_941_nl, mux_tmp_415, or_1050_cse);
  and_942_nl <= nand_84_cse AND mux_tmp_416;
  mux_tmp_417 <= MUX_s_1_2_2(and_942_nl, mux_tmp_416, or_1045_cse);
  nor_341_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_417));
  mux_420_nl <= MUX_s_1_2_2(nor_341_nl, mux_tmp_417, nand_57_cse);
  and_dcpl_693 <= mux_420_nl AND and_dcpl_31 AND and_dcpl_50 AND (rem_12cyc_st_9_1_0(0));
  nor_333_nl <= NOT(and_dcpl_30 OR (NOT or_tmp_1021));
  nand_12_nl <= NOT(CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11")) AND CONV_SL_1_1(rem_12cyc_st_9_3_2=STD_LOGIC_VECTOR'("10")));
  mux_tmp_419 <= MUX_s_1_2_2(nor_333_nl, or_tmp_1021, nand_12_nl);
  nor_334_nl <= NOT(and_dcpl_57 OR (NOT mux_tmp_419));
  mux_tmp_420 <= MUX_s_1_2_2(nor_334_nl, mux_tmp_419, nand_21_cse);
  nor_335_nl <= NOT(and_dcpl_84 OR (NOT mux_tmp_420));
  mux_tmp_421 <= MUX_s_1_2_2(nor_335_nl, mux_tmp_420, nand_29_cse);
  nor_336_nl <= NOT(and_dcpl_111 OR (NOT mux_tmp_421));
  mux_tmp_422 <= MUX_s_1_2_2(nor_336_nl, mux_tmp_421, nand_36_cse);
  and_935_nl <= nand_267_cse AND mux_tmp_422;
  mux_tmp_423 <= MUX_s_1_2_2(and_935_nl, mux_tmp_422, or_1066_cse);
  and_936_nl <= nand_79_cse AND mux_tmp_423;
  mux_tmp_424 <= MUX_s_1_2_2(and_936_nl, mux_tmp_423, or_1057_cse);
  and_937_nl <= nand_274_cse AND mux_tmp_424;
  mux_tmp_425 <= MUX_s_1_2_2(and_937_nl, mux_tmp_424, or_1050_cse);
  and_938_nl <= nand_84_cse AND mux_tmp_425;
  mux_tmp_426 <= MUX_s_1_2_2(and_938_nl, mux_tmp_425, or_1045_cse);
  nor_337_nl <= NOT(ccs_ccore_start_rsci_idat OR (NOT mux_tmp_426));
  mux_429_nl <= MUX_s_1_2_2(nor_337_nl, mux_tmp_426, nand_57_cse);
  and_dcpl_696 <= mux_429_nl AND and_dcpl_4 AND and_dcpl_23 AND (rem_12cyc_st_10_1_0(0));
  or_tmp_1122 <= CONV_SL_1_1(acc_tmp/=STD_LOGIC_VECTOR'("10")) OR nand_222_cse;
  nor_324_nl <= NOT((rem_12cyc_st_10_3_2(1)) OR (NOT or_tmp_1122));
  nand_1_nl <= NOT(main_stage_0_11 AND asn_itm_10 AND CONV_SL_1_1(rem_12cyc_st_10_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_10_3_2(0))));
  mux_tmp_428 <= MUX_s_1_2_2(nor_324_nl, or_tmp_1122, nand_1_nl);
  nor_325_nl <= NOT((rem_12cyc_st_6_3_2(1)) OR (NOT mux_tmp_428));
  nand_2_nl <= NOT(main_stage_0_7 AND asn_itm_6 AND CONV_SL_1_1(rem_12cyc_st_6_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_6_3_2(0))));
  mux_tmp_429 <= MUX_s_1_2_2(nor_325_nl, mux_tmp_428, nand_2_nl);
  nor_326_nl <= NOT((rem_12cyc_st_5_3_2(1)) OR (NOT mux_tmp_429));
  nand_3_nl <= NOT(main_stage_0_6 AND asn_itm_5 AND CONV_SL_1_1(rem_12cyc_st_5_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_5_3_2(0))));
  mux_tmp_430 <= MUX_s_1_2_2(nor_326_nl, mux_tmp_429, nand_3_nl);
  nor_327_nl <= NOT((rem_12cyc_st_4_3_2(1)) OR (NOT mux_tmp_430));
  nand_4_nl <= NOT(main_stage_0_5 AND asn_itm_4 AND CONV_SL_1_1(rem_12cyc_st_4_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_4_3_2(0))));
  mux_tmp_431 <= MUX_s_1_2_2(nor_327_nl, mux_tmp_430, nand_4_nl);
  nor_328_nl <= NOT((rem_12cyc_st_3_3_2(1)) OR (NOT mux_tmp_431));
  nand_5_nl <= NOT(main_stage_0_4 AND asn_itm_3 AND CONV_SL_1_1(rem_12cyc_st_3_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_3_3_2(0))));
  mux_tmp_432 <= MUX_s_1_2_2(nor_328_nl, mux_tmp_431, nand_5_nl);
  nor_329_nl <= NOT((rem_12cyc_st_2_3_2(1)) OR (NOT mux_tmp_432));
  nand_6_nl <= NOT(main_stage_0_3 AND asn_itm_2 AND CONV_SL_1_1(rem_12cyc_st_2_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_2_3_2(0))));
  mux_tmp_433 <= MUX_s_1_2_2(nor_329_nl, mux_tmp_432, nand_6_nl);
  nor_330_nl <= NOT((rem_12cyc_st_9_3_2(1)) OR (NOT mux_tmp_433));
  nand_7_nl <= NOT(main_stage_0_10 AND asn_itm_9 AND CONV_SL_1_1(rem_12cyc_st_9_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_9_3_2(0))));
  mux_tmp_434 <= MUX_s_1_2_2(nor_330_nl, mux_tmp_433, nand_7_nl);
  nor_331_nl <= NOT((rem_12cyc_st_8_3_2(1)) OR (NOT mux_tmp_434));
  nand_8_nl <= NOT(main_stage_0_9 AND asn_itm_8 AND CONV_SL_1_1(rem_12cyc_st_8_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_8_3_2(0))));
  mux_tmp_435 <= MUX_s_1_2_2(nor_331_nl, mux_tmp_434, nand_8_nl);
  nor_332_nl <= NOT((rem_12cyc_st_7_3_2(1)) OR (NOT mux_tmp_435));
  nand_9_nl <= NOT(main_stage_0_8 AND asn_itm_7 AND CONV_SL_1_1(rem_12cyc_st_7_1_0=STD_LOGIC_VECTOR'("11"))
      AND (NOT (rem_12cyc_st_7_3_2(0))));
  mux_tmp_436 <= MUX_s_1_2_2(nor_332_nl, mux_tmp_435, nand_9_nl);
  and_934_nl <= nand_223_cse AND mux_tmp_436;
  nand_11_nl <= NOT(main_stage_0_2 AND asn_itm_1 AND CONV_SL_1_1(rem_12cyc_3_2=STD_LOGIC_VECTOR'("10")));
  mux_tmp_437 <= MUX_s_1_2_2(and_934_nl, mux_tmp_436, nand_11_nl);
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( ccs_ccore_en = '1' ) THEN
        return_rsci_d <= MUX_v_64_2_2(result_sva_duc_mx0, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(qelse_acc_nl),
            64)), mux_13_nl);
        m_buf_sva_12 <= m_buf_sva_11;
        m_buf_sva_11 <= m_buf_sva_10;
        m_buf_sva_10 <= m_buf_sva_9;
        m_buf_sva_9 <= m_buf_sva_8;
        m_buf_sva_8 <= m_buf_sva_7;
        m_buf_sva_7 <= m_buf_sva_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        asn_itm_12 <= '0';
        asn_itm_11 <= '0';
        asn_itm_10 <= '0';
        asn_itm_9 <= '0';
        asn_itm_8 <= '0';
        asn_itm_7 <= '0';
        asn_itm_6 <= '0';
        asn_itm_5 <= '0';
        asn_itm_4 <= '0';
        asn_itm_3 <= '0';
        asn_itm_2 <= '0';
        asn_itm_1 <= '0';
        main_stage_0_2 <= '0';
        main_stage_0_3 <= '0';
        main_stage_0_4 <= '0';
        main_stage_0_5 <= '0';
        main_stage_0_6 <= '0';
        main_stage_0_7 <= '0';
        main_stage_0_8 <= '0';
        main_stage_0_9 <= '0';
        main_stage_0_10 <= '0';
        main_stage_0_11 <= '0';
        main_stage_0_12 <= '0';
        main_stage_0_13 <= '0';
      ELSIF ( ccs_ccore_en = '1' ) THEN
        asn_itm_12 <= asn_itm_11;
        asn_itm_11 <= asn_itm_10;
        asn_itm_10 <= asn_itm_9;
        asn_itm_9 <= asn_itm_8;
        asn_itm_8 <= asn_itm_7;
        asn_itm_7 <= asn_itm_6;
        asn_itm_6 <= asn_itm_5;
        asn_itm_5 <= asn_itm_4;
        asn_itm_4 <= asn_itm_3;
        asn_itm_3 <= asn_itm_2;
        asn_itm_2 <= asn_itm_1;
        asn_itm_1 <= ccs_ccore_start_rsci_idat;
        main_stage_0_2 <= '1';
        main_stage_0_3 <= main_stage_0_2;
        main_stage_0_4 <= main_stage_0_3;
        main_stage_0_5 <= main_stage_0_4;
        main_stage_0_6 <= main_stage_0_5;
        main_stage_0_7 <= main_stage_0_6;
        main_stage_0_8 <= main_stage_0_7;
        main_stage_0_9 <= main_stage_0_8;
        main_stage_0_10 <= main_stage_0_9;
        main_stage_0_11 <= main_stage_0_10;
        main_stage_0_12 <= main_stage_0_11;
        main_stage_0_13 <= main_stage_0_12;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        result_sva_duc <= STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000000");
      ELSIF ( (asn_itm_12 AND main_stage_0_13 AND ccs_ccore_en AND (NOT(CONV_SL_1_1(rem_12cyc_st_12_3_2=STD_LOGIC_VECTOR'("11")))))
          = '1' ) THEN
        result_sva_duc <= result_sva_duc_mx0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_12_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_12_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1203_cse = '1' ) THEN
        rem_12cyc_st_12_3_2 <= rem_12cyc_st_11_3_2;
        rem_12cyc_st_12_1_0 <= rem_12cyc_st_11_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1173_cse = '1' ) THEN
        rem_13_cmp_1_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_3_2_63_0, mut_3_3_63_0,
            mut_3_4_63_0, mut_3_5_63_0, mut_3_6_63_0, mut_3_7_63_0, mut_3_8_63_0,
            mut_3_9_63_0, mut_3_10_63_0, mut_3_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_294
            & and_dcpl_300 & and_dcpl_306 & and_dcpl_312 & and_dcpl_318 & and_dcpl_324
            & and_dcpl_330 & and_dcpl_336 & and_dcpl_342 & and_dcpl_348 & and_tmp_35));
        rem_13_cmp_1_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_2_63_0, mut_2_3_63_0,
            mut_2_4_63_0, mut_2_5_63_0, mut_2_6_63_0, mut_2_7_63_0, mut_2_8_63_0,
            mut_2_9_63_0, mut_2_10_63_0, mut_2_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_294
            & and_dcpl_300 & and_dcpl_306 & and_dcpl_312 & and_dcpl_318 & and_dcpl_324
            & and_dcpl_330 & and_dcpl_336 & and_dcpl_342 & and_dcpl_348 & and_tmp_35));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1175_cse = '1' ) THEN
        rem_13_cmp_2_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_5_2_63_0, mut_5_3_63_0,
            mut_5_4_63_0, mut_5_5_63_0, mut_5_6_63_0, mut_5_7_63_0, mut_5_8_63_0,
            mut_5_9_63_0, mut_5_10_63_0, mut_5_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_356
            & and_dcpl_360 & and_dcpl_364 & and_dcpl_368 & and_dcpl_372 & and_dcpl_376
            & and_dcpl_379 & and_dcpl_382 & and_dcpl_385 & and_dcpl_388 & mux_tmp_76));
        rem_13_cmp_2_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_4_2_63_0, mut_4_3_63_0,
            mut_4_4_63_0, mut_4_5_63_0, mut_4_6_63_0, mut_4_7_63_0, mut_4_8_63_0,
            mut_4_9_63_0, mut_4_10_63_0, mut_4_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_356
            & and_dcpl_360 & and_dcpl_364 & and_dcpl_368 & and_dcpl_372 & and_dcpl_376
            & and_dcpl_379 & and_dcpl_382 & and_dcpl_385 & and_dcpl_388 & mux_tmp_76));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1177_cse = '1' ) THEN
        rem_13_cmp_3_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_7_2_63_0, mut_7_3_63_0,
            mut_7_4_63_0, mut_7_5_63_0, mut_7_6_63_0, mut_7_7_63_0, mut_7_8_63_0,
            mut_7_9_63_0, mut_7_10_63_0, mut_7_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_394
            & and_dcpl_397 & and_dcpl_400 & and_dcpl_403 & and_dcpl_406 & and_dcpl_409
            & and_dcpl_413 & and_dcpl_417 & and_dcpl_421 & and_dcpl_425 & and_tmp_80));
        rem_13_cmp_3_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_6_2_63_0, mut_6_3_63_0,
            mut_6_4_63_0, mut_6_5_63_0, mut_6_6_63_0, mut_6_7_63_0, mut_6_8_63_0,
            mut_6_9_63_0, mut_6_10_63_0, mut_6_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_394
            & and_dcpl_397 & and_dcpl_400 & and_dcpl_403 & and_dcpl_406 & and_dcpl_409
            & and_dcpl_413 & and_dcpl_417 & and_dcpl_421 & and_dcpl_425 & and_tmp_80));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1179_cse = '1' ) THEN
        rem_13_cmp_4_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_9_2_63_0, mut_9_3_63_0,
            mut_9_4_63_0, mut_9_5_63_0, mut_9_6_63_0, mut_9_7_63_0, mut_9_8_63_0,
            mut_9_9_63_0, mut_9_10_63_0, mut_9_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_431
            & and_dcpl_433 & and_dcpl_435 & and_dcpl_437 & and_dcpl_439 & and_dcpl_442
            & and_dcpl_445 & and_dcpl_448 & and_dcpl_451 & and_dcpl_454 & mux_tmp_141));
        rem_13_cmp_4_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_8_2_63_0, mut_8_3_63_0,
            mut_8_4_63_0, mut_8_5_63_0, mut_8_6_63_0, mut_8_7_63_0, mut_8_8_63_0,
            mut_8_9_63_0, mut_8_10_63_0, mut_8_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_431
            & and_dcpl_433 & and_dcpl_435 & and_dcpl_437 & and_dcpl_439 & and_dcpl_442
            & and_dcpl_445 & and_dcpl_448 & and_dcpl_451 & and_dcpl_454 & mux_tmp_141));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1181_cse = '1' ) THEN
        rem_13_cmp_5_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_11_2_63_0, mut_11_3_63_0,
            mut_11_4_63_0, mut_11_5_63_0, mut_11_6_63_0, mut_11_7_63_0, mut_11_8_63_0,
            mut_11_9_63_0, mut_11_10_63_0, mut_11_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_461
            & and_dcpl_465 & and_dcpl_469 & and_dcpl_473 & and_dcpl_477 & and_dcpl_480
            & and_dcpl_483 & and_dcpl_486 & and_dcpl_489 & and_dcpl_492 & and_tmp_125));
        rem_13_cmp_5_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_10_2_63_0, mut_10_3_63_0,
            mut_10_4_63_0, mut_10_5_63_0, mut_10_6_63_0, mut_10_7_63_0, mut_10_8_63_0,
            mut_10_9_63_0, mut_10_10_63_0, mut_10_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_461
            & and_dcpl_465 & and_dcpl_469 & and_dcpl_473 & and_dcpl_477 & and_dcpl_480
            & and_dcpl_483 & and_dcpl_486 & and_dcpl_489 & and_dcpl_492 & and_tmp_125));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1183_cse = '1' ) THEN
        rem_13_cmp_6_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_13_2_63_0, mut_13_3_63_0,
            mut_13_4_63_0, mut_13_5_63_0, mut_13_6_63_0, mut_13_7_63_0, mut_13_8_63_0,
            mut_13_9_63_0, mut_13_10_63_0, mut_13_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_498
            & and_dcpl_500 & and_dcpl_502 & and_dcpl_504 & and_dcpl_506 & and_dcpl_508
            & and_dcpl_510 & and_dcpl_512 & and_dcpl_514 & and_dcpl_516 & mux_tmp_206));
        rem_13_cmp_6_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_12_2_63_0, mut_12_3_63_0,
            mut_12_4_63_0, mut_12_5_63_0, mut_12_6_63_0, mut_12_7_63_0, mut_12_8_63_0,
            mut_12_9_63_0, mut_12_10_63_0, mut_12_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_498
            & and_dcpl_500 & and_dcpl_502 & and_dcpl_504 & and_dcpl_506 & and_dcpl_508
            & and_dcpl_510 & and_dcpl_512 & and_dcpl_514 & and_dcpl_516 & mux_tmp_206));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1185_cse = '1' ) THEN
        rem_13_cmp_7_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_15_2_63_0, mut_15_3_63_0,
            mut_15_4_63_0, mut_15_5_63_0, mut_15_6_63_0, mut_15_7_63_0, mut_15_8_63_0,
            mut_15_9_63_0, mut_15_10_63_0, mut_15_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_520
            & and_dcpl_523 & and_dcpl_526 & and_dcpl_529 & and_dcpl_532 & and_dcpl_534
            & and_dcpl_536 & and_dcpl_538 & and_dcpl_540 & and_dcpl_542 & and_tmp_170));
        rem_13_cmp_7_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_14_2_63_0, mut_14_3_63_0,
            mut_14_4_63_0, mut_14_5_63_0, mut_14_6_63_0, mut_14_7_63_0, mut_14_8_63_0,
            mut_14_9_63_0, mut_14_10_63_0, mut_14_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_520
            & and_dcpl_523 & and_dcpl_526 & and_dcpl_529 & and_dcpl_532 & and_dcpl_534
            & and_dcpl_536 & and_dcpl_538 & and_dcpl_540 & and_dcpl_542 & and_tmp_170));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1187_cse = '1' ) THEN
        rem_13_cmp_8_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_17_2_63_0, mut_17_3_63_0,
            mut_17_4_63_0, mut_17_5_63_0, mut_17_6_63_0, mut_17_7_63_0, mut_17_8_63_0,
            mut_17_9_63_0, mut_17_10_63_0, mut_17_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_546
            & and_dcpl_548 & and_dcpl_550 & and_dcpl_552 & and_dcpl_554 & and_dcpl_556
            & and_dcpl_558 & and_dcpl_560 & and_dcpl_562 & and_dcpl_564 & mux_tmp_271));
        rem_13_cmp_8_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_16_2_63_0, mut_16_3_63_0,
            mut_16_4_63_0, mut_16_5_63_0, mut_16_6_63_0, mut_16_7_63_0, mut_16_8_63_0,
            mut_16_9_63_0, mut_16_10_63_0, mut_16_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_546
            & and_dcpl_548 & and_dcpl_550 & and_dcpl_552 & and_dcpl_554 & and_dcpl_556
            & and_dcpl_558 & and_dcpl_560 & and_dcpl_562 & and_dcpl_564 & mux_tmp_271));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1189_cse = '1' ) THEN
        rem_13_cmp_9_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_19_2_63_0, mut_19_3_63_0,
            mut_19_4_63_0, mut_19_5_63_0, mut_19_6_63_0, mut_19_7_63_0, mut_19_8_63_0,
            mut_19_9_63_0, mut_19_10_63_0, mut_19_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_569
            & and_dcpl_573 & and_dcpl_577 & and_dcpl_581 & and_dcpl_585 & and_dcpl_589
            & and_dcpl_593 & and_dcpl_597 & and_dcpl_601 & and_dcpl_605 & and_tmp_206));
        rem_13_cmp_9_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_18_2_63_0, mut_18_3_63_0,
            mut_18_4_63_0, mut_18_5_63_0, mut_18_6_63_0, mut_18_7_63_0, mut_18_8_63_0,
            mut_18_9_63_0, mut_18_10_63_0, mut_18_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_569
            & and_dcpl_573 & and_dcpl_577 & and_dcpl_581 & and_dcpl_585 & and_dcpl_589
            & and_dcpl_593 & and_dcpl_597 & and_dcpl_601 & and_dcpl_605 & and_tmp_206));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1191_cse = '1' ) THEN
        rem_13_cmp_10_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_21_2_63_0, mut_21_3_63_0,
            mut_21_4_63_0, mut_21_5_63_0, mut_21_6_63_0, mut_21_7_63_0, mut_21_8_63_0,
            mut_21_9_63_0, mut_21_10_63_0, mut_21_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_610
            & and_dcpl_612 & and_dcpl_614 & and_dcpl_616 & and_dcpl_618 & and_dcpl_622
            & and_dcpl_625 & and_dcpl_628 & and_dcpl_631 & and_dcpl_634 & mux_tmp_354));
        rem_13_cmp_10_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_20_2_63_0,
            mut_20_3_63_0, mut_20_4_63_0, mut_20_5_63_0, mut_20_6_63_0, mut_20_7_63_0,
            mut_20_8_63_0, mut_20_9_63_0, mut_20_10_63_0, mut_20_11_63_0, STD_LOGIC_VECTOR'(
            and_dcpl_610 & and_dcpl_612 & and_dcpl_614 & and_dcpl_616 & and_dcpl_618
            & and_dcpl_622 & and_dcpl_625 & and_dcpl_628 & and_dcpl_631 & and_dcpl_634
            & mux_tmp_354));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1193_cse = '1' ) THEN
        rem_13_cmp_11_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_23_2_63_0, mut_23_3_63_0,
            mut_23_4_63_0, mut_23_5_63_0, mut_23_6_63_0, mut_23_7_63_0, mut_23_8_63_0,
            mut_23_9_63_0, mut_23_10_63_0, mut_23_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_638
            & and_dcpl_641 & and_dcpl_644 & and_dcpl_647 & and_dcpl_650 & and_dcpl_653
            & and_dcpl_657 & and_dcpl_661 & and_dcpl_665 & and_dcpl_669 & and_tmp_233));
        rem_13_cmp_11_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_22_2_63_0,
            mut_22_3_63_0, mut_22_4_63_0, mut_22_5_63_0, mut_22_6_63_0, mut_22_7_63_0,
            mut_22_8_63_0, mut_22_9_63_0, mut_22_10_63_0, mut_22_11_63_0, STD_LOGIC_VECTOR'(
            and_dcpl_638 & and_dcpl_641 & and_dcpl_644 & and_dcpl_647 & and_dcpl_650
            & and_dcpl_653 & and_dcpl_657 & and_dcpl_661 & and_dcpl_665 & and_dcpl_669
            & and_tmp_233));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1195_cse = '1' ) THEN
        rem_13_cmp_b_63_0 <= MUX1HOT_v_64_11_2(m_rsci_idat, mut_1_2_63_0, mut_1_3_63_0,
            mut_1_4_63_0, mut_1_5_63_0, mut_1_6_63_0, mut_1_7_63_0, mut_1_8_63_0,
            mut_1_9_63_0, mut_1_10_63_0, mut_1_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_673
            & and_dcpl_675 & and_dcpl_677 & and_dcpl_679 & and_dcpl_681 & and_dcpl_684
            & and_dcpl_687 & and_dcpl_690 & and_dcpl_693 & and_dcpl_696 & mux_tmp_437));
        rem_13_cmp_a_63_0 <= MUX1HOT_v_64_11_2(base_rsci_idat, mut_2_63_0, mut_3_63_0,
            mut_4_63_0, mut_5_63_0, mut_6_63_0, mut_7_63_0, mut_8_63_0, mut_9_63_0,
            mut_10_63_0, mut_11_63_0, STD_LOGIC_VECTOR'( and_dcpl_673 & and_dcpl_675
            & and_dcpl_677 & and_dcpl_679 & and_dcpl_681 & and_dcpl_684 & and_dcpl_687
            & and_dcpl_690 & and_dcpl_693 & and_dcpl_696 & mux_tmp_437));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1205_cse = '1' ) THEN
        mut_3_11_63_0 <= mut_3_10_63_0;
        mut_2_11_63_0 <= mut_2_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1207_cse = '1' ) THEN
        mut_5_11_63_0 <= mut_5_10_63_0;
        mut_4_11_63_0 <= mut_4_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1209_cse = '1' ) THEN
        mut_7_11_63_0 <= mut_7_10_63_0;
        mut_6_11_63_0 <= mut_6_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1211_cse = '1' ) THEN
        mut_9_11_63_0 <= mut_9_10_63_0;
        mut_8_11_63_0 <= mut_8_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1213_cse = '1' ) THEN
        mut_11_11_63_0 <= mut_11_10_63_0;
        mut_10_11_63_0 <= mut_10_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1215_cse = '1' ) THEN
        mut_13_11_63_0 <= mut_13_10_63_0;
        mut_12_11_63_0 <= mut_12_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1217_cse = '1' ) THEN
        mut_15_11_63_0 <= mut_15_10_63_0;
        mut_14_11_63_0 <= mut_14_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1219_cse = '1' ) THEN
        mut_17_11_63_0 <= mut_17_10_63_0;
        mut_16_11_63_0 <= mut_16_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1221_cse = '1' ) THEN
        mut_19_11_63_0 <= mut_19_10_63_0;
        mut_18_11_63_0 <= mut_18_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1223_cse = '1' ) THEN
        mut_21_11_63_0 <= mut_21_10_63_0;
        mut_20_11_63_0 <= mut_20_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1225_cse = '1' ) THEN
        mut_23_11_63_0 <= mut_23_10_63_0;
        mut_22_11_63_0 <= mut_22_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1227_cse = '1' ) THEN
        mut_1_11_63_0 <= mut_1_10_63_0;
        mut_11_63_0 <= mut_10_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_11_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_11_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1229_cse = '1' ) THEN
        rem_12cyc_st_11_3_2 <= rem_12cyc_st_10_3_2;
        rem_12cyc_st_11_1_0 <= rem_12cyc_st_10_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1231_cse = '1' ) THEN
        mut_3_10_63_0 <= mut_3_9_63_0;
        mut_2_10_63_0 <= mut_2_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1233_cse = '1' ) THEN
        mut_5_10_63_0 <= mut_5_9_63_0;
        mut_4_10_63_0 <= mut_4_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1235_cse = '1' ) THEN
        mut_7_10_63_0 <= mut_7_9_63_0;
        mut_6_10_63_0 <= mut_6_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1237_cse = '1' ) THEN
        mut_9_10_63_0 <= mut_9_9_63_0;
        mut_8_10_63_0 <= mut_8_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1239_cse = '1' ) THEN
        mut_11_10_63_0 <= mut_11_9_63_0;
        mut_10_10_63_0 <= mut_10_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1241_cse = '1' ) THEN
        mut_13_10_63_0 <= mut_13_9_63_0;
        mut_12_10_63_0 <= mut_12_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1243_cse = '1' ) THEN
        mut_15_10_63_0 <= mut_15_9_63_0;
        mut_14_10_63_0 <= mut_14_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1245_cse = '1' ) THEN
        mut_17_10_63_0 <= mut_17_9_63_0;
        mut_16_10_63_0 <= mut_16_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1247_cse = '1' ) THEN
        mut_19_10_63_0 <= mut_19_9_63_0;
        mut_18_10_63_0 <= mut_18_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1249_cse = '1' ) THEN
        mut_21_10_63_0 <= mut_21_9_63_0;
        mut_20_10_63_0 <= mut_20_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1251_cse = '1' ) THEN
        mut_23_10_63_0 <= mut_23_9_63_0;
        mut_22_10_63_0 <= mut_22_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1253_cse = '1' ) THEN
        mut_1_10_63_0 <= mut_1_9_63_0;
        mut_10_63_0 <= mut_9_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_10_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_10_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1255_cse = '1' ) THEN
        rem_12cyc_st_10_3_2 <= rem_12cyc_st_9_3_2;
        rem_12cyc_st_10_1_0 <= rem_12cyc_st_9_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1257_cse = '1' ) THEN
        mut_3_9_63_0 <= mut_3_8_63_0;
        mut_2_9_63_0 <= mut_2_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1259_cse = '1' ) THEN
        mut_5_9_63_0 <= mut_5_8_63_0;
        mut_4_9_63_0 <= mut_4_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1261_cse = '1' ) THEN
        mut_7_9_63_0 <= mut_7_8_63_0;
        mut_6_9_63_0 <= mut_6_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1263_cse = '1' ) THEN
        mut_9_9_63_0 <= mut_9_8_63_0;
        mut_8_9_63_0 <= mut_8_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1265_cse = '1' ) THEN
        mut_11_9_63_0 <= mut_11_8_63_0;
        mut_10_9_63_0 <= mut_10_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1267_cse = '1' ) THEN
        mut_13_9_63_0 <= mut_13_8_63_0;
        mut_12_9_63_0 <= mut_12_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1269_cse = '1' ) THEN
        mut_15_9_63_0 <= mut_15_8_63_0;
        mut_14_9_63_0 <= mut_14_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1271_cse = '1' ) THEN
        mut_17_9_63_0 <= mut_17_8_63_0;
        mut_16_9_63_0 <= mut_16_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1273_cse = '1' ) THEN
        mut_19_9_63_0 <= mut_19_8_63_0;
        mut_18_9_63_0 <= mut_18_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1275_cse = '1' ) THEN
        mut_21_9_63_0 <= mut_21_8_63_0;
        mut_20_9_63_0 <= mut_20_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1277_cse = '1' ) THEN
        mut_23_9_63_0 <= mut_23_8_63_0;
        mut_22_9_63_0 <= mut_22_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1279_cse = '1' ) THEN
        mut_1_9_63_0 <= mut_1_8_63_0;
        mut_9_63_0 <= mut_8_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_9_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_9_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1281_cse = '1' ) THEN
        rem_12cyc_st_9_3_2 <= rem_12cyc_st_8_3_2;
        rem_12cyc_st_9_1_0 <= rem_12cyc_st_8_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1283_cse = '1' ) THEN
        mut_3_8_63_0 <= mut_3_7_63_0;
        mut_2_8_63_0 <= mut_2_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1285_cse = '1' ) THEN
        mut_5_8_63_0 <= mut_5_7_63_0;
        mut_4_8_63_0 <= mut_4_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1287_cse = '1' ) THEN
        mut_7_8_63_0 <= mut_7_7_63_0;
        mut_6_8_63_0 <= mut_6_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1289_cse = '1' ) THEN
        mut_9_8_63_0 <= mut_9_7_63_0;
        mut_8_8_63_0 <= mut_8_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1291_cse = '1' ) THEN
        mut_11_8_63_0 <= mut_11_7_63_0;
        mut_10_8_63_0 <= mut_10_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1293_cse = '1' ) THEN
        mut_13_8_63_0 <= mut_13_7_63_0;
        mut_12_8_63_0 <= mut_12_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1295_cse = '1' ) THEN
        mut_15_8_63_0 <= mut_15_7_63_0;
        mut_14_8_63_0 <= mut_14_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1297_cse = '1' ) THEN
        mut_17_8_63_0 <= mut_17_7_63_0;
        mut_16_8_63_0 <= mut_16_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1299_cse = '1' ) THEN
        mut_19_8_63_0 <= mut_19_7_63_0;
        mut_18_8_63_0 <= mut_18_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1301_cse = '1' ) THEN
        mut_21_8_63_0 <= mut_21_7_63_0;
        mut_20_8_63_0 <= mut_20_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1303_cse = '1' ) THEN
        mut_23_8_63_0 <= mut_23_7_63_0;
        mut_22_8_63_0 <= mut_22_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1305_cse = '1' ) THEN
        mut_1_8_63_0 <= mut_1_7_63_0;
        mut_8_63_0 <= mut_7_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_8_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_8_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1307_cse = '1' ) THEN
        rem_12cyc_st_8_3_2 <= rem_12cyc_st_7_3_2;
        rem_12cyc_st_8_1_0 <= rem_12cyc_st_7_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1309_cse = '1' ) THEN
        mut_3_7_63_0 <= mut_3_6_63_0;
        mut_2_7_63_0 <= mut_2_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1311_cse = '1' ) THEN
        mut_5_7_63_0 <= mut_5_6_63_0;
        mut_4_7_63_0 <= mut_4_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1313_cse = '1' ) THEN
        mut_7_7_63_0 <= mut_7_6_63_0;
        mut_6_7_63_0 <= mut_6_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1315_cse = '1' ) THEN
        mut_9_7_63_0 <= mut_9_6_63_0;
        mut_8_7_63_0 <= mut_8_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1317_cse = '1' ) THEN
        mut_11_7_63_0 <= mut_11_6_63_0;
        mut_10_7_63_0 <= mut_10_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1319_cse = '1' ) THEN
        mut_13_7_63_0 <= mut_13_6_63_0;
        mut_12_7_63_0 <= mut_12_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1321_cse = '1' ) THEN
        mut_15_7_63_0 <= mut_15_6_63_0;
        mut_14_7_63_0 <= mut_14_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1323_cse = '1' ) THEN
        mut_17_7_63_0 <= mut_17_6_63_0;
        mut_16_7_63_0 <= mut_16_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1325_cse = '1' ) THEN
        mut_19_7_63_0 <= mut_19_6_63_0;
        mut_18_7_63_0 <= mut_18_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1327_cse = '1' ) THEN
        mut_21_7_63_0 <= mut_21_6_63_0;
        mut_20_7_63_0 <= mut_20_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1329_cse = '1' ) THEN
        mut_23_7_63_0 <= mut_23_6_63_0;
        mut_22_7_63_0 <= mut_22_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1331_cse = '1' ) THEN
        mut_1_7_63_0 <= mut_1_6_63_0;
        mut_7_63_0 <= mut_6_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_7_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_7_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1333_cse = '1' ) THEN
        rem_12cyc_st_7_3_2 <= rem_12cyc_st_6_3_2;
        rem_12cyc_st_7_1_0 <= rem_12cyc_st_6_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1335_cse = '1' ) THEN
        mut_3_6_63_0 <= mut_3_5_63_0;
        mut_2_6_63_0 <= mut_2_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1337_cse = '1' ) THEN
        mut_5_6_63_0 <= mut_5_5_63_0;
        mut_4_6_63_0 <= mut_4_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1339_cse = '1' ) THEN
        mut_7_6_63_0 <= mut_7_5_63_0;
        mut_6_6_63_0 <= mut_6_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1341_cse = '1' ) THEN
        mut_9_6_63_0 <= mut_9_5_63_0;
        mut_8_6_63_0 <= mut_8_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1343_cse = '1' ) THEN
        mut_11_6_63_0 <= mut_11_5_63_0;
        mut_10_6_63_0 <= mut_10_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1345_cse = '1' ) THEN
        mut_13_6_63_0 <= mut_13_5_63_0;
        mut_12_6_63_0 <= mut_12_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1347_cse = '1' ) THEN
        mut_15_6_63_0 <= mut_15_5_63_0;
        mut_14_6_63_0 <= mut_14_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1349_cse = '1' ) THEN
        mut_17_6_63_0 <= mut_17_5_63_0;
        mut_16_6_63_0 <= mut_16_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1351_cse = '1' ) THEN
        mut_19_6_63_0 <= mut_19_5_63_0;
        mut_18_6_63_0 <= mut_18_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1353_cse = '1' ) THEN
        mut_21_6_63_0 <= mut_21_5_63_0;
        mut_20_6_63_0 <= mut_20_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1355_cse = '1' ) THEN
        mut_23_6_63_0 <= mut_23_5_63_0;
        mut_22_6_63_0 <= mut_22_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1357_cse = '1' ) THEN
        mut_1_6_63_0 <= mut_1_5_63_0;
        mut_6_63_0 <= mut_5_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1359_cse = '1' ) THEN
        m_buf_sva_6 <= m_buf_sva_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_6_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_6_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1359_cse = '1' ) THEN
        rem_12cyc_st_6_3_2 <= rem_12cyc_st_5_3_2;
        rem_12cyc_st_6_1_0 <= rem_12cyc_st_5_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1361_cse = '1' ) THEN
        mut_3_5_63_0 <= mut_3_4_63_0;
        mut_2_5_63_0 <= mut_2_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1363_cse = '1' ) THEN
        mut_5_5_63_0 <= mut_5_4_63_0;
        mut_4_5_63_0 <= mut_4_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1365_cse = '1' ) THEN
        mut_7_5_63_0 <= mut_7_4_63_0;
        mut_6_5_63_0 <= mut_6_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1367_cse = '1' ) THEN
        mut_9_5_63_0 <= mut_9_4_63_0;
        mut_8_5_63_0 <= mut_8_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1369_cse = '1' ) THEN
        mut_11_5_63_0 <= mut_11_4_63_0;
        mut_10_5_63_0 <= mut_10_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1371_cse = '1' ) THEN
        mut_13_5_63_0 <= mut_13_4_63_0;
        mut_12_5_63_0 <= mut_12_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1373_cse = '1' ) THEN
        mut_15_5_63_0 <= mut_15_4_63_0;
        mut_14_5_63_0 <= mut_14_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1375_cse = '1' ) THEN
        mut_17_5_63_0 <= mut_17_4_63_0;
        mut_16_5_63_0 <= mut_16_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1377_cse = '1' ) THEN
        mut_19_5_63_0 <= mut_19_4_63_0;
        mut_18_5_63_0 <= mut_18_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1379_cse = '1' ) THEN
        mut_21_5_63_0 <= mut_21_4_63_0;
        mut_20_5_63_0 <= mut_20_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1381_cse = '1' ) THEN
        mut_23_5_63_0 <= mut_23_4_63_0;
        mut_22_5_63_0 <= mut_22_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1383_cse = '1' ) THEN
        mut_1_5_63_0 <= mut_1_4_63_0;
        mut_5_63_0 <= mut_4_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1385_cse = '1' ) THEN
        m_buf_sva_5 <= m_buf_sva_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_5_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_5_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1385_cse = '1' ) THEN
        rem_12cyc_st_5_3_2 <= rem_12cyc_st_4_3_2;
        rem_12cyc_st_5_1_0 <= rem_12cyc_st_4_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1387_cse = '1' ) THEN
        mut_3_4_63_0 <= mut_3_3_63_0;
        mut_2_4_63_0 <= mut_2_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1389_cse = '1' ) THEN
        mut_5_4_63_0 <= mut_5_3_63_0;
        mut_4_4_63_0 <= mut_4_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1391_cse = '1' ) THEN
        mut_7_4_63_0 <= mut_7_3_63_0;
        mut_6_4_63_0 <= mut_6_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1393_cse = '1' ) THEN
        mut_9_4_63_0 <= mut_9_3_63_0;
        mut_8_4_63_0 <= mut_8_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1395_cse = '1' ) THEN
        mut_11_4_63_0 <= mut_11_3_63_0;
        mut_10_4_63_0 <= mut_10_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1397_cse = '1' ) THEN
        mut_13_4_63_0 <= mut_13_3_63_0;
        mut_12_4_63_0 <= mut_12_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1399_cse = '1' ) THEN
        mut_15_4_63_0 <= mut_15_3_63_0;
        mut_14_4_63_0 <= mut_14_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1401_cse = '1' ) THEN
        mut_17_4_63_0 <= mut_17_3_63_0;
        mut_16_4_63_0 <= mut_16_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1403_cse = '1' ) THEN
        mut_19_4_63_0 <= mut_19_3_63_0;
        mut_18_4_63_0 <= mut_18_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1405_cse = '1' ) THEN
        mut_21_4_63_0 <= mut_21_3_63_0;
        mut_20_4_63_0 <= mut_20_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1407_cse = '1' ) THEN
        mut_23_4_63_0 <= mut_23_3_63_0;
        mut_22_4_63_0 <= mut_22_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1409_cse = '1' ) THEN
        mut_1_4_63_0 <= mut_1_3_63_0;
        mut_4_63_0 <= mut_3_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1411_cse = '1' ) THEN
        m_buf_sva_4 <= m_buf_sva_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_4_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_4_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1411_cse = '1' ) THEN
        rem_12cyc_st_4_3_2 <= rem_12cyc_st_3_3_2;
        rem_12cyc_st_4_1_0 <= rem_12cyc_st_3_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1413_cse = '1' ) THEN
        mut_3_3_63_0 <= mut_3_2_63_0;
        mut_2_3_63_0 <= mut_2_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1415_cse = '1' ) THEN
        mut_5_3_63_0 <= mut_5_2_63_0;
        mut_4_3_63_0 <= mut_4_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1417_cse = '1' ) THEN
        mut_7_3_63_0 <= mut_7_2_63_0;
        mut_6_3_63_0 <= mut_6_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1419_cse = '1' ) THEN
        mut_9_3_63_0 <= mut_9_2_63_0;
        mut_8_3_63_0 <= mut_8_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1421_cse = '1' ) THEN
        mut_11_3_63_0 <= mut_11_2_63_0;
        mut_10_3_63_0 <= mut_10_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1423_cse = '1' ) THEN
        mut_13_3_63_0 <= mut_13_2_63_0;
        mut_12_3_63_0 <= mut_12_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1425_cse = '1' ) THEN
        mut_15_3_63_0 <= mut_15_2_63_0;
        mut_14_3_63_0 <= mut_14_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1427_cse = '1' ) THEN
        mut_17_3_63_0 <= mut_17_2_63_0;
        mut_16_3_63_0 <= mut_16_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1429_cse = '1' ) THEN
        mut_19_3_63_0 <= mut_19_2_63_0;
        mut_18_3_63_0 <= mut_18_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1431_cse = '1' ) THEN
        mut_21_3_63_0 <= mut_21_2_63_0;
        mut_20_3_63_0 <= mut_20_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1433_cse = '1' ) THEN
        mut_23_3_63_0 <= mut_23_2_63_0;
        mut_22_3_63_0 <= mut_22_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1435_cse = '1' ) THEN
        mut_1_3_63_0 <= mut_1_2_63_0;
        mut_3_63_0 <= mut_2_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1437_cse = '1' ) THEN
        m_buf_sva_3 <= m_buf_sva_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_3_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_3_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1437_cse = '1' ) THEN
        rem_12cyc_st_3_3_2 <= rem_12cyc_st_2_3_2;
        rem_12cyc_st_3_1_0 <= rem_12cyc_st_2_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1439_cse = '1' ) THEN
        mut_3_2_63_0 <= rem_13_cmp_1_b_63_0;
        mut_2_2_63_0 <= rem_13_cmp_1_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1441_cse = '1' ) THEN
        mut_5_2_63_0 <= rem_13_cmp_2_b_63_0;
        mut_4_2_63_0 <= rem_13_cmp_2_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1443_cse = '1' ) THEN
        mut_7_2_63_0 <= rem_13_cmp_3_b_63_0;
        mut_6_2_63_0 <= rem_13_cmp_3_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1445_cse = '1' ) THEN
        mut_9_2_63_0 <= rem_13_cmp_4_b_63_0;
        mut_8_2_63_0 <= rem_13_cmp_4_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1447_cse = '1' ) THEN
        mut_11_2_63_0 <= rem_13_cmp_5_b_63_0;
        mut_10_2_63_0 <= rem_13_cmp_5_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1449_cse = '1' ) THEN
        mut_13_2_63_0 <= rem_13_cmp_6_b_63_0;
        mut_12_2_63_0 <= rem_13_cmp_6_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1451_cse = '1' ) THEN
        mut_15_2_63_0 <= rem_13_cmp_7_b_63_0;
        mut_14_2_63_0 <= rem_13_cmp_7_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1453_cse = '1' ) THEN
        mut_17_2_63_0 <= rem_13_cmp_8_b_63_0;
        mut_16_2_63_0 <= rem_13_cmp_8_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1455_cse = '1' ) THEN
        mut_19_2_63_0 <= rem_13_cmp_9_b_63_0;
        mut_18_2_63_0 <= rem_13_cmp_9_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1457_cse = '1' ) THEN
        mut_21_2_63_0 <= rem_13_cmp_10_b_63_0;
        mut_20_2_63_0 <= rem_13_cmp_10_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1459_cse = '1' ) THEN
        mut_23_2_63_0 <= rem_13_cmp_11_b_63_0;
        mut_22_2_63_0 <= rem_13_cmp_11_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1461_cse = '1' ) THEN
        mut_1_2_63_0 <= rem_13_cmp_b_63_0;
        mut_2_63_0 <= rem_13_cmp_a_63_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1463_cse = '1' ) THEN
        m_buf_sva_2 <= m_buf_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_st_2_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_st_2_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1463_cse = '1' ) THEN
        rem_12cyc_st_2_3_2 <= rem_12cyc_3_2;
        rem_12cyc_st_2_1_0 <= rem_12cyc_1_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF ( and_1197_cse = '1' ) THEN
        m_buf_sva_1 <= m_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (ccs_ccore_clk)
  BEGIN
    IF ccs_ccore_clk'EVENT AND ( ccs_ccore_clk = '1' ) THEN
      IF (ccs_ccore_srst = '1') THEN
        rem_12cyc_3_2 <= STD_LOGIC_VECTOR'( "00");
        rem_12cyc_1_0 <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( and_1197_cse = '1' ) THEN
        rem_12cyc_3_2 <= acc_tmp;
        rem_12cyc_1_0 <= acc_1_tmp(1 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  qelse_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(result_sva_duc_mx0) + UNSIGNED(m_buf_sva_12),
      64));
  mux_10_nl <= MUX_s_1_2_2((rem_13_cmp_1_z(63)), (rem_13_cmp_3_z(63)), rem_12cyc_st_12_1_0(1));
  mux_9_nl <= MUX_s_1_2_2((rem_13_cmp_2_z(63)), (rem_13_cmp_4_z(63)), rem_12cyc_st_12_1_0(1));
  mux_11_nl <= MUX_s_1_2_2(mux_10_nl, mux_9_nl, rem_12cyc_st_12_1_0(0));
  mux_7_nl <= MUX_s_1_2_2((rem_13_cmp_9_z(63)), (rem_13_cmp_11_z(63)), rem_12cyc_st_12_1_0(1));
  mux_6_nl <= MUX_s_1_2_2((rem_13_cmp_10_z(63)), (rem_13_cmp_z(63)), rem_12cyc_st_12_1_0(1));
  mux_8_nl <= MUX_s_1_2_2(mux_7_nl, mux_6_nl, rem_12cyc_st_12_1_0(0));
  mux_12_nl <= MUX_s_1_2_2(mux_11_nl, mux_8_nl, rem_12cyc_st_12_3_2(1));
  mux_3_nl <= MUX_s_1_2_2((rem_13_cmp_5_z(63)), (rem_13_cmp_7_z(63)), rem_12cyc_st_12_1_0(1));
  mux_2_nl <= MUX_s_1_2_2((rem_13_cmp_6_z(63)), (rem_13_cmp_8_z(63)), rem_12cyc_st_12_1_0(1));
  mux_4_nl <= MUX_s_1_2_2(mux_3_nl, mux_2_nl, rem_12cyc_st_12_1_0(0));
  mux_5_nl <= MUX_s_1_2_2(mux_4_nl, (result_sva_duc(63)), rem_12cyc_st_12_3_2(1));
  mux_13_nl <= MUX_s_1_2_2(mux_12_nl, mux_5_nl, rem_12cyc_st_12_3_2(0));
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    modulo_dev
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_out_dreg_pkg_v2.ALL;
USE work.mgc_comps.ALL;


ENTITY modulo_dev IS
  PORT(
    base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    ccs_ccore_start_rsc_dat : IN STD_LOGIC;
    ccs_ccore_clk : IN STD_LOGIC;
    ccs_ccore_srst : IN STD_LOGIC;
    ccs_ccore_en : IN STD_LOGIC
  );
END modulo_dev;

ARCHITECTURE v1 OF modulo_dev IS
  -- Default Constants

  COMPONENT modulo_dev_core
    PORT(
      base_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_dev_core_inst_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_core_inst_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_core_inst_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  modulo_dev_core_inst : modulo_dev_core
    PORT MAP(
      base_rsc_dat => modulo_dev_core_inst_base_rsc_dat,
      m_rsc_dat => modulo_dev_core_inst_m_rsc_dat,
      return_rsc_z => modulo_dev_core_inst_return_rsc_z,
      ccs_ccore_start_rsc_dat => ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => ccs_ccore_clk,
      ccs_ccore_srst => ccs_ccore_srst,
      ccs_ccore_en => ccs_ccore_en
    );
  modulo_dev_core_inst_base_rsc_dat <= base_rsc_dat;
  modulo_dev_core_inst_m_rsc_dat <= m_rsc_dat;
  return_rsc_z <= modulo_dev_core_inst_return_rsc_z;

END v1;




--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_div IS
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END mgc_div;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

USE work.funcs.all;

ARCHITECTURE beh OF mgc_div IS
BEGIN
  z <= std_logic_vector(unsigned(a) / unsigned(b)) WHEN signd = 0 ELSE
       std_logic_vector(  signed(a) /   signed(b));
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   yl7897@newnano.poly.edu
--  Generated date: Thu Aug  5 01:55:06 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen;

ARCHITECTURE v11 OF inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen
    IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    STAGE_LOOP_C_3_tr0 : IN STD_LOGIC;
    modExp_dev_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_1_tr0 : IN STD_LOGIC;
    COMP_LOOP_1_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_32_tr0 : IN STD_LOGIC;
    COMP_LOOP_2_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_64_tr0 : IN STD_LOGIC;
    COMP_LOOP_3_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_96_tr0 : IN STD_LOGIC;
    COMP_LOOP_4_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_128_tr0 : IN STD_LOGIC;
    COMP_LOOP_5_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_160_tr0 : IN STD_LOGIC;
    COMP_LOOP_6_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_192_tr0 : IN STD_LOGIC;
    COMP_LOOP_7_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_224_tr0 : IN STD_LOGIC;
    COMP_LOOP_8_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_256_tr0 : IN STD_LOGIC;
    COMP_LOOP_9_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_288_tr0 : IN STD_LOGIC;
    COMP_LOOP_10_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_320_tr0 : IN STD_LOGIC;
    COMP_LOOP_11_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_352_tr0 : IN STD_LOGIC;
    COMP_LOOP_12_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_384_tr0 : IN STD_LOGIC;
    COMP_LOOP_13_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_416_tr0 : IN STD_LOGIC;
    COMP_LOOP_14_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_448_tr0 : IN STD_LOGIC;
    COMP_LOOP_15_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_480_tr0 : IN STD_LOGIC;
    COMP_LOOP_16_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
    COMP_LOOP_C_512_tr0 : IN STD_LOGIC;
    VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
    STAGE_LOOP_C_4_tr0 : IN STD_LOGIC
  );
END inPlaceNTT_DIT_core_core_fsm;

ARCHITECTURE v11 OF inPlaceNTT_DIT_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  TYPE inPlaceNTT_DIT_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, STAGE_LOOP_C_1,
      STAGE_LOOP_C_2, STAGE_LOOP_C_3, modExp_dev_while_C_0, modExp_dev_while_C_1,
      modExp_dev_while_C_2, modExp_dev_while_C_3, modExp_dev_while_C_4, modExp_dev_while_C_5,
      modExp_dev_while_C_6, modExp_dev_while_C_7, modExp_dev_while_C_8, modExp_dev_while_C_9,
      modExp_dev_while_C_10, modExp_dev_while_C_11, modExp_dev_while_C_12, modExp_dev_while_C_13,
      modExp_dev_while_C_14, COMP_LOOP_C_0, COMP_LOOP_C_1, COMP_LOOP_1_modExp_dev_1_while_C_0,
      COMP_LOOP_1_modExp_dev_1_while_C_1, COMP_LOOP_1_modExp_dev_1_while_C_2, COMP_LOOP_1_modExp_dev_1_while_C_3,
      COMP_LOOP_1_modExp_dev_1_while_C_4, COMP_LOOP_1_modExp_dev_1_while_C_5, COMP_LOOP_1_modExp_dev_1_while_C_6,
      COMP_LOOP_1_modExp_dev_1_while_C_7, COMP_LOOP_1_modExp_dev_1_while_C_8, COMP_LOOP_1_modExp_dev_1_while_C_9,
      COMP_LOOP_1_modExp_dev_1_while_C_10, COMP_LOOP_1_modExp_dev_1_while_C_11, COMP_LOOP_1_modExp_dev_1_while_C_12,
      COMP_LOOP_1_modExp_dev_1_while_C_13, COMP_LOOP_1_modExp_dev_1_while_C_14, COMP_LOOP_C_2,
      COMP_LOOP_C_3, COMP_LOOP_C_4, COMP_LOOP_C_5, COMP_LOOP_C_6, COMP_LOOP_C_7,
      COMP_LOOP_C_8, COMP_LOOP_C_9, COMP_LOOP_C_10, COMP_LOOP_C_11, COMP_LOOP_C_12,
      COMP_LOOP_C_13, COMP_LOOP_C_14, COMP_LOOP_C_15, COMP_LOOP_C_16, COMP_LOOP_C_17,
      COMP_LOOP_C_18, COMP_LOOP_C_19, COMP_LOOP_C_20, COMP_LOOP_C_21, COMP_LOOP_C_22,
      COMP_LOOP_C_23, COMP_LOOP_C_24, COMP_LOOP_C_25, COMP_LOOP_C_26, COMP_LOOP_C_27,
      COMP_LOOP_C_28, COMP_LOOP_C_29, COMP_LOOP_C_30, COMP_LOOP_C_31, COMP_LOOP_C_32,
      COMP_LOOP_C_33, COMP_LOOP_2_modExp_dev_1_while_C_0, COMP_LOOP_2_modExp_dev_1_while_C_1,
      COMP_LOOP_2_modExp_dev_1_while_C_2, COMP_LOOP_2_modExp_dev_1_while_C_3, COMP_LOOP_2_modExp_dev_1_while_C_4,
      COMP_LOOP_2_modExp_dev_1_while_C_5, COMP_LOOP_2_modExp_dev_1_while_C_6, COMP_LOOP_2_modExp_dev_1_while_C_7,
      COMP_LOOP_2_modExp_dev_1_while_C_8, COMP_LOOP_2_modExp_dev_1_while_C_9, COMP_LOOP_2_modExp_dev_1_while_C_10,
      COMP_LOOP_2_modExp_dev_1_while_C_11, COMP_LOOP_2_modExp_dev_1_while_C_12, COMP_LOOP_2_modExp_dev_1_while_C_13,
      COMP_LOOP_2_modExp_dev_1_while_C_14, COMP_LOOP_C_34, COMP_LOOP_C_35, COMP_LOOP_C_36,
      COMP_LOOP_C_37, COMP_LOOP_C_38, COMP_LOOP_C_39, COMP_LOOP_C_40, COMP_LOOP_C_41,
      COMP_LOOP_C_42, COMP_LOOP_C_43, COMP_LOOP_C_44, COMP_LOOP_C_45, COMP_LOOP_C_46,
      COMP_LOOP_C_47, COMP_LOOP_C_48, COMP_LOOP_C_49, COMP_LOOP_C_50, COMP_LOOP_C_51,
      COMP_LOOP_C_52, COMP_LOOP_C_53, COMP_LOOP_C_54, COMP_LOOP_C_55, COMP_LOOP_C_56,
      COMP_LOOP_C_57, COMP_LOOP_C_58, COMP_LOOP_C_59, COMP_LOOP_C_60, COMP_LOOP_C_61,
      COMP_LOOP_C_62, COMP_LOOP_C_63, COMP_LOOP_C_64, COMP_LOOP_C_65, COMP_LOOP_3_modExp_dev_1_while_C_0,
      COMP_LOOP_3_modExp_dev_1_while_C_1, COMP_LOOP_3_modExp_dev_1_while_C_2, COMP_LOOP_3_modExp_dev_1_while_C_3,
      COMP_LOOP_3_modExp_dev_1_while_C_4, COMP_LOOP_3_modExp_dev_1_while_C_5, COMP_LOOP_3_modExp_dev_1_while_C_6,
      COMP_LOOP_3_modExp_dev_1_while_C_7, COMP_LOOP_3_modExp_dev_1_while_C_8, COMP_LOOP_3_modExp_dev_1_while_C_9,
      COMP_LOOP_3_modExp_dev_1_while_C_10, COMP_LOOP_3_modExp_dev_1_while_C_11, COMP_LOOP_3_modExp_dev_1_while_C_12,
      COMP_LOOP_3_modExp_dev_1_while_C_13, COMP_LOOP_3_modExp_dev_1_while_C_14, COMP_LOOP_C_66,
      COMP_LOOP_C_67, COMP_LOOP_C_68, COMP_LOOP_C_69, COMP_LOOP_C_70, COMP_LOOP_C_71,
      COMP_LOOP_C_72, COMP_LOOP_C_73, COMP_LOOP_C_74, COMP_LOOP_C_75, COMP_LOOP_C_76,
      COMP_LOOP_C_77, COMP_LOOP_C_78, COMP_LOOP_C_79, COMP_LOOP_C_80, COMP_LOOP_C_81,
      COMP_LOOP_C_82, COMP_LOOP_C_83, COMP_LOOP_C_84, COMP_LOOP_C_85, COMP_LOOP_C_86,
      COMP_LOOP_C_87, COMP_LOOP_C_88, COMP_LOOP_C_89, COMP_LOOP_C_90, COMP_LOOP_C_91,
      COMP_LOOP_C_92, COMP_LOOP_C_93, COMP_LOOP_C_94, COMP_LOOP_C_95, COMP_LOOP_C_96,
      COMP_LOOP_C_97, COMP_LOOP_4_modExp_dev_1_while_C_0, COMP_LOOP_4_modExp_dev_1_while_C_1,
      COMP_LOOP_4_modExp_dev_1_while_C_2, COMP_LOOP_4_modExp_dev_1_while_C_3, COMP_LOOP_4_modExp_dev_1_while_C_4,
      COMP_LOOP_4_modExp_dev_1_while_C_5, COMP_LOOP_4_modExp_dev_1_while_C_6, COMP_LOOP_4_modExp_dev_1_while_C_7,
      COMP_LOOP_4_modExp_dev_1_while_C_8, COMP_LOOP_4_modExp_dev_1_while_C_9, COMP_LOOP_4_modExp_dev_1_while_C_10,
      COMP_LOOP_4_modExp_dev_1_while_C_11, COMP_LOOP_4_modExp_dev_1_while_C_12, COMP_LOOP_4_modExp_dev_1_while_C_13,
      COMP_LOOP_4_modExp_dev_1_while_C_14, COMP_LOOP_C_98, COMP_LOOP_C_99, COMP_LOOP_C_100,
      COMP_LOOP_C_101, COMP_LOOP_C_102, COMP_LOOP_C_103, COMP_LOOP_C_104, COMP_LOOP_C_105,
      COMP_LOOP_C_106, COMP_LOOP_C_107, COMP_LOOP_C_108, COMP_LOOP_C_109, COMP_LOOP_C_110,
      COMP_LOOP_C_111, COMP_LOOP_C_112, COMP_LOOP_C_113, COMP_LOOP_C_114, COMP_LOOP_C_115,
      COMP_LOOP_C_116, COMP_LOOP_C_117, COMP_LOOP_C_118, COMP_LOOP_C_119, COMP_LOOP_C_120,
      COMP_LOOP_C_121, COMP_LOOP_C_122, COMP_LOOP_C_123, COMP_LOOP_C_124, COMP_LOOP_C_125,
      COMP_LOOP_C_126, COMP_LOOP_C_127, COMP_LOOP_C_128, COMP_LOOP_C_129, COMP_LOOP_5_modExp_dev_1_while_C_0,
      COMP_LOOP_5_modExp_dev_1_while_C_1, COMP_LOOP_5_modExp_dev_1_while_C_2, COMP_LOOP_5_modExp_dev_1_while_C_3,
      COMP_LOOP_5_modExp_dev_1_while_C_4, COMP_LOOP_5_modExp_dev_1_while_C_5, COMP_LOOP_5_modExp_dev_1_while_C_6,
      COMP_LOOP_5_modExp_dev_1_while_C_7, COMP_LOOP_5_modExp_dev_1_while_C_8, COMP_LOOP_5_modExp_dev_1_while_C_9,
      COMP_LOOP_5_modExp_dev_1_while_C_10, COMP_LOOP_5_modExp_dev_1_while_C_11, COMP_LOOP_5_modExp_dev_1_while_C_12,
      COMP_LOOP_5_modExp_dev_1_while_C_13, COMP_LOOP_5_modExp_dev_1_while_C_14, COMP_LOOP_C_130,
      COMP_LOOP_C_131, COMP_LOOP_C_132, COMP_LOOP_C_133, COMP_LOOP_C_134, COMP_LOOP_C_135,
      COMP_LOOP_C_136, COMP_LOOP_C_137, COMP_LOOP_C_138, COMP_LOOP_C_139, COMP_LOOP_C_140,
      COMP_LOOP_C_141, COMP_LOOP_C_142, COMP_LOOP_C_143, COMP_LOOP_C_144, COMP_LOOP_C_145,
      COMP_LOOP_C_146, COMP_LOOP_C_147, COMP_LOOP_C_148, COMP_LOOP_C_149, COMP_LOOP_C_150,
      COMP_LOOP_C_151, COMP_LOOP_C_152, COMP_LOOP_C_153, COMP_LOOP_C_154, COMP_LOOP_C_155,
      COMP_LOOP_C_156, COMP_LOOP_C_157, COMP_LOOP_C_158, COMP_LOOP_C_159, COMP_LOOP_C_160,
      COMP_LOOP_C_161, COMP_LOOP_6_modExp_dev_1_while_C_0, COMP_LOOP_6_modExp_dev_1_while_C_1,
      COMP_LOOP_6_modExp_dev_1_while_C_2, COMP_LOOP_6_modExp_dev_1_while_C_3, COMP_LOOP_6_modExp_dev_1_while_C_4,
      COMP_LOOP_6_modExp_dev_1_while_C_5, COMP_LOOP_6_modExp_dev_1_while_C_6, COMP_LOOP_6_modExp_dev_1_while_C_7,
      COMP_LOOP_6_modExp_dev_1_while_C_8, COMP_LOOP_6_modExp_dev_1_while_C_9, COMP_LOOP_6_modExp_dev_1_while_C_10,
      COMP_LOOP_6_modExp_dev_1_while_C_11, COMP_LOOP_6_modExp_dev_1_while_C_12, COMP_LOOP_6_modExp_dev_1_while_C_13,
      COMP_LOOP_6_modExp_dev_1_while_C_14, COMP_LOOP_C_162, COMP_LOOP_C_163, COMP_LOOP_C_164,
      COMP_LOOP_C_165, COMP_LOOP_C_166, COMP_LOOP_C_167, COMP_LOOP_C_168, COMP_LOOP_C_169,
      COMP_LOOP_C_170, COMP_LOOP_C_171, COMP_LOOP_C_172, COMP_LOOP_C_173, COMP_LOOP_C_174,
      COMP_LOOP_C_175, COMP_LOOP_C_176, COMP_LOOP_C_177, COMP_LOOP_C_178, COMP_LOOP_C_179,
      COMP_LOOP_C_180, COMP_LOOP_C_181, COMP_LOOP_C_182, COMP_LOOP_C_183, COMP_LOOP_C_184,
      COMP_LOOP_C_185, COMP_LOOP_C_186, COMP_LOOP_C_187, COMP_LOOP_C_188, COMP_LOOP_C_189,
      COMP_LOOP_C_190, COMP_LOOP_C_191, COMP_LOOP_C_192, COMP_LOOP_C_193, COMP_LOOP_7_modExp_dev_1_while_C_0,
      COMP_LOOP_7_modExp_dev_1_while_C_1, COMP_LOOP_7_modExp_dev_1_while_C_2, COMP_LOOP_7_modExp_dev_1_while_C_3,
      COMP_LOOP_7_modExp_dev_1_while_C_4, COMP_LOOP_7_modExp_dev_1_while_C_5, COMP_LOOP_7_modExp_dev_1_while_C_6,
      COMP_LOOP_7_modExp_dev_1_while_C_7, COMP_LOOP_7_modExp_dev_1_while_C_8, COMP_LOOP_7_modExp_dev_1_while_C_9,
      COMP_LOOP_7_modExp_dev_1_while_C_10, COMP_LOOP_7_modExp_dev_1_while_C_11, COMP_LOOP_7_modExp_dev_1_while_C_12,
      COMP_LOOP_7_modExp_dev_1_while_C_13, COMP_LOOP_7_modExp_dev_1_while_C_14, COMP_LOOP_C_194,
      COMP_LOOP_C_195, COMP_LOOP_C_196, COMP_LOOP_C_197, COMP_LOOP_C_198, COMP_LOOP_C_199,
      COMP_LOOP_C_200, COMP_LOOP_C_201, COMP_LOOP_C_202, COMP_LOOP_C_203, COMP_LOOP_C_204,
      COMP_LOOP_C_205, COMP_LOOP_C_206, COMP_LOOP_C_207, COMP_LOOP_C_208, COMP_LOOP_C_209,
      COMP_LOOP_C_210, COMP_LOOP_C_211, COMP_LOOP_C_212, COMP_LOOP_C_213, COMP_LOOP_C_214,
      COMP_LOOP_C_215, COMP_LOOP_C_216, COMP_LOOP_C_217, COMP_LOOP_C_218, COMP_LOOP_C_219,
      COMP_LOOP_C_220, COMP_LOOP_C_221, COMP_LOOP_C_222, COMP_LOOP_C_223, COMP_LOOP_C_224,
      COMP_LOOP_C_225, COMP_LOOP_8_modExp_dev_1_while_C_0, COMP_LOOP_8_modExp_dev_1_while_C_1,
      COMP_LOOP_8_modExp_dev_1_while_C_2, COMP_LOOP_8_modExp_dev_1_while_C_3, COMP_LOOP_8_modExp_dev_1_while_C_4,
      COMP_LOOP_8_modExp_dev_1_while_C_5, COMP_LOOP_8_modExp_dev_1_while_C_6, COMP_LOOP_8_modExp_dev_1_while_C_7,
      COMP_LOOP_8_modExp_dev_1_while_C_8, COMP_LOOP_8_modExp_dev_1_while_C_9, COMP_LOOP_8_modExp_dev_1_while_C_10,
      COMP_LOOP_8_modExp_dev_1_while_C_11, COMP_LOOP_8_modExp_dev_1_while_C_12, COMP_LOOP_8_modExp_dev_1_while_C_13,
      COMP_LOOP_8_modExp_dev_1_while_C_14, COMP_LOOP_C_226, COMP_LOOP_C_227, COMP_LOOP_C_228,
      COMP_LOOP_C_229, COMP_LOOP_C_230, COMP_LOOP_C_231, COMP_LOOP_C_232, COMP_LOOP_C_233,
      COMP_LOOP_C_234, COMP_LOOP_C_235, COMP_LOOP_C_236, COMP_LOOP_C_237, COMP_LOOP_C_238,
      COMP_LOOP_C_239, COMP_LOOP_C_240, COMP_LOOP_C_241, COMP_LOOP_C_242, COMP_LOOP_C_243,
      COMP_LOOP_C_244, COMP_LOOP_C_245, COMP_LOOP_C_246, COMP_LOOP_C_247, COMP_LOOP_C_248,
      COMP_LOOP_C_249, COMP_LOOP_C_250, COMP_LOOP_C_251, COMP_LOOP_C_252, COMP_LOOP_C_253,
      COMP_LOOP_C_254, COMP_LOOP_C_255, COMP_LOOP_C_256, COMP_LOOP_C_257, COMP_LOOP_9_modExp_dev_1_while_C_0,
      COMP_LOOP_9_modExp_dev_1_while_C_1, COMP_LOOP_9_modExp_dev_1_while_C_2, COMP_LOOP_9_modExp_dev_1_while_C_3,
      COMP_LOOP_9_modExp_dev_1_while_C_4, COMP_LOOP_9_modExp_dev_1_while_C_5, COMP_LOOP_9_modExp_dev_1_while_C_6,
      COMP_LOOP_9_modExp_dev_1_while_C_7, COMP_LOOP_9_modExp_dev_1_while_C_8, COMP_LOOP_9_modExp_dev_1_while_C_9,
      COMP_LOOP_9_modExp_dev_1_while_C_10, COMP_LOOP_9_modExp_dev_1_while_C_11, COMP_LOOP_9_modExp_dev_1_while_C_12,
      COMP_LOOP_9_modExp_dev_1_while_C_13, COMP_LOOP_9_modExp_dev_1_while_C_14, COMP_LOOP_C_258,
      COMP_LOOP_C_259, COMP_LOOP_C_260, COMP_LOOP_C_261, COMP_LOOP_C_262, COMP_LOOP_C_263,
      COMP_LOOP_C_264, COMP_LOOP_C_265, COMP_LOOP_C_266, COMP_LOOP_C_267, COMP_LOOP_C_268,
      COMP_LOOP_C_269, COMP_LOOP_C_270, COMP_LOOP_C_271, COMP_LOOP_C_272, COMP_LOOP_C_273,
      COMP_LOOP_C_274, COMP_LOOP_C_275, COMP_LOOP_C_276, COMP_LOOP_C_277, COMP_LOOP_C_278,
      COMP_LOOP_C_279, COMP_LOOP_C_280, COMP_LOOP_C_281, COMP_LOOP_C_282, COMP_LOOP_C_283,
      COMP_LOOP_C_284, COMP_LOOP_C_285, COMP_LOOP_C_286, COMP_LOOP_C_287, COMP_LOOP_C_288,
      COMP_LOOP_C_289, COMP_LOOP_10_modExp_dev_1_while_C_0, COMP_LOOP_10_modExp_dev_1_while_C_1,
      COMP_LOOP_10_modExp_dev_1_while_C_2, COMP_LOOP_10_modExp_dev_1_while_C_3, COMP_LOOP_10_modExp_dev_1_while_C_4,
      COMP_LOOP_10_modExp_dev_1_while_C_5, COMP_LOOP_10_modExp_dev_1_while_C_6, COMP_LOOP_10_modExp_dev_1_while_C_7,
      COMP_LOOP_10_modExp_dev_1_while_C_8, COMP_LOOP_10_modExp_dev_1_while_C_9, COMP_LOOP_10_modExp_dev_1_while_C_10,
      COMP_LOOP_10_modExp_dev_1_while_C_11, COMP_LOOP_10_modExp_dev_1_while_C_12,
      COMP_LOOP_10_modExp_dev_1_while_C_13, COMP_LOOP_10_modExp_dev_1_while_C_14,
      COMP_LOOP_C_290, COMP_LOOP_C_291, COMP_LOOP_C_292, COMP_LOOP_C_293, COMP_LOOP_C_294,
      COMP_LOOP_C_295, COMP_LOOP_C_296, COMP_LOOP_C_297, COMP_LOOP_C_298, COMP_LOOP_C_299,
      COMP_LOOP_C_300, COMP_LOOP_C_301, COMP_LOOP_C_302, COMP_LOOP_C_303, COMP_LOOP_C_304,
      COMP_LOOP_C_305, COMP_LOOP_C_306, COMP_LOOP_C_307, COMP_LOOP_C_308, COMP_LOOP_C_309,
      COMP_LOOP_C_310, COMP_LOOP_C_311, COMP_LOOP_C_312, COMP_LOOP_C_313, COMP_LOOP_C_314,
      COMP_LOOP_C_315, COMP_LOOP_C_316, COMP_LOOP_C_317, COMP_LOOP_C_318, COMP_LOOP_C_319,
      COMP_LOOP_C_320, COMP_LOOP_C_321, COMP_LOOP_11_modExp_dev_1_while_C_0, COMP_LOOP_11_modExp_dev_1_while_C_1,
      COMP_LOOP_11_modExp_dev_1_while_C_2, COMP_LOOP_11_modExp_dev_1_while_C_3, COMP_LOOP_11_modExp_dev_1_while_C_4,
      COMP_LOOP_11_modExp_dev_1_while_C_5, COMP_LOOP_11_modExp_dev_1_while_C_6, COMP_LOOP_11_modExp_dev_1_while_C_7,
      COMP_LOOP_11_modExp_dev_1_while_C_8, COMP_LOOP_11_modExp_dev_1_while_C_9, COMP_LOOP_11_modExp_dev_1_while_C_10,
      COMP_LOOP_11_modExp_dev_1_while_C_11, COMP_LOOP_11_modExp_dev_1_while_C_12,
      COMP_LOOP_11_modExp_dev_1_while_C_13, COMP_LOOP_11_modExp_dev_1_while_C_14,
      COMP_LOOP_C_322, COMP_LOOP_C_323, COMP_LOOP_C_324, COMP_LOOP_C_325, COMP_LOOP_C_326,
      COMP_LOOP_C_327, COMP_LOOP_C_328, COMP_LOOP_C_329, COMP_LOOP_C_330, COMP_LOOP_C_331,
      COMP_LOOP_C_332, COMP_LOOP_C_333, COMP_LOOP_C_334, COMP_LOOP_C_335, COMP_LOOP_C_336,
      COMP_LOOP_C_337, COMP_LOOP_C_338, COMP_LOOP_C_339, COMP_LOOP_C_340, COMP_LOOP_C_341,
      COMP_LOOP_C_342, COMP_LOOP_C_343, COMP_LOOP_C_344, COMP_LOOP_C_345, COMP_LOOP_C_346,
      COMP_LOOP_C_347, COMP_LOOP_C_348, COMP_LOOP_C_349, COMP_LOOP_C_350, COMP_LOOP_C_351,
      COMP_LOOP_C_352, COMP_LOOP_C_353, COMP_LOOP_12_modExp_dev_1_while_C_0, COMP_LOOP_12_modExp_dev_1_while_C_1,
      COMP_LOOP_12_modExp_dev_1_while_C_2, COMP_LOOP_12_modExp_dev_1_while_C_3, COMP_LOOP_12_modExp_dev_1_while_C_4,
      COMP_LOOP_12_modExp_dev_1_while_C_5, COMP_LOOP_12_modExp_dev_1_while_C_6, COMP_LOOP_12_modExp_dev_1_while_C_7,
      COMP_LOOP_12_modExp_dev_1_while_C_8, COMP_LOOP_12_modExp_dev_1_while_C_9, COMP_LOOP_12_modExp_dev_1_while_C_10,
      COMP_LOOP_12_modExp_dev_1_while_C_11, COMP_LOOP_12_modExp_dev_1_while_C_12,
      COMP_LOOP_12_modExp_dev_1_while_C_13, COMP_LOOP_12_modExp_dev_1_while_C_14,
      COMP_LOOP_C_354, COMP_LOOP_C_355, COMP_LOOP_C_356, COMP_LOOP_C_357, COMP_LOOP_C_358,
      COMP_LOOP_C_359, COMP_LOOP_C_360, COMP_LOOP_C_361, COMP_LOOP_C_362, COMP_LOOP_C_363,
      COMP_LOOP_C_364, COMP_LOOP_C_365, COMP_LOOP_C_366, COMP_LOOP_C_367, COMP_LOOP_C_368,
      COMP_LOOP_C_369, COMP_LOOP_C_370, COMP_LOOP_C_371, COMP_LOOP_C_372, COMP_LOOP_C_373,
      COMP_LOOP_C_374, COMP_LOOP_C_375, COMP_LOOP_C_376, COMP_LOOP_C_377, COMP_LOOP_C_378,
      COMP_LOOP_C_379, COMP_LOOP_C_380, COMP_LOOP_C_381, COMP_LOOP_C_382, COMP_LOOP_C_383,
      COMP_LOOP_C_384, COMP_LOOP_C_385, COMP_LOOP_13_modExp_dev_1_while_C_0, COMP_LOOP_13_modExp_dev_1_while_C_1,
      COMP_LOOP_13_modExp_dev_1_while_C_2, COMP_LOOP_13_modExp_dev_1_while_C_3, COMP_LOOP_13_modExp_dev_1_while_C_4,
      COMP_LOOP_13_modExp_dev_1_while_C_5, COMP_LOOP_13_modExp_dev_1_while_C_6, COMP_LOOP_13_modExp_dev_1_while_C_7,
      COMP_LOOP_13_modExp_dev_1_while_C_8, COMP_LOOP_13_modExp_dev_1_while_C_9, COMP_LOOP_13_modExp_dev_1_while_C_10,
      COMP_LOOP_13_modExp_dev_1_while_C_11, COMP_LOOP_13_modExp_dev_1_while_C_12,
      COMP_LOOP_13_modExp_dev_1_while_C_13, COMP_LOOP_13_modExp_dev_1_while_C_14,
      COMP_LOOP_C_386, COMP_LOOP_C_387, COMP_LOOP_C_388, COMP_LOOP_C_389, COMP_LOOP_C_390,
      COMP_LOOP_C_391, COMP_LOOP_C_392, COMP_LOOP_C_393, COMP_LOOP_C_394, COMP_LOOP_C_395,
      COMP_LOOP_C_396, COMP_LOOP_C_397, COMP_LOOP_C_398, COMP_LOOP_C_399, COMP_LOOP_C_400,
      COMP_LOOP_C_401, COMP_LOOP_C_402, COMP_LOOP_C_403, COMP_LOOP_C_404, COMP_LOOP_C_405,
      COMP_LOOP_C_406, COMP_LOOP_C_407, COMP_LOOP_C_408, COMP_LOOP_C_409, COMP_LOOP_C_410,
      COMP_LOOP_C_411, COMP_LOOP_C_412, COMP_LOOP_C_413, COMP_LOOP_C_414, COMP_LOOP_C_415,
      COMP_LOOP_C_416, COMP_LOOP_C_417, COMP_LOOP_14_modExp_dev_1_while_C_0, COMP_LOOP_14_modExp_dev_1_while_C_1,
      COMP_LOOP_14_modExp_dev_1_while_C_2, COMP_LOOP_14_modExp_dev_1_while_C_3, COMP_LOOP_14_modExp_dev_1_while_C_4,
      COMP_LOOP_14_modExp_dev_1_while_C_5, COMP_LOOP_14_modExp_dev_1_while_C_6, COMP_LOOP_14_modExp_dev_1_while_C_7,
      COMP_LOOP_14_modExp_dev_1_while_C_8, COMP_LOOP_14_modExp_dev_1_while_C_9, COMP_LOOP_14_modExp_dev_1_while_C_10,
      COMP_LOOP_14_modExp_dev_1_while_C_11, COMP_LOOP_14_modExp_dev_1_while_C_12,
      COMP_LOOP_14_modExp_dev_1_while_C_13, COMP_LOOP_14_modExp_dev_1_while_C_14,
      COMP_LOOP_C_418, COMP_LOOP_C_419, COMP_LOOP_C_420, COMP_LOOP_C_421, COMP_LOOP_C_422,
      COMP_LOOP_C_423, COMP_LOOP_C_424, COMP_LOOP_C_425, COMP_LOOP_C_426, COMP_LOOP_C_427,
      COMP_LOOP_C_428, COMP_LOOP_C_429, COMP_LOOP_C_430, COMP_LOOP_C_431, COMP_LOOP_C_432,
      COMP_LOOP_C_433, COMP_LOOP_C_434, COMP_LOOP_C_435, COMP_LOOP_C_436, COMP_LOOP_C_437,
      COMP_LOOP_C_438, COMP_LOOP_C_439, COMP_LOOP_C_440, COMP_LOOP_C_441, COMP_LOOP_C_442,
      COMP_LOOP_C_443, COMP_LOOP_C_444, COMP_LOOP_C_445, COMP_LOOP_C_446, COMP_LOOP_C_447,
      COMP_LOOP_C_448, COMP_LOOP_C_449, COMP_LOOP_15_modExp_dev_1_while_C_0, COMP_LOOP_15_modExp_dev_1_while_C_1,
      COMP_LOOP_15_modExp_dev_1_while_C_2, COMP_LOOP_15_modExp_dev_1_while_C_3, COMP_LOOP_15_modExp_dev_1_while_C_4,
      COMP_LOOP_15_modExp_dev_1_while_C_5, COMP_LOOP_15_modExp_dev_1_while_C_6, COMP_LOOP_15_modExp_dev_1_while_C_7,
      COMP_LOOP_15_modExp_dev_1_while_C_8, COMP_LOOP_15_modExp_dev_1_while_C_9, COMP_LOOP_15_modExp_dev_1_while_C_10,
      COMP_LOOP_15_modExp_dev_1_while_C_11, COMP_LOOP_15_modExp_dev_1_while_C_12,
      COMP_LOOP_15_modExp_dev_1_while_C_13, COMP_LOOP_15_modExp_dev_1_while_C_14,
      COMP_LOOP_C_450, COMP_LOOP_C_451, COMP_LOOP_C_452, COMP_LOOP_C_453, COMP_LOOP_C_454,
      COMP_LOOP_C_455, COMP_LOOP_C_456, COMP_LOOP_C_457, COMP_LOOP_C_458, COMP_LOOP_C_459,
      COMP_LOOP_C_460, COMP_LOOP_C_461, COMP_LOOP_C_462, COMP_LOOP_C_463, COMP_LOOP_C_464,
      COMP_LOOP_C_465, COMP_LOOP_C_466, COMP_LOOP_C_467, COMP_LOOP_C_468, COMP_LOOP_C_469,
      COMP_LOOP_C_470, COMP_LOOP_C_471, COMP_LOOP_C_472, COMP_LOOP_C_473, COMP_LOOP_C_474,
      COMP_LOOP_C_475, COMP_LOOP_C_476, COMP_LOOP_C_477, COMP_LOOP_C_478, COMP_LOOP_C_479,
      COMP_LOOP_C_480, COMP_LOOP_C_481, COMP_LOOP_16_modExp_dev_1_while_C_0, COMP_LOOP_16_modExp_dev_1_while_C_1,
      COMP_LOOP_16_modExp_dev_1_while_C_2, COMP_LOOP_16_modExp_dev_1_while_C_3, COMP_LOOP_16_modExp_dev_1_while_C_4,
      COMP_LOOP_16_modExp_dev_1_while_C_5, COMP_LOOP_16_modExp_dev_1_while_C_6, COMP_LOOP_16_modExp_dev_1_while_C_7,
      COMP_LOOP_16_modExp_dev_1_while_C_8, COMP_LOOP_16_modExp_dev_1_while_C_9, COMP_LOOP_16_modExp_dev_1_while_C_10,
      COMP_LOOP_16_modExp_dev_1_while_C_11, COMP_LOOP_16_modExp_dev_1_while_C_12,
      COMP_LOOP_16_modExp_dev_1_while_C_13, COMP_LOOP_16_modExp_dev_1_while_C_14,
      COMP_LOOP_C_482, COMP_LOOP_C_483, COMP_LOOP_C_484, COMP_LOOP_C_485, COMP_LOOP_C_486,
      COMP_LOOP_C_487, COMP_LOOP_C_488, COMP_LOOP_C_489, COMP_LOOP_C_490, COMP_LOOP_C_491,
      COMP_LOOP_C_492, COMP_LOOP_C_493, COMP_LOOP_C_494, COMP_LOOP_C_495, COMP_LOOP_C_496,
      COMP_LOOP_C_497, COMP_LOOP_C_498, COMP_LOOP_C_499, COMP_LOOP_C_500, COMP_LOOP_C_501,
      COMP_LOOP_C_502, COMP_LOOP_C_503, COMP_LOOP_C_504, COMP_LOOP_C_505, COMP_LOOP_C_506,
      COMP_LOOP_C_507, COMP_LOOP_C_508, COMP_LOOP_C_509, COMP_LOOP_C_510, COMP_LOOP_C_511,
      COMP_LOOP_C_512, VEC_LOOP_C_0, STAGE_LOOP_C_4, main_C_1);

  SIGNAL state_var : inPlaceNTT_DIT_core_core_fsm_1_ST;
  SIGNAL state_var_NS : inPlaceNTT_DIT_core_core_fsm_1_ST;

BEGIN
  inPlaceNTT_DIT_core_core_fsm_1 : PROCESS (STAGE_LOOP_C_3_tr0, modExp_dev_while_C_14_tr0,
      COMP_LOOP_C_1_tr0, COMP_LOOP_1_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_32_tr0,
      COMP_LOOP_2_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_64_tr0, COMP_LOOP_3_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_96_tr0, COMP_LOOP_4_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_128_tr0,
      COMP_LOOP_5_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_160_tr0, COMP_LOOP_6_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_192_tr0, COMP_LOOP_7_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_224_tr0,
      COMP_LOOP_8_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_256_tr0, COMP_LOOP_9_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_288_tr0, COMP_LOOP_10_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_320_tr0,
      COMP_LOOP_11_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_352_tr0, COMP_LOOP_12_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_384_tr0, COMP_LOOP_13_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_416_tr0,
      COMP_LOOP_14_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_448_tr0, COMP_LOOP_15_modExp_dev_1_while_C_14_tr0,
      COMP_LOOP_C_480_tr0, COMP_LOOP_16_modExp_dev_1_while_C_14_tr0, COMP_LOOP_C_512_tr0,
      VEC_LOOP_C_0_tr0, STAGE_LOOP_C_4_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000001");
        state_var_NS <= STAGE_LOOP_C_1;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000010");
        state_var_NS <= STAGE_LOOP_C_2;
      WHEN STAGE_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000011");
        state_var_NS <= STAGE_LOOP_C_3;
      WHEN STAGE_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000100");
        IF ( STAGE_LOOP_C_3_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_dev_while_C_0;
        END IF;
      WHEN modExp_dev_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000101");
        state_var_NS <= modExp_dev_while_C_1;
      WHEN modExp_dev_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000110");
        state_var_NS <= modExp_dev_while_C_2;
      WHEN modExp_dev_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000111");
        state_var_NS <= modExp_dev_while_C_3;
      WHEN modExp_dev_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001000");
        state_var_NS <= modExp_dev_while_C_4;
      WHEN modExp_dev_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001001");
        state_var_NS <= modExp_dev_while_C_5;
      WHEN modExp_dev_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001010");
        state_var_NS <= modExp_dev_while_C_6;
      WHEN modExp_dev_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001011");
        state_var_NS <= modExp_dev_while_C_7;
      WHEN modExp_dev_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001100");
        state_var_NS <= modExp_dev_while_C_8;
      WHEN modExp_dev_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001101");
        state_var_NS <= modExp_dev_while_C_9;
      WHEN modExp_dev_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001110");
        state_var_NS <= modExp_dev_while_C_10;
      WHEN modExp_dev_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001111");
        state_var_NS <= modExp_dev_while_C_11;
      WHEN modExp_dev_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010000");
        state_var_NS <= modExp_dev_while_C_12;
      WHEN modExp_dev_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010001");
        state_var_NS <= modExp_dev_while_C_13;
      WHEN modExp_dev_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010010");
        state_var_NS <= modExp_dev_while_C_14;
      WHEN modExp_dev_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010011");
        IF ( modExp_dev_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_0;
        ELSE
          state_var_NS <= modExp_dev_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010100");
        state_var_NS <= COMP_LOOP_C_1;
      WHEN COMP_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010101");
        IF ( COMP_LOOP_C_1_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_2;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010110");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010111");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011000");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011001");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011010");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011011");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011100");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011101");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011110");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000011111");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100000");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100001");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100010");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100011");
        state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_1_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100100");
        IF ( COMP_LOOP_1_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_2;
        ELSE
          state_var_NS <= COMP_LOOP_1_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100101");
        state_var_NS <= COMP_LOOP_C_3;
      WHEN COMP_LOOP_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100110");
        state_var_NS <= COMP_LOOP_C_4;
      WHEN COMP_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100111");
        state_var_NS <= COMP_LOOP_C_5;
      WHEN COMP_LOOP_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101000");
        state_var_NS <= COMP_LOOP_C_6;
      WHEN COMP_LOOP_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101001");
        state_var_NS <= COMP_LOOP_C_7;
      WHEN COMP_LOOP_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101010");
        state_var_NS <= COMP_LOOP_C_8;
      WHEN COMP_LOOP_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101011");
        state_var_NS <= COMP_LOOP_C_9;
      WHEN COMP_LOOP_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101100");
        state_var_NS <= COMP_LOOP_C_10;
      WHEN COMP_LOOP_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101101");
        state_var_NS <= COMP_LOOP_C_11;
      WHEN COMP_LOOP_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101110");
        state_var_NS <= COMP_LOOP_C_12;
      WHEN COMP_LOOP_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000101111");
        state_var_NS <= COMP_LOOP_C_13;
      WHEN COMP_LOOP_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110000");
        state_var_NS <= COMP_LOOP_C_14;
      WHEN COMP_LOOP_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110001");
        state_var_NS <= COMP_LOOP_C_15;
      WHEN COMP_LOOP_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110010");
        state_var_NS <= COMP_LOOP_C_16;
      WHEN COMP_LOOP_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110011");
        state_var_NS <= COMP_LOOP_C_17;
      WHEN COMP_LOOP_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110100");
        state_var_NS <= COMP_LOOP_C_18;
      WHEN COMP_LOOP_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110101");
        state_var_NS <= COMP_LOOP_C_19;
      WHEN COMP_LOOP_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110110");
        state_var_NS <= COMP_LOOP_C_20;
      WHEN COMP_LOOP_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000110111");
        state_var_NS <= COMP_LOOP_C_21;
      WHEN COMP_LOOP_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111000");
        state_var_NS <= COMP_LOOP_C_22;
      WHEN COMP_LOOP_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111001");
        state_var_NS <= COMP_LOOP_C_23;
      WHEN COMP_LOOP_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111010");
        state_var_NS <= COMP_LOOP_C_24;
      WHEN COMP_LOOP_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111011");
        state_var_NS <= COMP_LOOP_C_25;
      WHEN COMP_LOOP_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111100");
        state_var_NS <= COMP_LOOP_C_26;
      WHEN COMP_LOOP_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111101");
        state_var_NS <= COMP_LOOP_C_27;
      WHEN COMP_LOOP_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111110");
        state_var_NS <= COMP_LOOP_C_28;
      WHEN COMP_LOOP_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000111111");
        state_var_NS <= COMP_LOOP_C_29;
      WHEN COMP_LOOP_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000000");
        state_var_NS <= COMP_LOOP_C_30;
      WHEN COMP_LOOP_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000001");
        state_var_NS <= COMP_LOOP_C_31;
      WHEN COMP_LOOP_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000010");
        state_var_NS <= COMP_LOOP_C_32;
      WHEN COMP_LOOP_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000011");
        IF ( COMP_LOOP_C_32_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_33;
        END IF;
      WHEN COMP_LOOP_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000100");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000101");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000110");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000111");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001000");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001001");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001010");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001011");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001100");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001101");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001110");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001001111");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010000");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010001");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010010");
        state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_2_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010011");
        IF ( COMP_LOOP_2_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_34;
        ELSE
          state_var_NS <= COMP_LOOP_2_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_34 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010100");
        state_var_NS <= COMP_LOOP_C_35;
      WHEN COMP_LOOP_C_35 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010101");
        state_var_NS <= COMP_LOOP_C_36;
      WHEN COMP_LOOP_C_36 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010110");
        state_var_NS <= COMP_LOOP_C_37;
      WHEN COMP_LOOP_C_37 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001010111");
        state_var_NS <= COMP_LOOP_C_38;
      WHEN COMP_LOOP_C_38 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011000");
        state_var_NS <= COMP_LOOP_C_39;
      WHEN COMP_LOOP_C_39 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011001");
        state_var_NS <= COMP_LOOP_C_40;
      WHEN COMP_LOOP_C_40 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011010");
        state_var_NS <= COMP_LOOP_C_41;
      WHEN COMP_LOOP_C_41 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011011");
        state_var_NS <= COMP_LOOP_C_42;
      WHEN COMP_LOOP_C_42 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011100");
        state_var_NS <= COMP_LOOP_C_43;
      WHEN COMP_LOOP_C_43 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011101");
        state_var_NS <= COMP_LOOP_C_44;
      WHEN COMP_LOOP_C_44 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011110");
        state_var_NS <= COMP_LOOP_C_45;
      WHEN COMP_LOOP_C_45 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001011111");
        state_var_NS <= COMP_LOOP_C_46;
      WHEN COMP_LOOP_C_46 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100000");
        state_var_NS <= COMP_LOOP_C_47;
      WHEN COMP_LOOP_C_47 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100001");
        state_var_NS <= COMP_LOOP_C_48;
      WHEN COMP_LOOP_C_48 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100010");
        state_var_NS <= COMP_LOOP_C_49;
      WHEN COMP_LOOP_C_49 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100011");
        state_var_NS <= COMP_LOOP_C_50;
      WHEN COMP_LOOP_C_50 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100100");
        state_var_NS <= COMP_LOOP_C_51;
      WHEN COMP_LOOP_C_51 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100101");
        state_var_NS <= COMP_LOOP_C_52;
      WHEN COMP_LOOP_C_52 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100110");
        state_var_NS <= COMP_LOOP_C_53;
      WHEN COMP_LOOP_C_53 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001100111");
        state_var_NS <= COMP_LOOP_C_54;
      WHEN COMP_LOOP_C_54 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101000");
        state_var_NS <= COMP_LOOP_C_55;
      WHEN COMP_LOOP_C_55 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101001");
        state_var_NS <= COMP_LOOP_C_56;
      WHEN COMP_LOOP_C_56 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101010");
        state_var_NS <= COMP_LOOP_C_57;
      WHEN COMP_LOOP_C_57 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101011");
        state_var_NS <= COMP_LOOP_C_58;
      WHEN COMP_LOOP_C_58 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101100");
        state_var_NS <= COMP_LOOP_C_59;
      WHEN COMP_LOOP_C_59 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101101");
        state_var_NS <= COMP_LOOP_C_60;
      WHEN COMP_LOOP_C_60 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101110");
        state_var_NS <= COMP_LOOP_C_61;
      WHEN COMP_LOOP_C_61 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001101111");
        state_var_NS <= COMP_LOOP_C_62;
      WHEN COMP_LOOP_C_62 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110000");
        state_var_NS <= COMP_LOOP_C_63;
      WHEN COMP_LOOP_C_63 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110001");
        state_var_NS <= COMP_LOOP_C_64;
      WHEN COMP_LOOP_C_64 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110010");
        IF ( COMP_LOOP_C_64_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_65;
        END IF;
      WHEN COMP_LOOP_C_65 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110011");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110100");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110101");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110110");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001110111");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111000");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111001");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111010");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111011");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111100");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111101");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111110");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001111111");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000000");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000001");
        state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_3_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000010");
        IF ( COMP_LOOP_3_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_66;
        ELSE
          state_var_NS <= COMP_LOOP_3_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_66 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000011");
        state_var_NS <= COMP_LOOP_C_67;
      WHEN COMP_LOOP_C_67 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000100");
        state_var_NS <= COMP_LOOP_C_68;
      WHEN COMP_LOOP_C_68 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000101");
        state_var_NS <= COMP_LOOP_C_69;
      WHEN COMP_LOOP_C_69 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000110");
        state_var_NS <= COMP_LOOP_C_70;
      WHEN COMP_LOOP_C_70 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000111");
        state_var_NS <= COMP_LOOP_C_71;
      WHEN COMP_LOOP_C_71 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001000");
        state_var_NS <= COMP_LOOP_C_72;
      WHEN COMP_LOOP_C_72 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001001");
        state_var_NS <= COMP_LOOP_C_73;
      WHEN COMP_LOOP_C_73 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001010");
        state_var_NS <= COMP_LOOP_C_74;
      WHEN COMP_LOOP_C_74 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001011");
        state_var_NS <= COMP_LOOP_C_75;
      WHEN COMP_LOOP_C_75 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001100");
        state_var_NS <= COMP_LOOP_C_76;
      WHEN COMP_LOOP_C_76 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001101");
        state_var_NS <= COMP_LOOP_C_77;
      WHEN COMP_LOOP_C_77 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001110");
        state_var_NS <= COMP_LOOP_C_78;
      WHEN COMP_LOOP_C_78 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010001111");
        state_var_NS <= COMP_LOOP_C_79;
      WHEN COMP_LOOP_C_79 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010000");
        state_var_NS <= COMP_LOOP_C_80;
      WHEN COMP_LOOP_C_80 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010001");
        state_var_NS <= COMP_LOOP_C_81;
      WHEN COMP_LOOP_C_81 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010010");
        state_var_NS <= COMP_LOOP_C_82;
      WHEN COMP_LOOP_C_82 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010011");
        state_var_NS <= COMP_LOOP_C_83;
      WHEN COMP_LOOP_C_83 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010100");
        state_var_NS <= COMP_LOOP_C_84;
      WHEN COMP_LOOP_C_84 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010101");
        state_var_NS <= COMP_LOOP_C_85;
      WHEN COMP_LOOP_C_85 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010110");
        state_var_NS <= COMP_LOOP_C_86;
      WHEN COMP_LOOP_C_86 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010010111");
        state_var_NS <= COMP_LOOP_C_87;
      WHEN COMP_LOOP_C_87 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011000");
        state_var_NS <= COMP_LOOP_C_88;
      WHEN COMP_LOOP_C_88 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011001");
        state_var_NS <= COMP_LOOP_C_89;
      WHEN COMP_LOOP_C_89 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011010");
        state_var_NS <= COMP_LOOP_C_90;
      WHEN COMP_LOOP_C_90 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011011");
        state_var_NS <= COMP_LOOP_C_91;
      WHEN COMP_LOOP_C_91 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011100");
        state_var_NS <= COMP_LOOP_C_92;
      WHEN COMP_LOOP_C_92 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011101");
        state_var_NS <= COMP_LOOP_C_93;
      WHEN COMP_LOOP_C_93 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011110");
        state_var_NS <= COMP_LOOP_C_94;
      WHEN COMP_LOOP_C_94 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010011111");
        state_var_NS <= COMP_LOOP_C_95;
      WHEN COMP_LOOP_C_95 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100000");
        state_var_NS <= COMP_LOOP_C_96;
      WHEN COMP_LOOP_C_96 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100001");
        IF ( COMP_LOOP_C_96_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_97;
        END IF;
      WHEN COMP_LOOP_C_97 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100010");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100011");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100100");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100101");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100110");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010100111");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101000");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101001");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101010");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101011");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101100");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101101");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101110");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010101111");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110000");
        state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_4_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110001");
        IF ( COMP_LOOP_4_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_98;
        ELSE
          state_var_NS <= COMP_LOOP_4_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_98 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110010");
        state_var_NS <= COMP_LOOP_C_99;
      WHEN COMP_LOOP_C_99 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110011");
        state_var_NS <= COMP_LOOP_C_100;
      WHEN COMP_LOOP_C_100 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110100");
        state_var_NS <= COMP_LOOP_C_101;
      WHEN COMP_LOOP_C_101 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110101");
        state_var_NS <= COMP_LOOP_C_102;
      WHEN COMP_LOOP_C_102 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110110");
        state_var_NS <= COMP_LOOP_C_103;
      WHEN COMP_LOOP_C_103 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010110111");
        state_var_NS <= COMP_LOOP_C_104;
      WHEN COMP_LOOP_C_104 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111000");
        state_var_NS <= COMP_LOOP_C_105;
      WHEN COMP_LOOP_C_105 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111001");
        state_var_NS <= COMP_LOOP_C_106;
      WHEN COMP_LOOP_C_106 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111010");
        state_var_NS <= COMP_LOOP_C_107;
      WHEN COMP_LOOP_C_107 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111011");
        state_var_NS <= COMP_LOOP_C_108;
      WHEN COMP_LOOP_C_108 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111100");
        state_var_NS <= COMP_LOOP_C_109;
      WHEN COMP_LOOP_C_109 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111101");
        state_var_NS <= COMP_LOOP_C_110;
      WHEN COMP_LOOP_C_110 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111110");
        state_var_NS <= COMP_LOOP_C_111;
      WHEN COMP_LOOP_C_111 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010111111");
        state_var_NS <= COMP_LOOP_C_112;
      WHEN COMP_LOOP_C_112 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000000");
        state_var_NS <= COMP_LOOP_C_113;
      WHEN COMP_LOOP_C_113 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000001");
        state_var_NS <= COMP_LOOP_C_114;
      WHEN COMP_LOOP_C_114 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000010");
        state_var_NS <= COMP_LOOP_C_115;
      WHEN COMP_LOOP_C_115 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000011");
        state_var_NS <= COMP_LOOP_C_116;
      WHEN COMP_LOOP_C_116 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000100");
        state_var_NS <= COMP_LOOP_C_117;
      WHEN COMP_LOOP_C_117 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000101");
        state_var_NS <= COMP_LOOP_C_118;
      WHEN COMP_LOOP_C_118 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000110");
        state_var_NS <= COMP_LOOP_C_119;
      WHEN COMP_LOOP_C_119 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011000111");
        state_var_NS <= COMP_LOOP_C_120;
      WHEN COMP_LOOP_C_120 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001000");
        state_var_NS <= COMP_LOOP_C_121;
      WHEN COMP_LOOP_C_121 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001001");
        state_var_NS <= COMP_LOOP_C_122;
      WHEN COMP_LOOP_C_122 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001010");
        state_var_NS <= COMP_LOOP_C_123;
      WHEN COMP_LOOP_C_123 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001011");
        state_var_NS <= COMP_LOOP_C_124;
      WHEN COMP_LOOP_C_124 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001100");
        state_var_NS <= COMP_LOOP_C_125;
      WHEN COMP_LOOP_C_125 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001101");
        state_var_NS <= COMP_LOOP_C_126;
      WHEN COMP_LOOP_C_126 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001110");
        state_var_NS <= COMP_LOOP_C_127;
      WHEN COMP_LOOP_C_127 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011001111");
        state_var_NS <= COMP_LOOP_C_128;
      WHEN COMP_LOOP_C_128 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010000");
        IF ( COMP_LOOP_C_128_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_129;
        END IF;
      WHEN COMP_LOOP_C_129 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010001");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010010");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010011");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010100");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010101");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010110");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011010111");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011000");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011001");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011010");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011011");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011100");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011101");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011110");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011011111");
        state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_5_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100000");
        IF ( COMP_LOOP_5_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_130;
        ELSE
          state_var_NS <= COMP_LOOP_5_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_130 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100001");
        state_var_NS <= COMP_LOOP_C_131;
      WHEN COMP_LOOP_C_131 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100010");
        state_var_NS <= COMP_LOOP_C_132;
      WHEN COMP_LOOP_C_132 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100011");
        state_var_NS <= COMP_LOOP_C_133;
      WHEN COMP_LOOP_C_133 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100100");
        state_var_NS <= COMP_LOOP_C_134;
      WHEN COMP_LOOP_C_134 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100101");
        state_var_NS <= COMP_LOOP_C_135;
      WHEN COMP_LOOP_C_135 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100110");
        state_var_NS <= COMP_LOOP_C_136;
      WHEN COMP_LOOP_C_136 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011100111");
        state_var_NS <= COMP_LOOP_C_137;
      WHEN COMP_LOOP_C_137 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101000");
        state_var_NS <= COMP_LOOP_C_138;
      WHEN COMP_LOOP_C_138 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101001");
        state_var_NS <= COMP_LOOP_C_139;
      WHEN COMP_LOOP_C_139 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101010");
        state_var_NS <= COMP_LOOP_C_140;
      WHEN COMP_LOOP_C_140 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101011");
        state_var_NS <= COMP_LOOP_C_141;
      WHEN COMP_LOOP_C_141 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101100");
        state_var_NS <= COMP_LOOP_C_142;
      WHEN COMP_LOOP_C_142 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101101");
        state_var_NS <= COMP_LOOP_C_143;
      WHEN COMP_LOOP_C_143 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101110");
        state_var_NS <= COMP_LOOP_C_144;
      WHEN COMP_LOOP_C_144 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011101111");
        state_var_NS <= COMP_LOOP_C_145;
      WHEN COMP_LOOP_C_145 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110000");
        state_var_NS <= COMP_LOOP_C_146;
      WHEN COMP_LOOP_C_146 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110001");
        state_var_NS <= COMP_LOOP_C_147;
      WHEN COMP_LOOP_C_147 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110010");
        state_var_NS <= COMP_LOOP_C_148;
      WHEN COMP_LOOP_C_148 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110011");
        state_var_NS <= COMP_LOOP_C_149;
      WHEN COMP_LOOP_C_149 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110100");
        state_var_NS <= COMP_LOOP_C_150;
      WHEN COMP_LOOP_C_150 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110101");
        state_var_NS <= COMP_LOOP_C_151;
      WHEN COMP_LOOP_C_151 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110110");
        state_var_NS <= COMP_LOOP_C_152;
      WHEN COMP_LOOP_C_152 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011110111");
        state_var_NS <= COMP_LOOP_C_153;
      WHEN COMP_LOOP_C_153 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111000");
        state_var_NS <= COMP_LOOP_C_154;
      WHEN COMP_LOOP_C_154 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111001");
        state_var_NS <= COMP_LOOP_C_155;
      WHEN COMP_LOOP_C_155 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111010");
        state_var_NS <= COMP_LOOP_C_156;
      WHEN COMP_LOOP_C_156 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111011");
        state_var_NS <= COMP_LOOP_C_157;
      WHEN COMP_LOOP_C_157 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111100");
        state_var_NS <= COMP_LOOP_C_158;
      WHEN COMP_LOOP_C_158 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111101");
        state_var_NS <= COMP_LOOP_C_159;
      WHEN COMP_LOOP_C_159 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111110");
        state_var_NS <= COMP_LOOP_C_160;
      WHEN COMP_LOOP_C_160 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0011111111");
        IF ( COMP_LOOP_C_160_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_161;
        END IF;
      WHEN COMP_LOOP_C_161 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000000");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000001");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000010");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000011");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000100");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000101");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000110");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000111");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001000");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001001");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001010");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001011");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001100");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001101");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001110");
        state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_6_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100001111");
        IF ( COMP_LOOP_6_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_162;
        ELSE
          state_var_NS <= COMP_LOOP_6_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_162 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010000");
        state_var_NS <= COMP_LOOP_C_163;
      WHEN COMP_LOOP_C_163 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010001");
        state_var_NS <= COMP_LOOP_C_164;
      WHEN COMP_LOOP_C_164 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010010");
        state_var_NS <= COMP_LOOP_C_165;
      WHEN COMP_LOOP_C_165 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010011");
        state_var_NS <= COMP_LOOP_C_166;
      WHEN COMP_LOOP_C_166 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010100");
        state_var_NS <= COMP_LOOP_C_167;
      WHEN COMP_LOOP_C_167 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010101");
        state_var_NS <= COMP_LOOP_C_168;
      WHEN COMP_LOOP_C_168 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010110");
        state_var_NS <= COMP_LOOP_C_169;
      WHEN COMP_LOOP_C_169 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100010111");
        state_var_NS <= COMP_LOOP_C_170;
      WHEN COMP_LOOP_C_170 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011000");
        state_var_NS <= COMP_LOOP_C_171;
      WHEN COMP_LOOP_C_171 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011001");
        state_var_NS <= COMP_LOOP_C_172;
      WHEN COMP_LOOP_C_172 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011010");
        state_var_NS <= COMP_LOOP_C_173;
      WHEN COMP_LOOP_C_173 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011011");
        state_var_NS <= COMP_LOOP_C_174;
      WHEN COMP_LOOP_C_174 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011100");
        state_var_NS <= COMP_LOOP_C_175;
      WHEN COMP_LOOP_C_175 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011101");
        state_var_NS <= COMP_LOOP_C_176;
      WHEN COMP_LOOP_C_176 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011110");
        state_var_NS <= COMP_LOOP_C_177;
      WHEN COMP_LOOP_C_177 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100011111");
        state_var_NS <= COMP_LOOP_C_178;
      WHEN COMP_LOOP_C_178 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100000");
        state_var_NS <= COMP_LOOP_C_179;
      WHEN COMP_LOOP_C_179 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100001");
        state_var_NS <= COMP_LOOP_C_180;
      WHEN COMP_LOOP_C_180 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100010");
        state_var_NS <= COMP_LOOP_C_181;
      WHEN COMP_LOOP_C_181 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100011");
        state_var_NS <= COMP_LOOP_C_182;
      WHEN COMP_LOOP_C_182 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100100");
        state_var_NS <= COMP_LOOP_C_183;
      WHEN COMP_LOOP_C_183 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100101");
        state_var_NS <= COMP_LOOP_C_184;
      WHEN COMP_LOOP_C_184 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100110");
        state_var_NS <= COMP_LOOP_C_185;
      WHEN COMP_LOOP_C_185 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100100111");
        state_var_NS <= COMP_LOOP_C_186;
      WHEN COMP_LOOP_C_186 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101000");
        state_var_NS <= COMP_LOOP_C_187;
      WHEN COMP_LOOP_C_187 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101001");
        state_var_NS <= COMP_LOOP_C_188;
      WHEN COMP_LOOP_C_188 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101010");
        state_var_NS <= COMP_LOOP_C_189;
      WHEN COMP_LOOP_C_189 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101011");
        state_var_NS <= COMP_LOOP_C_190;
      WHEN COMP_LOOP_C_190 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101100");
        state_var_NS <= COMP_LOOP_C_191;
      WHEN COMP_LOOP_C_191 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101101");
        state_var_NS <= COMP_LOOP_C_192;
      WHEN COMP_LOOP_C_192 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101110");
        IF ( COMP_LOOP_C_192_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_193;
        END IF;
      WHEN COMP_LOOP_C_193 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100101111");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110000");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110001");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110010");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110011");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110100");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110101");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110110");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100110111");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111000");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111001");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111010");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111011");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111100");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111101");
        state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_7_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111110");
        IF ( COMP_LOOP_7_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_194;
        ELSE
          state_var_NS <= COMP_LOOP_7_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_194 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100111111");
        state_var_NS <= COMP_LOOP_C_195;
      WHEN COMP_LOOP_C_195 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000000");
        state_var_NS <= COMP_LOOP_C_196;
      WHEN COMP_LOOP_C_196 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000001");
        state_var_NS <= COMP_LOOP_C_197;
      WHEN COMP_LOOP_C_197 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000010");
        state_var_NS <= COMP_LOOP_C_198;
      WHEN COMP_LOOP_C_198 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000011");
        state_var_NS <= COMP_LOOP_C_199;
      WHEN COMP_LOOP_C_199 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000100");
        state_var_NS <= COMP_LOOP_C_200;
      WHEN COMP_LOOP_C_200 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000101");
        state_var_NS <= COMP_LOOP_C_201;
      WHEN COMP_LOOP_C_201 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000110");
        state_var_NS <= COMP_LOOP_C_202;
      WHEN COMP_LOOP_C_202 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101000111");
        state_var_NS <= COMP_LOOP_C_203;
      WHEN COMP_LOOP_C_203 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001000");
        state_var_NS <= COMP_LOOP_C_204;
      WHEN COMP_LOOP_C_204 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001001");
        state_var_NS <= COMP_LOOP_C_205;
      WHEN COMP_LOOP_C_205 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001010");
        state_var_NS <= COMP_LOOP_C_206;
      WHEN COMP_LOOP_C_206 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001011");
        state_var_NS <= COMP_LOOP_C_207;
      WHEN COMP_LOOP_C_207 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001100");
        state_var_NS <= COMP_LOOP_C_208;
      WHEN COMP_LOOP_C_208 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001101");
        state_var_NS <= COMP_LOOP_C_209;
      WHEN COMP_LOOP_C_209 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001110");
        state_var_NS <= COMP_LOOP_C_210;
      WHEN COMP_LOOP_C_210 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101001111");
        state_var_NS <= COMP_LOOP_C_211;
      WHEN COMP_LOOP_C_211 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010000");
        state_var_NS <= COMP_LOOP_C_212;
      WHEN COMP_LOOP_C_212 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010001");
        state_var_NS <= COMP_LOOP_C_213;
      WHEN COMP_LOOP_C_213 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010010");
        state_var_NS <= COMP_LOOP_C_214;
      WHEN COMP_LOOP_C_214 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010011");
        state_var_NS <= COMP_LOOP_C_215;
      WHEN COMP_LOOP_C_215 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010100");
        state_var_NS <= COMP_LOOP_C_216;
      WHEN COMP_LOOP_C_216 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010101");
        state_var_NS <= COMP_LOOP_C_217;
      WHEN COMP_LOOP_C_217 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010110");
        state_var_NS <= COMP_LOOP_C_218;
      WHEN COMP_LOOP_C_218 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101010111");
        state_var_NS <= COMP_LOOP_C_219;
      WHEN COMP_LOOP_C_219 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011000");
        state_var_NS <= COMP_LOOP_C_220;
      WHEN COMP_LOOP_C_220 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011001");
        state_var_NS <= COMP_LOOP_C_221;
      WHEN COMP_LOOP_C_221 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011010");
        state_var_NS <= COMP_LOOP_C_222;
      WHEN COMP_LOOP_C_222 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011011");
        state_var_NS <= COMP_LOOP_C_223;
      WHEN COMP_LOOP_C_223 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011100");
        state_var_NS <= COMP_LOOP_C_224;
      WHEN COMP_LOOP_C_224 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011101");
        IF ( COMP_LOOP_C_224_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_225;
        END IF;
      WHEN COMP_LOOP_C_225 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011110");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101011111");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100000");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100001");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100010");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100011");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100100");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100101");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100110");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101100111");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101000");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101001");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101010");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101011");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101100");
        state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_8_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101101");
        IF ( COMP_LOOP_8_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_226;
        ELSE
          state_var_NS <= COMP_LOOP_8_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_226 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101110");
        state_var_NS <= COMP_LOOP_C_227;
      WHEN COMP_LOOP_C_227 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101101111");
        state_var_NS <= COMP_LOOP_C_228;
      WHEN COMP_LOOP_C_228 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110000");
        state_var_NS <= COMP_LOOP_C_229;
      WHEN COMP_LOOP_C_229 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110001");
        state_var_NS <= COMP_LOOP_C_230;
      WHEN COMP_LOOP_C_230 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110010");
        state_var_NS <= COMP_LOOP_C_231;
      WHEN COMP_LOOP_C_231 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110011");
        state_var_NS <= COMP_LOOP_C_232;
      WHEN COMP_LOOP_C_232 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110100");
        state_var_NS <= COMP_LOOP_C_233;
      WHEN COMP_LOOP_C_233 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110101");
        state_var_NS <= COMP_LOOP_C_234;
      WHEN COMP_LOOP_C_234 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110110");
        state_var_NS <= COMP_LOOP_C_235;
      WHEN COMP_LOOP_C_235 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101110111");
        state_var_NS <= COMP_LOOP_C_236;
      WHEN COMP_LOOP_C_236 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111000");
        state_var_NS <= COMP_LOOP_C_237;
      WHEN COMP_LOOP_C_237 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111001");
        state_var_NS <= COMP_LOOP_C_238;
      WHEN COMP_LOOP_C_238 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111010");
        state_var_NS <= COMP_LOOP_C_239;
      WHEN COMP_LOOP_C_239 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111011");
        state_var_NS <= COMP_LOOP_C_240;
      WHEN COMP_LOOP_C_240 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111100");
        state_var_NS <= COMP_LOOP_C_241;
      WHEN COMP_LOOP_C_241 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111101");
        state_var_NS <= COMP_LOOP_C_242;
      WHEN COMP_LOOP_C_242 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111110");
        state_var_NS <= COMP_LOOP_C_243;
      WHEN COMP_LOOP_C_243 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0101111111");
        state_var_NS <= COMP_LOOP_C_244;
      WHEN COMP_LOOP_C_244 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000000");
        state_var_NS <= COMP_LOOP_C_245;
      WHEN COMP_LOOP_C_245 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000001");
        state_var_NS <= COMP_LOOP_C_246;
      WHEN COMP_LOOP_C_246 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000010");
        state_var_NS <= COMP_LOOP_C_247;
      WHEN COMP_LOOP_C_247 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000011");
        state_var_NS <= COMP_LOOP_C_248;
      WHEN COMP_LOOP_C_248 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000100");
        state_var_NS <= COMP_LOOP_C_249;
      WHEN COMP_LOOP_C_249 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000101");
        state_var_NS <= COMP_LOOP_C_250;
      WHEN COMP_LOOP_C_250 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000110");
        state_var_NS <= COMP_LOOP_C_251;
      WHEN COMP_LOOP_C_251 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110000111");
        state_var_NS <= COMP_LOOP_C_252;
      WHEN COMP_LOOP_C_252 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001000");
        state_var_NS <= COMP_LOOP_C_253;
      WHEN COMP_LOOP_C_253 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001001");
        state_var_NS <= COMP_LOOP_C_254;
      WHEN COMP_LOOP_C_254 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001010");
        state_var_NS <= COMP_LOOP_C_255;
      WHEN COMP_LOOP_C_255 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001011");
        state_var_NS <= COMP_LOOP_C_256;
      WHEN COMP_LOOP_C_256 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001100");
        IF ( COMP_LOOP_C_256_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_257;
        END IF;
      WHEN COMP_LOOP_C_257 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001101");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001110");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110001111");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010000");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010001");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010010");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010011");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010100");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010101");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010110");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110010111");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011000");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011001");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011010");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011011");
        state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_9_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011100");
        IF ( COMP_LOOP_9_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_258;
        ELSE
          state_var_NS <= COMP_LOOP_9_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_258 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011101");
        state_var_NS <= COMP_LOOP_C_259;
      WHEN COMP_LOOP_C_259 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011110");
        state_var_NS <= COMP_LOOP_C_260;
      WHEN COMP_LOOP_C_260 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110011111");
        state_var_NS <= COMP_LOOP_C_261;
      WHEN COMP_LOOP_C_261 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100000");
        state_var_NS <= COMP_LOOP_C_262;
      WHEN COMP_LOOP_C_262 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100001");
        state_var_NS <= COMP_LOOP_C_263;
      WHEN COMP_LOOP_C_263 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100010");
        state_var_NS <= COMP_LOOP_C_264;
      WHEN COMP_LOOP_C_264 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100011");
        state_var_NS <= COMP_LOOP_C_265;
      WHEN COMP_LOOP_C_265 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100100");
        state_var_NS <= COMP_LOOP_C_266;
      WHEN COMP_LOOP_C_266 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100101");
        state_var_NS <= COMP_LOOP_C_267;
      WHEN COMP_LOOP_C_267 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100110");
        state_var_NS <= COMP_LOOP_C_268;
      WHEN COMP_LOOP_C_268 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110100111");
        state_var_NS <= COMP_LOOP_C_269;
      WHEN COMP_LOOP_C_269 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101000");
        state_var_NS <= COMP_LOOP_C_270;
      WHEN COMP_LOOP_C_270 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101001");
        state_var_NS <= COMP_LOOP_C_271;
      WHEN COMP_LOOP_C_271 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101010");
        state_var_NS <= COMP_LOOP_C_272;
      WHEN COMP_LOOP_C_272 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101011");
        state_var_NS <= COMP_LOOP_C_273;
      WHEN COMP_LOOP_C_273 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101100");
        state_var_NS <= COMP_LOOP_C_274;
      WHEN COMP_LOOP_C_274 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101101");
        state_var_NS <= COMP_LOOP_C_275;
      WHEN COMP_LOOP_C_275 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101110");
        state_var_NS <= COMP_LOOP_C_276;
      WHEN COMP_LOOP_C_276 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110101111");
        state_var_NS <= COMP_LOOP_C_277;
      WHEN COMP_LOOP_C_277 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110000");
        state_var_NS <= COMP_LOOP_C_278;
      WHEN COMP_LOOP_C_278 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110001");
        state_var_NS <= COMP_LOOP_C_279;
      WHEN COMP_LOOP_C_279 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110010");
        state_var_NS <= COMP_LOOP_C_280;
      WHEN COMP_LOOP_C_280 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110011");
        state_var_NS <= COMP_LOOP_C_281;
      WHEN COMP_LOOP_C_281 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110100");
        state_var_NS <= COMP_LOOP_C_282;
      WHEN COMP_LOOP_C_282 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110101");
        state_var_NS <= COMP_LOOP_C_283;
      WHEN COMP_LOOP_C_283 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110110");
        state_var_NS <= COMP_LOOP_C_284;
      WHEN COMP_LOOP_C_284 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110110111");
        state_var_NS <= COMP_LOOP_C_285;
      WHEN COMP_LOOP_C_285 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111000");
        state_var_NS <= COMP_LOOP_C_286;
      WHEN COMP_LOOP_C_286 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111001");
        state_var_NS <= COMP_LOOP_C_287;
      WHEN COMP_LOOP_C_287 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111010");
        state_var_NS <= COMP_LOOP_C_288;
      WHEN COMP_LOOP_C_288 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111011");
        IF ( COMP_LOOP_C_288_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_289;
        END IF;
      WHEN COMP_LOOP_C_289 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111100");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111101");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111110");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0110111111");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000000");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000001");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000010");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000011");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000100");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000101");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000110");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111000111");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001000");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001001");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001010");
        state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_10_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001011");
        IF ( COMP_LOOP_10_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_290;
        ELSE
          state_var_NS <= COMP_LOOP_10_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_290 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001100");
        state_var_NS <= COMP_LOOP_C_291;
      WHEN COMP_LOOP_C_291 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001101");
        state_var_NS <= COMP_LOOP_C_292;
      WHEN COMP_LOOP_C_292 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001110");
        state_var_NS <= COMP_LOOP_C_293;
      WHEN COMP_LOOP_C_293 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111001111");
        state_var_NS <= COMP_LOOP_C_294;
      WHEN COMP_LOOP_C_294 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010000");
        state_var_NS <= COMP_LOOP_C_295;
      WHEN COMP_LOOP_C_295 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010001");
        state_var_NS <= COMP_LOOP_C_296;
      WHEN COMP_LOOP_C_296 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010010");
        state_var_NS <= COMP_LOOP_C_297;
      WHEN COMP_LOOP_C_297 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010011");
        state_var_NS <= COMP_LOOP_C_298;
      WHEN COMP_LOOP_C_298 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010100");
        state_var_NS <= COMP_LOOP_C_299;
      WHEN COMP_LOOP_C_299 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010101");
        state_var_NS <= COMP_LOOP_C_300;
      WHEN COMP_LOOP_C_300 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010110");
        state_var_NS <= COMP_LOOP_C_301;
      WHEN COMP_LOOP_C_301 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111010111");
        state_var_NS <= COMP_LOOP_C_302;
      WHEN COMP_LOOP_C_302 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011000");
        state_var_NS <= COMP_LOOP_C_303;
      WHEN COMP_LOOP_C_303 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011001");
        state_var_NS <= COMP_LOOP_C_304;
      WHEN COMP_LOOP_C_304 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011010");
        state_var_NS <= COMP_LOOP_C_305;
      WHEN COMP_LOOP_C_305 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011011");
        state_var_NS <= COMP_LOOP_C_306;
      WHEN COMP_LOOP_C_306 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011100");
        state_var_NS <= COMP_LOOP_C_307;
      WHEN COMP_LOOP_C_307 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011101");
        state_var_NS <= COMP_LOOP_C_308;
      WHEN COMP_LOOP_C_308 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011110");
        state_var_NS <= COMP_LOOP_C_309;
      WHEN COMP_LOOP_C_309 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111011111");
        state_var_NS <= COMP_LOOP_C_310;
      WHEN COMP_LOOP_C_310 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100000");
        state_var_NS <= COMP_LOOP_C_311;
      WHEN COMP_LOOP_C_311 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100001");
        state_var_NS <= COMP_LOOP_C_312;
      WHEN COMP_LOOP_C_312 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100010");
        state_var_NS <= COMP_LOOP_C_313;
      WHEN COMP_LOOP_C_313 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100011");
        state_var_NS <= COMP_LOOP_C_314;
      WHEN COMP_LOOP_C_314 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100100");
        state_var_NS <= COMP_LOOP_C_315;
      WHEN COMP_LOOP_C_315 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100101");
        state_var_NS <= COMP_LOOP_C_316;
      WHEN COMP_LOOP_C_316 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100110");
        state_var_NS <= COMP_LOOP_C_317;
      WHEN COMP_LOOP_C_317 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111100111");
        state_var_NS <= COMP_LOOP_C_318;
      WHEN COMP_LOOP_C_318 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101000");
        state_var_NS <= COMP_LOOP_C_319;
      WHEN COMP_LOOP_C_319 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101001");
        state_var_NS <= COMP_LOOP_C_320;
      WHEN COMP_LOOP_C_320 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101010");
        IF ( COMP_LOOP_C_320_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_321;
        END IF;
      WHEN COMP_LOOP_C_321 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101011");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101100");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101101");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101110");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111101111");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110000");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110001");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110010");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110011");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110100");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110101");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110110");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111110111");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111000");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111001");
        state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_11_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111010");
        IF ( COMP_LOOP_11_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_322;
        ELSE
          state_var_NS <= COMP_LOOP_11_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_322 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111011");
        state_var_NS <= COMP_LOOP_C_323;
      WHEN COMP_LOOP_C_323 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111100");
        state_var_NS <= COMP_LOOP_C_324;
      WHEN COMP_LOOP_C_324 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111101");
        state_var_NS <= COMP_LOOP_C_325;
      WHEN COMP_LOOP_C_325 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111110");
        state_var_NS <= COMP_LOOP_C_326;
      WHEN COMP_LOOP_C_326 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0111111111");
        state_var_NS <= COMP_LOOP_C_327;
      WHEN COMP_LOOP_C_327 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000000");
        state_var_NS <= COMP_LOOP_C_328;
      WHEN COMP_LOOP_C_328 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000001");
        state_var_NS <= COMP_LOOP_C_329;
      WHEN COMP_LOOP_C_329 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000010");
        state_var_NS <= COMP_LOOP_C_330;
      WHEN COMP_LOOP_C_330 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000011");
        state_var_NS <= COMP_LOOP_C_331;
      WHEN COMP_LOOP_C_331 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000100");
        state_var_NS <= COMP_LOOP_C_332;
      WHEN COMP_LOOP_C_332 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000101");
        state_var_NS <= COMP_LOOP_C_333;
      WHEN COMP_LOOP_C_333 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000110");
        state_var_NS <= COMP_LOOP_C_334;
      WHEN COMP_LOOP_C_334 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000111");
        state_var_NS <= COMP_LOOP_C_335;
      WHEN COMP_LOOP_C_335 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001000");
        state_var_NS <= COMP_LOOP_C_336;
      WHEN COMP_LOOP_C_336 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001001");
        state_var_NS <= COMP_LOOP_C_337;
      WHEN COMP_LOOP_C_337 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001010");
        state_var_NS <= COMP_LOOP_C_338;
      WHEN COMP_LOOP_C_338 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001011");
        state_var_NS <= COMP_LOOP_C_339;
      WHEN COMP_LOOP_C_339 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001100");
        state_var_NS <= COMP_LOOP_C_340;
      WHEN COMP_LOOP_C_340 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001101");
        state_var_NS <= COMP_LOOP_C_341;
      WHEN COMP_LOOP_C_341 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001110");
        state_var_NS <= COMP_LOOP_C_342;
      WHEN COMP_LOOP_C_342 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000001111");
        state_var_NS <= COMP_LOOP_C_343;
      WHEN COMP_LOOP_C_343 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010000");
        state_var_NS <= COMP_LOOP_C_344;
      WHEN COMP_LOOP_C_344 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010001");
        state_var_NS <= COMP_LOOP_C_345;
      WHEN COMP_LOOP_C_345 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010010");
        state_var_NS <= COMP_LOOP_C_346;
      WHEN COMP_LOOP_C_346 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010011");
        state_var_NS <= COMP_LOOP_C_347;
      WHEN COMP_LOOP_C_347 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010100");
        state_var_NS <= COMP_LOOP_C_348;
      WHEN COMP_LOOP_C_348 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010101");
        state_var_NS <= COMP_LOOP_C_349;
      WHEN COMP_LOOP_C_349 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010110");
        state_var_NS <= COMP_LOOP_C_350;
      WHEN COMP_LOOP_C_350 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000010111");
        state_var_NS <= COMP_LOOP_C_351;
      WHEN COMP_LOOP_C_351 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011000");
        state_var_NS <= COMP_LOOP_C_352;
      WHEN COMP_LOOP_C_352 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011001");
        IF ( COMP_LOOP_C_352_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_353;
        END IF;
      WHEN COMP_LOOP_C_353 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011010");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011011");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011100");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011101");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011110");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000011111");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100000");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100001");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100010");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100011");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100100");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100101");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100110");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000100111");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101000");
        state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_12_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101001");
        IF ( COMP_LOOP_12_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_354;
        ELSE
          state_var_NS <= COMP_LOOP_12_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_354 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101010");
        state_var_NS <= COMP_LOOP_C_355;
      WHEN COMP_LOOP_C_355 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101011");
        state_var_NS <= COMP_LOOP_C_356;
      WHEN COMP_LOOP_C_356 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101100");
        state_var_NS <= COMP_LOOP_C_357;
      WHEN COMP_LOOP_C_357 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101101");
        state_var_NS <= COMP_LOOP_C_358;
      WHEN COMP_LOOP_C_358 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101110");
        state_var_NS <= COMP_LOOP_C_359;
      WHEN COMP_LOOP_C_359 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000101111");
        state_var_NS <= COMP_LOOP_C_360;
      WHEN COMP_LOOP_C_360 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110000");
        state_var_NS <= COMP_LOOP_C_361;
      WHEN COMP_LOOP_C_361 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110001");
        state_var_NS <= COMP_LOOP_C_362;
      WHEN COMP_LOOP_C_362 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110010");
        state_var_NS <= COMP_LOOP_C_363;
      WHEN COMP_LOOP_C_363 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110011");
        state_var_NS <= COMP_LOOP_C_364;
      WHEN COMP_LOOP_C_364 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110100");
        state_var_NS <= COMP_LOOP_C_365;
      WHEN COMP_LOOP_C_365 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110101");
        state_var_NS <= COMP_LOOP_C_366;
      WHEN COMP_LOOP_C_366 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110110");
        state_var_NS <= COMP_LOOP_C_367;
      WHEN COMP_LOOP_C_367 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000110111");
        state_var_NS <= COMP_LOOP_C_368;
      WHEN COMP_LOOP_C_368 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111000");
        state_var_NS <= COMP_LOOP_C_369;
      WHEN COMP_LOOP_C_369 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111001");
        state_var_NS <= COMP_LOOP_C_370;
      WHEN COMP_LOOP_C_370 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111010");
        state_var_NS <= COMP_LOOP_C_371;
      WHEN COMP_LOOP_C_371 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111011");
        state_var_NS <= COMP_LOOP_C_372;
      WHEN COMP_LOOP_C_372 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111100");
        state_var_NS <= COMP_LOOP_C_373;
      WHEN COMP_LOOP_C_373 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111101");
        state_var_NS <= COMP_LOOP_C_374;
      WHEN COMP_LOOP_C_374 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111110");
        state_var_NS <= COMP_LOOP_C_375;
      WHEN COMP_LOOP_C_375 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000111111");
        state_var_NS <= COMP_LOOP_C_376;
      WHEN COMP_LOOP_C_376 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000000");
        state_var_NS <= COMP_LOOP_C_377;
      WHEN COMP_LOOP_C_377 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000001");
        state_var_NS <= COMP_LOOP_C_378;
      WHEN COMP_LOOP_C_378 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000010");
        state_var_NS <= COMP_LOOP_C_379;
      WHEN COMP_LOOP_C_379 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000011");
        state_var_NS <= COMP_LOOP_C_380;
      WHEN COMP_LOOP_C_380 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000100");
        state_var_NS <= COMP_LOOP_C_381;
      WHEN COMP_LOOP_C_381 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000101");
        state_var_NS <= COMP_LOOP_C_382;
      WHEN COMP_LOOP_C_382 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000110");
        state_var_NS <= COMP_LOOP_C_383;
      WHEN COMP_LOOP_C_383 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001000111");
        state_var_NS <= COMP_LOOP_C_384;
      WHEN COMP_LOOP_C_384 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001000");
        IF ( COMP_LOOP_C_384_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_385;
        END IF;
      WHEN COMP_LOOP_C_385 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001001");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001010");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001011");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001100");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001101");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001110");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001001111");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010000");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010001");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010010");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010011");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010100");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010101");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010110");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001010111");
        state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_13_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011000");
        IF ( COMP_LOOP_13_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_386;
        ELSE
          state_var_NS <= COMP_LOOP_13_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_386 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011001");
        state_var_NS <= COMP_LOOP_C_387;
      WHEN COMP_LOOP_C_387 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011010");
        state_var_NS <= COMP_LOOP_C_388;
      WHEN COMP_LOOP_C_388 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011011");
        state_var_NS <= COMP_LOOP_C_389;
      WHEN COMP_LOOP_C_389 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011100");
        state_var_NS <= COMP_LOOP_C_390;
      WHEN COMP_LOOP_C_390 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011101");
        state_var_NS <= COMP_LOOP_C_391;
      WHEN COMP_LOOP_C_391 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011110");
        state_var_NS <= COMP_LOOP_C_392;
      WHEN COMP_LOOP_C_392 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001011111");
        state_var_NS <= COMP_LOOP_C_393;
      WHEN COMP_LOOP_C_393 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100000");
        state_var_NS <= COMP_LOOP_C_394;
      WHEN COMP_LOOP_C_394 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100001");
        state_var_NS <= COMP_LOOP_C_395;
      WHEN COMP_LOOP_C_395 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100010");
        state_var_NS <= COMP_LOOP_C_396;
      WHEN COMP_LOOP_C_396 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100011");
        state_var_NS <= COMP_LOOP_C_397;
      WHEN COMP_LOOP_C_397 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100100");
        state_var_NS <= COMP_LOOP_C_398;
      WHEN COMP_LOOP_C_398 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100101");
        state_var_NS <= COMP_LOOP_C_399;
      WHEN COMP_LOOP_C_399 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100110");
        state_var_NS <= COMP_LOOP_C_400;
      WHEN COMP_LOOP_C_400 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001100111");
        state_var_NS <= COMP_LOOP_C_401;
      WHEN COMP_LOOP_C_401 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101000");
        state_var_NS <= COMP_LOOP_C_402;
      WHEN COMP_LOOP_C_402 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101001");
        state_var_NS <= COMP_LOOP_C_403;
      WHEN COMP_LOOP_C_403 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101010");
        state_var_NS <= COMP_LOOP_C_404;
      WHEN COMP_LOOP_C_404 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101011");
        state_var_NS <= COMP_LOOP_C_405;
      WHEN COMP_LOOP_C_405 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101100");
        state_var_NS <= COMP_LOOP_C_406;
      WHEN COMP_LOOP_C_406 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101101");
        state_var_NS <= COMP_LOOP_C_407;
      WHEN COMP_LOOP_C_407 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101110");
        state_var_NS <= COMP_LOOP_C_408;
      WHEN COMP_LOOP_C_408 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001101111");
        state_var_NS <= COMP_LOOP_C_409;
      WHEN COMP_LOOP_C_409 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110000");
        state_var_NS <= COMP_LOOP_C_410;
      WHEN COMP_LOOP_C_410 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110001");
        state_var_NS <= COMP_LOOP_C_411;
      WHEN COMP_LOOP_C_411 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110010");
        state_var_NS <= COMP_LOOP_C_412;
      WHEN COMP_LOOP_C_412 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110011");
        state_var_NS <= COMP_LOOP_C_413;
      WHEN COMP_LOOP_C_413 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110100");
        state_var_NS <= COMP_LOOP_C_414;
      WHEN COMP_LOOP_C_414 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110101");
        state_var_NS <= COMP_LOOP_C_415;
      WHEN COMP_LOOP_C_415 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110110");
        state_var_NS <= COMP_LOOP_C_416;
      WHEN COMP_LOOP_C_416 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001110111");
        IF ( COMP_LOOP_C_416_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_417;
        END IF;
      WHEN COMP_LOOP_C_417 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111000");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111001");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111010");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111011");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111100");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111101");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111110");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1001111111");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000000");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000001");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000010");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000011");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000100");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000101");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000110");
        state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_14_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010000111");
        IF ( COMP_LOOP_14_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_418;
        ELSE
          state_var_NS <= COMP_LOOP_14_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_418 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001000");
        state_var_NS <= COMP_LOOP_C_419;
      WHEN COMP_LOOP_C_419 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001001");
        state_var_NS <= COMP_LOOP_C_420;
      WHEN COMP_LOOP_C_420 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001010");
        state_var_NS <= COMP_LOOP_C_421;
      WHEN COMP_LOOP_C_421 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001011");
        state_var_NS <= COMP_LOOP_C_422;
      WHEN COMP_LOOP_C_422 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001100");
        state_var_NS <= COMP_LOOP_C_423;
      WHEN COMP_LOOP_C_423 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001101");
        state_var_NS <= COMP_LOOP_C_424;
      WHEN COMP_LOOP_C_424 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001110");
        state_var_NS <= COMP_LOOP_C_425;
      WHEN COMP_LOOP_C_425 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010001111");
        state_var_NS <= COMP_LOOP_C_426;
      WHEN COMP_LOOP_C_426 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010000");
        state_var_NS <= COMP_LOOP_C_427;
      WHEN COMP_LOOP_C_427 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010001");
        state_var_NS <= COMP_LOOP_C_428;
      WHEN COMP_LOOP_C_428 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010010");
        state_var_NS <= COMP_LOOP_C_429;
      WHEN COMP_LOOP_C_429 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010011");
        state_var_NS <= COMP_LOOP_C_430;
      WHEN COMP_LOOP_C_430 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010100");
        state_var_NS <= COMP_LOOP_C_431;
      WHEN COMP_LOOP_C_431 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010101");
        state_var_NS <= COMP_LOOP_C_432;
      WHEN COMP_LOOP_C_432 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010110");
        state_var_NS <= COMP_LOOP_C_433;
      WHEN COMP_LOOP_C_433 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010010111");
        state_var_NS <= COMP_LOOP_C_434;
      WHEN COMP_LOOP_C_434 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011000");
        state_var_NS <= COMP_LOOP_C_435;
      WHEN COMP_LOOP_C_435 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011001");
        state_var_NS <= COMP_LOOP_C_436;
      WHEN COMP_LOOP_C_436 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011010");
        state_var_NS <= COMP_LOOP_C_437;
      WHEN COMP_LOOP_C_437 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011011");
        state_var_NS <= COMP_LOOP_C_438;
      WHEN COMP_LOOP_C_438 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011100");
        state_var_NS <= COMP_LOOP_C_439;
      WHEN COMP_LOOP_C_439 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011101");
        state_var_NS <= COMP_LOOP_C_440;
      WHEN COMP_LOOP_C_440 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011110");
        state_var_NS <= COMP_LOOP_C_441;
      WHEN COMP_LOOP_C_441 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010011111");
        state_var_NS <= COMP_LOOP_C_442;
      WHEN COMP_LOOP_C_442 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100000");
        state_var_NS <= COMP_LOOP_C_443;
      WHEN COMP_LOOP_C_443 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100001");
        state_var_NS <= COMP_LOOP_C_444;
      WHEN COMP_LOOP_C_444 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100010");
        state_var_NS <= COMP_LOOP_C_445;
      WHEN COMP_LOOP_C_445 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100011");
        state_var_NS <= COMP_LOOP_C_446;
      WHEN COMP_LOOP_C_446 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100100");
        state_var_NS <= COMP_LOOP_C_447;
      WHEN COMP_LOOP_C_447 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100101");
        state_var_NS <= COMP_LOOP_C_448;
      WHEN COMP_LOOP_C_448 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100110");
        IF ( COMP_LOOP_C_448_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_449;
        END IF;
      WHEN COMP_LOOP_C_449 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010100111");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101000");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101001");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101010");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101011");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101100");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101101");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101110");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010101111");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110000");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110001");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110010");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110011");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110100");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110101");
        state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_15_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110110");
        IF ( COMP_LOOP_15_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_450;
        ELSE
          state_var_NS <= COMP_LOOP_15_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_450 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010110111");
        state_var_NS <= COMP_LOOP_C_451;
      WHEN COMP_LOOP_C_451 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111000");
        state_var_NS <= COMP_LOOP_C_452;
      WHEN COMP_LOOP_C_452 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111001");
        state_var_NS <= COMP_LOOP_C_453;
      WHEN COMP_LOOP_C_453 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111010");
        state_var_NS <= COMP_LOOP_C_454;
      WHEN COMP_LOOP_C_454 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111011");
        state_var_NS <= COMP_LOOP_C_455;
      WHEN COMP_LOOP_C_455 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111100");
        state_var_NS <= COMP_LOOP_C_456;
      WHEN COMP_LOOP_C_456 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111101");
        state_var_NS <= COMP_LOOP_C_457;
      WHEN COMP_LOOP_C_457 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111110");
        state_var_NS <= COMP_LOOP_C_458;
      WHEN COMP_LOOP_C_458 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1010111111");
        state_var_NS <= COMP_LOOP_C_459;
      WHEN COMP_LOOP_C_459 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000000");
        state_var_NS <= COMP_LOOP_C_460;
      WHEN COMP_LOOP_C_460 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000001");
        state_var_NS <= COMP_LOOP_C_461;
      WHEN COMP_LOOP_C_461 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000010");
        state_var_NS <= COMP_LOOP_C_462;
      WHEN COMP_LOOP_C_462 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000011");
        state_var_NS <= COMP_LOOP_C_463;
      WHEN COMP_LOOP_C_463 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000100");
        state_var_NS <= COMP_LOOP_C_464;
      WHEN COMP_LOOP_C_464 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000101");
        state_var_NS <= COMP_LOOP_C_465;
      WHEN COMP_LOOP_C_465 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000110");
        state_var_NS <= COMP_LOOP_C_466;
      WHEN COMP_LOOP_C_466 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011000111");
        state_var_NS <= COMP_LOOP_C_467;
      WHEN COMP_LOOP_C_467 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001000");
        state_var_NS <= COMP_LOOP_C_468;
      WHEN COMP_LOOP_C_468 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001001");
        state_var_NS <= COMP_LOOP_C_469;
      WHEN COMP_LOOP_C_469 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001010");
        state_var_NS <= COMP_LOOP_C_470;
      WHEN COMP_LOOP_C_470 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001011");
        state_var_NS <= COMP_LOOP_C_471;
      WHEN COMP_LOOP_C_471 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001100");
        state_var_NS <= COMP_LOOP_C_472;
      WHEN COMP_LOOP_C_472 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001101");
        state_var_NS <= COMP_LOOP_C_473;
      WHEN COMP_LOOP_C_473 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001110");
        state_var_NS <= COMP_LOOP_C_474;
      WHEN COMP_LOOP_C_474 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011001111");
        state_var_NS <= COMP_LOOP_C_475;
      WHEN COMP_LOOP_C_475 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010000");
        state_var_NS <= COMP_LOOP_C_476;
      WHEN COMP_LOOP_C_476 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010001");
        state_var_NS <= COMP_LOOP_C_477;
      WHEN COMP_LOOP_C_477 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010010");
        state_var_NS <= COMP_LOOP_C_478;
      WHEN COMP_LOOP_C_478 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010011");
        state_var_NS <= COMP_LOOP_C_479;
      WHEN COMP_LOOP_C_479 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010100");
        state_var_NS <= COMP_LOOP_C_480;
      WHEN COMP_LOOP_C_480 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010101");
        IF ( COMP_LOOP_C_480_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_481;
        END IF;
      WHEN COMP_LOOP_C_481 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010110");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_0;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011010111");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_1;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011000");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_2;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011001");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_3;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011010");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_4;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011011");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_5;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011100");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_6;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011101");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_7;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011110");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_8;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011011111");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_9;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100000");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_10;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100001");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_11;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100010");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_12;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100011");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_13;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100100");
        state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_14;
      WHEN COMP_LOOP_16_modExp_dev_1_while_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100101");
        IF ( COMP_LOOP_16_modExp_dev_1_while_C_14_tr0 = '1' ) THEN
          state_var_NS <= COMP_LOOP_C_482;
        ELSE
          state_var_NS <= COMP_LOOP_16_modExp_dev_1_while_C_0;
        END IF;
      WHEN COMP_LOOP_C_482 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100110");
        state_var_NS <= COMP_LOOP_C_483;
      WHEN COMP_LOOP_C_483 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011100111");
        state_var_NS <= COMP_LOOP_C_484;
      WHEN COMP_LOOP_C_484 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101000");
        state_var_NS <= COMP_LOOP_C_485;
      WHEN COMP_LOOP_C_485 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101001");
        state_var_NS <= COMP_LOOP_C_486;
      WHEN COMP_LOOP_C_486 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101010");
        state_var_NS <= COMP_LOOP_C_487;
      WHEN COMP_LOOP_C_487 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101011");
        state_var_NS <= COMP_LOOP_C_488;
      WHEN COMP_LOOP_C_488 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101100");
        state_var_NS <= COMP_LOOP_C_489;
      WHEN COMP_LOOP_C_489 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101101");
        state_var_NS <= COMP_LOOP_C_490;
      WHEN COMP_LOOP_C_490 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101110");
        state_var_NS <= COMP_LOOP_C_491;
      WHEN COMP_LOOP_C_491 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011101111");
        state_var_NS <= COMP_LOOP_C_492;
      WHEN COMP_LOOP_C_492 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110000");
        state_var_NS <= COMP_LOOP_C_493;
      WHEN COMP_LOOP_C_493 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110001");
        state_var_NS <= COMP_LOOP_C_494;
      WHEN COMP_LOOP_C_494 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110010");
        state_var_NS <= COMP_LOOP_C_495;
      WHEN COMP_LOOP_C_495 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110011");
        state_var_NS <= COMP_LOOP_C_496;
      WHEN COMP_LOOP_C_496 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110100");
        state_var_NS <= COMP_LOOP_C_497;
      WHEN COMP_LOOP_C_497 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110101");
        state_var_NS <= COMP_LOOP_C_498;
      WHEN COMP_LOOP_C_498 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110110");
        state_var_NS <= COMP_LOOP_C_499;
      WHEN COMP_LOOP_C_499 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011110111");
        state_var_NS <= COMP_LOOP_C_500;
      WHEN COMP_LOOP_C_500 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111000");
        state_var_NS <= COMP_LOOP_C_501;
      WHEN COMP_LOOP_C_501 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111001");
        state_var_NS <= COMP_LOOP_C_502;
      WHEN COMP_LOOP_C_502 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111010");
        state_var_NS <= COMP_LOOP_C_503;
      WHEN COMP_LOOP_C_503 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111011");
        state_var_NS <= COMP_LOOP_C_504;
      WHEN COMP_LOOP_C_504 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111100");
        state_var_NS <= COMP_LOOP_C_505;
      WHEN COMP_LOOP_C_505 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111101");
        state_var_NS <= COMP_LOOP_C_506;
      WHEN COMP_LOOP_C_506 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111110");
        state_var_NS <= COMP_LOOP_C_507;
      WHEN COMP_LOOP_C_507 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1011111111");
        state_var_NS <= COMP_LOOP_C_508;
      WHEN COMP_LOOP_C_508 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000000");
        state_var_NS <= COMP_LOOP_C_509;
      WHEN COMP_LOOP_C_509 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000001");
        state_var_NS <= COMP_LOOP_C_510;
      WHEN COMP_LOOP_C_510 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000010");
        state_var_NS <= COMP_LOOP_C_511;
      WHEN COMP_LOOP_C_511 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000011");
        state_var_NS <= COMP_LOOP_C_512;
      WHEN COMP_LOOP_C_512 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000100");
        IF ( COMP_LOOP_C_512_tr0 = '1' ) THEN
          state_var_NS <= VEC_LOOP_C_0;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN VEC_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000101");
        IF ( VEC_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_4;
        ELSE
          state_var_NS <= COMP_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000110");
        IF ( STAGE_LOOP_C_4_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1100000111");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS inPlaceNTT_DIT_core_core_fsm_1;

  inPlaceNTT_DIT_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS inPlaceNTT_DIT_core_core_fsm_1_REG;

END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core_wait_dp IS
  PORT(
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    modulo_dev_cmp_ccs_ccore_en : OUT STD_LOGIC
  );
END inPlaceNTT_DIT_core_wait_dp;

ARCHITECTURE v11 OF inPlaceNTT_DIT_core_wait_dp IS
  -- Default Constants

BEGIN
  modulo_dev_cmp_ccs_ccore_en <= ensig_cgo OR ensig_cgo_iro;
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    vec_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    vec_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_1_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_2_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_3_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_4_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_5_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_6_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_7_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_8_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_9_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_10_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_11_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_12_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_13_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_14_i_we_d_pff : OUT STD_LOGIC;
    vec_rsc_0_15_i_we_d_pff : OUT STD_LOGIC
  );
END inPlaceNTT_DIT_core;

ARCHITECTURE v11 OF inPlaceNTT_DIT_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_cmp_return_rsc_z : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_cmp_ccs_ccore_en : STD_LOGIC;
  SIGNAL operator_66_true_div_cmp_a : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_z : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_b_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL nand_tmp : STD_LOGIC;
  SIGNAL or_tmp_20 : STD_LOGIC;
  SIGNAL nor_tmp_14 : STD_LOGIC;
  SIGNAL or_tmp_74 : STD_LOGIC;
  SIGNAL nor_tmp_40 : STD_LOGIC;
  SIGNAL and_dcpl_13 : STD_LOGIC;
  SIGNAL and_dcpl_14 : STD_LOGIC;
  SIGNAL and_dcpl_15 : STD_LOGIC;
  SIGNAL and_dcpl_16 : STD_LOGIC;
  SIGNAL and_dcpl_17 : STD_LOGIC;
  SIGNAL and_dcpl_18 : STD_LOGIC;
  SIGNAL and_dcpl_19 : STD_LOGIC;
  SIGNAL and_dcpl_23 : STD_LOGIC;
  SIGNAL not_tmp_121 : STD_LOGIC;
  SIGNAL and_dcpl_26 : STD_LOGIC;
  SIGNAL and_dcpl_27 : STD_LOGIC;
  SIGNAL and_dcpl_28 : STD_LOGIC;
  SIGNAL and_dcpl_29 : STD_LOGIC;
  SIGNAL and_dcpl_30 : STD_LOGIC;
  SIGNAL and_dcpl_32 : STD_LOGIC;
  SIGNAL and_dcpl_33 : STD_LOGIC;
  SIGNAL and_dcpl_34 : STD_LOGIC;
  SIGNAL and_dcpl_35 : STD_LOGIC;
  SIGNAL and_dcpl_36 : STD_LOGIC;
  SIGNAL and_dcpl_37 : STD_LOGIC;
  SIGNAL and_dcpl_38 : STD_LOGIC;
  SIGNAL and_dcpl_39 : STD_LOGIC;
  SIGNAL and_dcpl_40 : STD_LOGIC;
  SIGNAL and_dcpl_42 : STD_LOGIC;
  SIGNAL and_dcpl_43 : STD_LOGIC;
  SIGNAL and_dcpl_44 : STD_LOGIC;
  SIGNAL and_dcpl_45 : STD_LOGIC;
  SIGNAL and_dcpl_47 : STD_LOGIC;
  SIGNAL and_dcpl_48 : STD_LOGIC;
  SIGNAL and_dcpl_49 : STD_LOGIC;
  SIGNAL and_dcpl_50 : STD_LOGIC;
  SIGNAL and_dcpl_51 : STD_LOGIC;
  SIGNAL and_dcpl_52 : STD_LOGIC;
  SIGNAL and_dcpl_54 : STD_LOGIC;
  SIGNAL and_dcpl_55 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_58 : STD_LOGIC;
  SIGNAL and_dcpl_59 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_61 : STD_LOGIC;
  SIGNAL and_dcpl_63 : STD_LOGIC;
  SIGNAL and_dcpl_64 : STD_LOGIC;
  SIGNAL and_dcpl_65 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_68 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL and_dcpl_71 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_73 : STD_LOGIC;
  SIGNAL and_dcpl_74 : STD_LOGIC;
  SIGNAL and_dcpl_75 : STD_LOGIC;
  SIGNAL and_dcpl_78 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL and_dcpl_80 : STD_LOGIC;
  SIGNAL and_dcpl_81 : STD_LOGIC;
  SIGNAL and_dcpl_83 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_85 : STD_LOGIC;
  SIGNAL and_dcpl_86 : STD_LOGIC;
  SIGNAL and_dcpl_87 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_90 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_93 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_95 : STD_LOGIC;
  SIGNAL and_dcpl_97 : STD_LOGIC;
  SIGNAL and_dcpl_98 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL and_dcpl_101 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_106 : STD_LOGIC;
  SIGNAL and_dcpl_107 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_116 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL or_tmp_237 : STD_LOGIC;
  SIGNAL nand_tmp_6 : STD_LOGIC;
  SIGNAL or_tmp_239 : STD_LOGIC;
  SIGNAL or_tmp_241 : STD_LOGIC;
  SIGNAL nand_tmp_7 : STD_LOGIC;
  SIGNAL and_dcpl_122 : STD_LOGIC;
  SIGNAL and_dcpl_130 : STD_LOGIC;
  SIGNAL and_dcpl_132 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_138 : STD_LOGIC;
  SIGNAL or_tmp_252 : STD_LOGIC;
  SIGNAL or_tmp_253 : STD_LOGIC;
  SIGNAL or_tmp_258 : STD_LOGIC;
  SIGNAL or_tmp_259 : STD_LOGIC;
  SIGNAL not_tmp_133 : STD_LOGIC;
  SIGNAL not_tmp_134 : STD_LOGIC;
  SIGNAL or_tmp_346 : STD_LOGIC;
  SIGNAL or_tmp_352 : STD_LOGIC;
  SIGNAL or_tmp_353 : STD_LOGIC;
  SIGNAL or_tmp_362 : STD_LOGIC;
  SIGNAL or_tmp_438 : STD_LOGIC;
  SIGNAL or_tmp_439 : STD_LOGIC;
  SIGNAL or_tmp_444 : STD_LOGIC;
  SIGNAL or_tmp_445 : STD_LOGIC;
  SIGNAL or_tmp_531 : STD_LOGIC;
  SIGNAL or_tmp_532 : STD_LOGIC;
  SIGNAL or_tmp_537 : STD_LOGIC;
  SIGNAL or_tmp_538 : STD_LOGIC;
  SIGNAL or_tmp_624 : STD_LOGIC;
  SIGNAL or_tmp_625 : STD_LOGIC;
  SIGNAL or_tmp_630 : STD_LOGIC;
  SIGNAL or_tmp_631 : STD_LOGIC;
  SIGNAL or_tmp_718 : STD_LOGIC;
  SIGNAL or_tmp_724 : STD_LOGIC;
  SIGNAL or_tmp_725 : STD_LOGIC;
  SIGNAL or_tmp_734 : STD_LOGIC;
  SIGNAL or_tmp_810 : STD_LOGIC;
  SIGNAL or_tmp_811 : STD_LOGIC;
  SIGNAL or_tmp_816 : STD_LOGIC;
  SIGNAL or_tmp_817 : STD_LOGIC;
  SIGNAL or_tmp_903 : STD_LOGIC;
  SIGNAL or_tmp_904 : STD_LOGIC;
  SIGNAL or_tmp_909 : STD_LOGIC;
  SIGNAL or_tmp_910 : STD_LOGIC;
  SIGNAL or_tmp_997 : STD_LOGIC;
  SIGNAL or_tmp_999 : STD_LOGIC;
  SIGNAL or_tmp_1005 : STD_LOGIC;
  SIGNAL or_tmp_1007 : STD_LOGIC;
  SIGNAL or_tmp_1097 : STD_LOGIC;
  SIGNAL or_tmp_1104 : STD_LOGIC;
  SIGNAL or_tmp_1106 : STD_LOGIC;
  SIGNAL or_tmp_1116 : STD_LOGIC;
  SIGNAL or_tmp_1195 : STD_LOGIC;
  SIGNAL or_tmp_1197 : STD_LOGIC;
  SIGNAL or_tmp_1203 : STD_LOGIC;
  SIGNAL or_tmp_1205 : STD_LOGIC;
  SIGNAL or_tmp_1294 : STD_LOGIC;
  SIGNAL or_tmp_1296 : STD_LOGIC;
  SIGNAL or_tmp_1302 : STD_LOGIC;
  SIGNAL or_tmp_1304 : STD_LOGIC;
  SIGNAL not_tmp_289 : STD_LOGIC;
  SIGNAL or_tmp_1393 : STD_LOGIC;
  SIGNAL or_tmp_1395 : STD_LOGIC;
  SIGNAL or_tmp_1401 : STD_LOGIC;
  SIGNAL or_tmp_1403 : STD_LOGIC;
  SIGNAL not_tmp_304 : STD_LOGIC;
  SIGNAL or_tmp_1493 : STD_LOGIC;
  SIGNAL or_tmp_1500 : STD_LOGIC;
  SIGNAL or_tmp_1502 : STD_LOGIC;
  SIGNAL or_tmp_1512 : STD_LOGIC;
  SIGNAL or_tmp_1590 : STD_LOGIC;
  SIGNAL or_tmp_1592 : STD_LOGIC;
  SIGNAL or_tmp_1598 : STD_LOGIC;
  SIGNAL or_tmp_1600 : STD_LOGIC;
  SIGNAL not_tmp_335 : STD_LOGIC;
  SIGNAL or_tmp_1687 : STD_LOGIC;
  SIGNAL or_tmp_1689 : STD_LOGIC;
  SIGNAL not_tmp_336 : STD_LOGIC;
  SIGNAL or_tmp_1694 : STD_LOGIC;
  SIGNAL nor_tmp_186 : STD_LOGIC;
  SIGNAL mux_tmp_1470 : STD_LOGIC;
  SIGNAL mux_tmp_1471 : STD_LOGIC;
  SIGNAL mux_tmp_1472 : STD_LOGIC;
  SIGNAL mux_tmp_1473 : STD_LOGIC;
  SIGNAL mux_tmp_1476 : STD_LOGIC;
  SIGNAL nor_tmp_188 : STD_LOGIC;
  SIGNAL mux_tmp_1477 : STD_LOGIC;
  SIGNAL nor_tmp_190 : STD_LOGIC;
  SIGNAL mux_tmp_1482 : STD_LOGIC;
  SIGNAL mux_tmp_1483 : STD_LOGIC;
  SIGNAL mux_tmp_1484 : STD_LOGIC;
  SIGNAL mux_tmp_1485 : STD_LOGIC;
  SIGNAL mux_tmp_1488 : STD_LOGIC;
  SIGNAL mux_tmp_1489 : STD_LOGIC;
  SIGNAL mux_tmp_1496 : STD_LOGIC;
  SIGNAL mux_tmp_1498 : STD_LOGIC;
  SIGNAL mux_tmp_1501 : STD_LOGIC;
  SIGNAL mux_tmp_1503 : STD_LOGIC;
  SIGNAL mux_tmp_1514 : STD_LOGIC;
  SIGNAL or_tmp_1788 : STD_LOGIC;
  SIGNAL or_tmp_1793 : STD_LOGIC;
  SIGNAL or_tmp_1794 : STD_LOGIC;
  SIGNAL mux_tmp_1534 : STD_LOGIC;
  SIGNAL or_tmp_1796 : STD_LOGIC;
  SIGNAL mux_tmp_1537 : STD_LOGIC;
  SIGNAL or_tmp_1799 : STD_LOGIC;
  SIGNAL nand_tmp_106 : STD_LOGIC;
  SIGNAL not_tmp_370 : STD_LOGIC;
  SIGNAL or_tmp_1816 : STD_LOGIC;
  SIGNAL or_tmp_1818 : STD_LOGIC;
  SIGNAL mux_tmp_1562 : STD_LOGIC;
  SIGNAL mux_tmp_1563 : STD_LOGIC;
  SIGNAL or_tmp_1823 : STD_LOGIC;
  SIGNAL or_tmp_1824 : STD_LOGIC;
  SIGNAL mux_tmp_1566 : STD_LOGIC;
  SIGNAL or_tmp_1825 : STD_LOGIC;
  SIGNAL or_tmp_1827 : STD_LOGIC;
  SIGNAL or_tmp_1830 : STD_LOGIC;
  SIGNAL or_tmp_1831 : STD_LOGIC;
  SIGNAL mux_tmp_1573 : STD_LOGIC;
  SIGNAL or_tmp_1835 : STD_LOGIC;
  SIGNAL mux_tmp_1579 : STD_LOGIC;
  SIGNAL or_tmp_1838 : STD_LOGIC;
  SIGNAL or_tmp_1840 : STD_LOGIC;
  SIGNAL or_tmp_1841 : STD_LOGIC;
  SIGNAL and_dcpl_169 : STD_LOGIC;
  SIGNAL or_tmp_1845 : STD_LOGIC;
  SIGNAL and_tmp_12 : STD_LOGIC;
  SIGNAL mux_tmp_1610 : STD_LOGIC;
  SIGNAL mux_tmp_1612 : STD_LOGIC;
  SIGNAL or_tmp_1854 : STD_LOGIC;
  SIGNAL mux_tmp_1615 : STD_LOGIC;
  SIGNAL or_tmp_1855 : STD_LOGIC;
  SIGNAL mux_tmp_1618 : STD_LOGIC;
  SIGNAL mux_tmp_1621 : STD_LOGIC;
  SIGNAL mux_tmp_1623 : STD_LOGIC;
  SIGNAL mux_tmp_1625 : STD_LOGIC;
  SIGNAL mux_tmp_1626 : STD_LOGIC;
  SIGNAL mux_tmp_1629 : STD_LOGIC;
  SIGNAL mux_tmp_1688 : STD_LOGIC;
  SIGNAL or_tmp_1899 : STD_LOGIC;
  SIGNAL and_dcpl_183 : STD_LOGIC;
  SIGNAL not_tmp_402 : STD_LOGIC;
  SIGNAL nor_tmp_203 : STD_LOGIC;
  SIGNAL not_tmp_418 : STD_LOGIC;
  SIGNAL or_tmp_1989 : STD_LOGIC;
  SIGNAL or_tmp_1990 : STD_LOGIC;
  SIGNAL mux_tmp_1782 : STD_LOGIC;
  SIGNAL mux_tmp_1786 : STD_LOGIC;
  SIGNAL mux_tmp_1793 : STD_LOGIC;
  SIGNAL mux_tmp_1799 : STD_LOGIC;
  SIGNAL mux_tmp_1801 : STD_LOGIC;
  SIGNAL mux_tmp_1803 : STD_LOGIC;
  SIGNAL mux_tmp_1808 : STD_LOGIC;
  SIGNAL mux_tmp_1809 : STD_LOGIC;
  SIGNAL not_tmp_431 : STD_LOGIC;
  SIGNAL nor_tmp_215 : STD_LOGIC;
  SIGNAL not_tmp_439 : STD_LOGIC;
  SIGNAL mux_tmp_1839 : STD_LOGIC;
  SIGNAL and_dcpl_199 : STD_LOGIC;
  SIGNAL and_dcpl_200 : STD_LOGIC;
  SIGNAL and_dcpl_201 : STD_LOGIC;
  SIGNAL and_dcpl_202 : STD_LOGIC;
  SIGNAL and_dcpl_203 : STD_LOGIC;
  SIGNAL and_dcpl_204 : STD_LOGIC;
  SIGNAL and_dcpl_206 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL and_dcpl_208 : STD_LOGIC;
  SIGNAL and_dcpl_210 : STD_LOGIC;
  SIGNAL and_dcpl_212 : STD_LOGIC;
  SIGNAL and_dcpl_214 : STD_LOGIC;
  SIGNAL and_dcpl_215 : STD_LOGIC;
  SIGNAL and_dcpl_217 : STD_LOGIC;
  SIGNAL and_dcpl_219 : STD_LOGIC;
  SIGNAL and_dcpl_220 : STD_LOGIC;
  SIGNAL and_dcpl_221 : STD_LOGIC;
  SIGNAL or_tmp_2035 : STD_LOGIC;
  SIGNAL mux_tmp_1861 : STD_LOGIC;
  SIGNAL or_tmp_2037 : STD_LOGIC;
  SIGNAL mux_tmp_1863 : STD_LOGIC;
  SIGNAL or_tmp_2040 : STD_LOGIC;
  SIGNAL or_tmp_2041 : STD_LOGIC;
  SIGNAL mux_tmp_1866 : STD_LOGIC;
  SIGNAL or_tmp_2043 : STD_LOGIC;
  SIGNAL or_tmp_2044 : STD_LOGIC;
  SIGNAL mux_tmp_1870 : STD_LOGIC;
  SIGNAL mux_tmp_1872 : STD_LOGIC;
  SIGNAL or_tmp_2047 : STD_LOGIC;
  SIGNAL mux_tmp_1874 : STD_LOGIC;
  SIGNAL mux_tmp_1875 : STD_LOGIC;
  SIGNAL nand_tmp_134 : STD_LOGIC;
  SIGNAL mux_tmp_1876 : STD_LOGIC;
  SIGNAL mux_tmp_1877 : STD_LOGIC;
  SIGNAL mux_tmp_1882 : STD_LOGIC;
  SIGNAL mux_tmp_1883 : STD_LOGIC;
  SIGNAL mux_tmp_1888 : STD_LOGIC;
  SIGNAL mux_tmp_1891 : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_itm : STD_LOGIC;
  SIGNAL VEC_LOOP_acc_1_psp_1 : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_nor_11_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_13_psp_sva_1 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_k_9_4_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL VEC_LOOP_j_sva_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_acc_1_cse_6_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_13_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_4_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_11_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_14_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_19_psp_sva : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_12_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_17_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_10_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_16_psp_sva : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_8_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_14_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_20_psp_sva : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_1_cse_2_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL nand_308_cse : STD_LOGIC;
  SIGNAL nand_264_cse : STD_LOGIC;
  SIGNAL reg_vec_rsc_triosy_0_15_obj_ld_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL or_1973_cse : STD_LOGIC;
  SIGNAL nor_256_cse : STD_LOGIC;
  SIGNAL or_1916_cse : STD_LOGIC;
  SIGNAL and_267_cse : STD_LOGIC;
  SIGNAL or_2186_cse : STD_LOGIC;
  SIGNAL and_418_cse : STD_LOGIC;
  SIGNAL or_2040_cse : STD_LOGIC;
  SIGNAL or_1982_cse : STD_LOGIC;
  SIGNAL or_1967_cse : STD_LOGIC;
  SIGNAL or_214_cse : STD_LOGIC;
  SIGNAL nor_697_cse : STD_LOGIC;
  SIGNAL or_279_cse : STD_LOGIC;
  SIGNAL or_1977_cse : STD_LOGIC;
  SIGNAL and_375_cse : STD_LOGIC;
  SIGNAL mux_424_cse : STD_LOGIC;
  SIGNAL or_212_cse : STD_LOGIC;
  SIGNAL nand_321_cse : STD_LOGIC;
  SIGNAL and_247_cse : STD_LOGIC;
  SIGNAL or_2151_cse : STD_LOGIC;
  SIGNAL and_376_cse : STD_LOGIC;
  SIGNAL nor_728_cse : STD_LOGIC;
  SIGNAL or_1820_cse : STD_LOGIC;
  SIGNAL or_2012_cse : STD_LOGIC;
  SIGNAL or_103_cse : STD_LOGIC;
  SIGNAL nand_357_cse : STD_LOGIC;
  SIGNAL mux_1802_cse : STD_LOGIC;
  SIGNAL mux_1788_cse : STD_LOGIC;
  SIGNAL mux_1797_cse : STD_LOGIC;
  SIGNAL mux_461_cse : STD_LOGIC;
  SIGNAL mux_460_cse : STD_LOGIC;
  SIGNAL mux_1789_cse : STD_LOGIC;
  SIGNAL mux_1583_cse : STD_LOGIC;
  SIGNAL mux_1784_cse : STD_LOGIC;
  SIGNAL or_1880_cse : STD_LOGIC;
  SIGNAL nor_760_cse : STD_LOGIC;
  SIGNAL mux_1602_cse : STD_LOGIC;
  SIGNAL mux_1785_cse : STD_LOGIC;
  SIGNAL and_259_cse : STD_LOGIC;
  SIGNAL mux_1726_cse : STD_LOGIC;
  SIGNAL mux_1909_cse : STD_LOGIC;
  SIGNAL mux_1911_cse : STD_LOGIC;
  SIGNAL COMP_LOOP_1_mul_itm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL tmp_10_lpi_4_dfm : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_psp_sva : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL mux_1581_itm : STD_LOGIC;
  SIGNAL mux_1832_itm : STD_LOGIC;
  SIGNAL mux_1834_itm : STD_LOGIC;
  SIGNAL mux_tmp_2006 : STD_LOGIC;
  SIGNAL and_dcpl_231 : STD_LOGIC;
  SIGNAL and_dcpl_232 : STD_LOGIC;
  SIGNAL and_dcpl_233 : STD_LOGIC;
  SIGNAL and_dcpl_234 : STD_LOGIC;
  SIGNAL and_dcpl_236 : STD_LOGIC;
  SIGNAL and_dcpl_237 : STD_LOGIC;
  SIGNAL and_dcpl_238 : STD_LOGIC;
  SIGNAL and_dcpl_242 : STD_LOGIC;
  SIGNAL and_dcpl_243 : STD_LOGIC;
  SIGNAL and_dcpl_244 : STD_LOGIC;
  SIGNAL and_dcpl_246 : STD_LOGIC;
  SIGNAL and_dcpl_248 : STD_LOGIC;
  SIGNAL and_dcpl_250 : STD_LOGIC;
  SIGNAL and_dcpl_251 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL and_dcpl_255 : STD_LOGIC;
  SIGNAL and_dcpl_256 : STD_LOGIC;
  SIGNAL and_dcpl_260 : STD_LOGIC;
  SIGNAL and_dcpl_265 : STD_LOGIC;
  SIGNAL and_dcpl_267 : STD_LOGIC;
  SIGNAL and_dcpl_271 : STD_LOGIC;
  SIGNAL and_dcpl_272 : STD_LOGIC;
  SIGNAL and_dcpl_274 : STD_LOGIC;
  SIGNAL and_dcpl_277 : STD_LOGIC;
  SIGNAL and_dcpl_278 : STD_LOGIC;
  SIGNAL and_dcpl_279 : STD_LOGIC;
  SIGNAL and_dcpl_281 : STD_LOGIC;
  SIGNAL and_dcpl_284 : STD_LOGIC;
  SIGNAL z_out_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL and_dcpl_300 : STD_LOGIC;
  SIGNAL and_dcpl_308 : STD_LOGIC;
  SIGNAL z_out_2 : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL and_dcpl_344 : STD_LOGIC;
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL and_dcpl_361 : STD_LOGIC;
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL and_dcpl_376 : STD_LOGIC;
  SIGNAL and_dcpl_382 : STD_LOGIC;
  SIGNAL and_dcpl_396 : STD_LOGIC;
  SIGNAL and_dcpl_398 : STD_LOGIC;
  SIGNAL and_dcpl_402 : STD_LOGIC;
  SIGNAL and_dcpl_403 : STD_LOGIC;
  SIGNAL and_dcpl_406 : STD_LOGIC;
  SIGNAL and_dcpl_407 : STD_LOGIC;
  SIGNAL and_dcpl_416 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL and_dcpl_425 : STD_LOGIC;
  SIGNAL and_dcpl_444 : STD_LOGIC;
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL and_dcpl_460 : STD_LOGIC;
  SIGNAL and_dcpl_464 : STD_LOGIC;
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL r_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_psp_sva : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL modExp_dev_exp_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_dev_result_sva : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_2_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_4_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_5_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_6_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_8_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_9_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_11_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_13_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_14_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_nor_1_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_12_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_62_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_64_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_68_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_139_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_140_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_141_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_143_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_144_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_145_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_146_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_147_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_148_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_149_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_134_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_137_itm : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_244_itm : STD_LOGIC;
  SIGNAL modExp_dev_exp_1_sva_63_9 : STD_LOGIC_VECTOR (54 DOWNTO 0);
  SIGNAL modExp_dev_exp_1_sva_3_0 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_i_3_0_sva_mx0c1 : STD_LOGIC;
  SIGNAL STAGE_LOOP_lshift_psp_sva_mx0w0 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL VEC_LOOP_j_sva_9_0_mx0c1 : STD_LOGIC;
  SIGNAL and_195_rgt : STD_LOGIC;
  SIGNAL and_551_ssc : STD_LOGIC;
  SIGNAL nand_270_cse_1 : STD_LOGIC;
  SIGNAL nand_260_cse_1 : STD_LOGIC;
  SIGNAL modExp_dev_while_or_2_cse : STD_LOGIC;
  SIGNAL nor_678_cse : STD_LOGIC;
  SIGNAL or_368_cse : STD_LOGIC;
  SIGNAL or_369_cse : STD_LOGIC;
  SIGNAL nor_650_cse : STD_LOGIC;
  SIGNAL or_462_cse : STD_LOGIC;
  SIGNAL nor_624_cse : STD_LOGIC;
  SIGNAL or_554_cse : STD_LOGIC;
  SIGNAL or_555_cse : STD_LOGIC;
  SIGNAL nor_598_cse : STD_LOGIC;
  SIGNAL or_648_cse : STD_LOGIC;
  SIGNAL nor_572_cse : STD_LOGIC;
  SIGNAL or_740_cse : STD_LOGIC;
  SIGNAL or_741_cse : STD_LOGIC;
  SIGNAL nor_544_cse : STD_LOGIC;
  SIGNAL or_834_cse : STD_LOGIC;
  SIGNAL nor_518_cse : STD_LOGIC;
  SIGNAL or_926_cse : STD_LOGIC;
  SIGNAL or_927_cse : STD_LOGIC;
  SIGNAL nor_492_cse : STD_LOGIC;
  SIGNAL nand_280_cse : STD_LOGIC;
  SIGNAL nand_275_cse : STD_LOGIC;
  SIGNAL nor_467_cse : STD_LOGIC;
  SIGNAL or_1119_cse : STD_LOGIC;
  SIGNAL nor_439_cse : STD_LOGIC;
  SIGNAL or_1218_cse : STD_LOGIC;
  SIGNAL nor_413_cse : STD_LOGIC;
  SIGNAL or_1317_cse : STD_LOGIC;
  SIGNAL nor_387_cse : STD_LOGIC;
  SIGNAL nand_241_cse : STD_LOGIC;
  SIGNAL nor_362_cse : STD_LOGIC;
  SIGNAL or_1515_cse : STD_LOGIC;
  SIGNAL nor_335_cse : STD_LOGIC;
  SIGNAL nand_217_cse : STD_LOGIC;
  SIGNAL nor_310_cse : STD_LOGIC;
  SIGNAL nand_202_cse : STD_LOGIC;
  SIGNAL nand_197_cse : STD_LOGIC;
  SIGNAL and_291_cse : STD_LOGIC;
  SIGNAL nand_161_cse : STD_LOGIC;
  SIGNAL nand_160_cse : STD_LOGIC;
  SIGNAL or_1995_cse : STD_LOGIC;
  SIGNAL or_1976_cse : STD_LOGIC;
  SIGNAL mux_1768_cse : STD_LOGIC;
  SIGNAL mux_2066_cse : STD_LOGIC;
  SIGNAL nand_tmp_139 : STD_LOGIC;
  SIGNAL or_tmp_2154 : STD_LOGIC;
  SIGNAL mux_tmp_2041 : STD_LOGIC;
  SIGNAL or_tmp_2156 : STD_LOGIC;
  SIGNAL mux_tmp_2043 : STD_LOGIC;
  SIGNAL mux_tmp_2046 : STD_LOGIC;
  SIGNAL or_tmp_2166 : STD_LOGIC;
  SIGNAL or_tmp_2168 : STD_LOGIC;
  SIGNAL mux_tmp_2052 : STD_LOGIC;
  SIGNAL or_tmp_2171 : STD_LOGIC;
  SIGNAL mux_tmp_2058 : STD_LOGIC;
  SIGNAL or_tmp_2183 : STD_LOGIC;
  SIGNAL mux_tmp_2072 : STD_LOGIC;
  SIGNAL not_tmp_571 : STD_LOGIC;
  SIGNAL or_tmp_2191 : STD_LOGIC;
  SIGNAL or_tmp_2193 : STD_LOGIC;
  SIGNAL mux_tmp_2081 : STD_LOGIC;
  SIGNAL mux_tmp_2083 : STD_LOGIC;
  SIGNAL operator_64_false_operator_64_false_mux_rgt : STD_LOGIC_VECTOR (64 DOWNTO
      0);
  SIGNAL mux_tmp_2108 : STD_LOGIC;
  SIGNAL or_tmp_2223 : STD_LOGIC;
  SIGNAL mux_tmp_2112 : STD_LOGIC;
  SIGNAL or_tmp_2227 : STD_LOGIC;
  SIGNAL mux_tmp_2119 : STD_LOGIC;
  SIGNAL mux_tmp_2124 : STD_LOGIC;
  SIGNAL mux_tmp_2128 : STD_LOGIC;
  SIGNAL or_tmp_2236 : STD_LOGIC;
  SIGNAL mux_tmp_2150 : STD_LOGIC;
  SIGNAL mux_tmp_2153 : STD_LOGIC;
  SIGNAL mux_tmp_2154 : STD_LOGIC;
  SIGNAL mux_tmp_2156 : STD_LOGIC;
  SIGNAL mux_tmp_2159 : STD_LOGIC;
  SIGNAL mux_tmp_2164 : STD_LOGIC;
  SIGNAL mux_tmp_2165 : STD_LOGIC;
  SIGNAL mux_tmp_2167 : STD_LOGIC;
  SIGNAL mux_tmp_2169 : STD_LOGIC;
  SIGNAL mux_tmp_2170 : STD_LOGIC;
  SIGNAL mux_tmp_2179 : STD_LOGIC;
  SIGNAL mux_tmp_2180 : STD_LOGIC;
  SIGNAL or_tmp_2243 : STD_LOGIC;
  SIGNAL or_tmp_2244 : STD_LOGIC;
  SIGNAL mux_tmp_2192 : STD_LOGIC;
  SIGNAL mux_tmp_2193 : STD_LOGIC;
  SIGNAL or_tmp_2245 : STD_LOGIC;
  SIGNAL mux_tmp_2196 : STD_LOGIC;
  SIGNAL mux_tmp_2199 : STD_LOGIC;
  SIGNAL mux_tmp_2204 : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_192_rgt : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_1_sva_9_5 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL COMP_LOOP_acc_10_cse_10_1_1_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL operator_64_false_acc_mut_64 : STD_LOGIC;
  SIGNAL operator_64_false_acc_mut_63_0 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL or_2306_cse : STD_LOGIC;
  SIGNAL or_2348_cse : STD_LOGIC;
  SIGNAL or_2336_cse : STD_LOGIC;
  SIGNAL nor_810_cse : STD_LOGIC;
  SIGNAL or_2086_cse : STD_LOGIC;
  SIGNAL or_2146_cse : STD_LOGIC;
  SIGNAL and_357_cse : STD_LOGIC;
  SIGNAL mux_1949_cse : STD_LOGIC;
  SIGNAL mux_1920_cse : STD_LOGIC;
  SIGNAL mux_1922_cse : STD_LOGIC;
  SIGNAL mux_1938_cse : STD_LOGIC;
  SIGNAL mux_2249_itm : STD_LOGIC;
  SIGNAL z_out_6_10_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL z_out_8_64_2 : STD_LOGIC_VECTOR (62 DOWNTO 0);
  SIGNAL nor_761_cse : STD_LOGIC;

  SIGNAL mux_1580_nl : STD_LOGIC;
  SIGNAL mux_1579_nl : STD_LOGIC;
  SIGNAL mux_1578_nl : STD_LOGIC;
  SIGNAL mux_1577_nl : STD_LOGIC;
  SIGNAL mux_1576_nl : STD_LOGIC;
  SIGNAL mux_1575_nl : STD_LOGIC;
  SIGNAL mux_1574_nl : STD_LOGIC;
  SIGNAL mux_1573_nl : STD_LOGIC;
  SIGNAL mux_1572_nl : STD_LOGIC;
  SIGNAL mux_1571_nl : STD_LOGIC;
  SIGNAL mux_1570_nl : STD_LOGIC;
  SIGNAL and_278_nl : STD_LOGIC;
  SIGNAL mux_1569_nl : STD_LOGIC;
  SIGNAL mux_1568_nl : STD_LOGIC;
  SIGNAL mux_1567_nl : STD_LOGIC;
  SIGNAL mux_1566_nl : STD_LOGIC;
  SIGNAL mux_1563_nl : STD_LOGIC;
  SIGNAL mux_1562_nl : STD_LOGIC;
  SIGNAL and_280_nl : STD_LOGIC;
  SIGNAL mux_1561_nl : STD_LOGIC;
  SIGNAL mux_1560_nl : STD_LOGIC;
  SIGNAL mux_1559_nl : STD_LOGIC;
  SIGNAL mux_1558_nl : STD_LOGIC;
  SIGNAL mux_1557_nl : STD_LOGIC;
  SIGNAL mux_1556_nl : STD_LOGIC;
  SIGNAL mux_1555_nl : STD_LOGIC;
  SIGNAL mux_1553_nl : STD_LOGIC;
  SIGNAL mux_1551_nl : STD_LOGIC;
  SIGNAL mux_1550_nl : STD_LOGIC;
  SIGNAL mux_1546_nl : STD_LOGIC;
  SIGNAL mux_1545_nl : STD_LOGIC;
  SIGNAL mux_1544_nl : STD_LOGIC;
  SIGNAL mux_1543_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL mux_1541_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL mux_1531_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL mux_1529_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL nor_271_nl : STD_LOGIC;
  SIGNAL or_1980_nl : STD_LOGIC;
  SIGNAL mux_1725_nl : STD_LOGIC;
  SIGNAL modExp_dev_while_mux1h_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL mul_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_dev_while_mux_2_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_dev_while_mux_3_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_1_acc_8_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modExp_dev_while_or_1_nl : STD_LOGIC;
  SIGNAL mux_1792_nl : STD_LOGIC;
  SIGNAL mux_1791_nl : STD_LOGIC;
  SIGNAL mux_1790_nl : STD_LOGIC;
  SIGNAL and_258_nl : STD_LOGIC;
  SIGNAL nor_255_nl : STD_LOGIC;
  SIGNAL mux_1787_nl : STD_LOGIC;
  SIGNAL mux_1786_nl : STD_LOGIC;
  SIGNAL and_260_nl : STD_LOGIC;
  SIGNAL nor_257_nl : STD_LOGIC;
  SIGNAL mux_1783_nl : STD_LOGIC;
  SIGNAL mux_1698_nl : STD_LOGIC;
  SIGNAL mux_1697_nl : STD_LOGIC;
  SIGNAL mux_1696_nl : STD_LOGIC;
  SIGNAL mux_1695_nl : STD_LOGIC;
  SIGNAL mux_1694_nl : STD_LOGIC;
  SIGNAL or_1896_nl : STD_LOGIC;
  SIGNAL mux_1693_nl : STD_LOGIC;
  SIGNAL mux_1692_nl : STD_LOGIC;
  SIGNAL mux_1691_nl : STD_LOGIC;
  SIGNAL mux_1690_nl : STD_LOGIC;
  SIGNAL mux_1689_nl : STD_LOGIC;
  SIGNAL mux_1688_nl : STD_LOGIC;
  SIGNAL mux_1727_nl : STD_LOGIC;
  SIGNAL mux_1686_nl : STD_LOGIC;
  SIGNAL mux_1685_nl : STD_LOGIC;
  SIGNAL mux_1684_nl : STD_LOGIC;
  SIGNAL mux_1683_nl : STD_LOGIC;
  SIGNAL mux_1678_nl : STD_LOGIC;
  SIGNAL mux_1713_nl : STD_LOGIC;
  SIGNAL mux_1673_nl : STD_LOGIC;
  SIGNAL mux_1668_nl : STD_LOGIC;
  SIGNAL mux_1667_nl : STD_LOGIC;
  SIGNAL mux_1703_nl : STD_LOGIC;
  SIGNAL mux_1664_nl : STD_LOGIC;
  SIGNAL mux_2121_nl : STD_LOGIC;
  SIGNAL mux_2120_nl : STD_LOGIC;
  SIGNAL mux_2119_nl : STD_LOGIC;
  SIGNAL mux_2118_nl : STD_LOGIC;
  SIGNAL mux_2117_nl : STD_LOGIC;
  SIGNAL or_2287_nl : STD_LOGIC;
  SIGNAL mux_2116_nl : STD_LOGIC;
  SIGNAL or_2286_nl : STD_LOGIC;
  SIGNAL or_2284_nl : STD_LOGIC;
  SIGNAL mux_2115_nl : STD_LOGIC;
  SIGNAL mux_2114_nl : STD_LOGIC;
  SIGNAL mux_2113_nl : STD_LOGIC;
  SIGNAL or_2283_nl : STD_LOGIC;
  SIGNAL mux_2112_nl : STD_LOGIC;
  SIGNAL mux_2111_nl : STD_LOGIC;
  SIGNAL mux_2109_nl : STD_LOGIC;
  SIGNAL or_2280_nl : STD_LOGIC;
  SIGNAL mux_2108_nl : STD_LOGIC;
  SIGNAL mux_2107_nl : STD_LOGIC;
  SIGNAL mux_2106_nl : STD_LOGIC;
  SIGNAL mux_2105_nl : STD_LOGIC;
  SIGNAL nand_390_nl : STD_LOGIC;
  SIGNAL mux_2100_nl : STD_LOGIC;
  SIGNAL mux_2099_nl : STD_LOGIC;
  SIGNAL mux_2096_nl : STD_LOGIC;
  SIGNAL or_2265_nl : STD_LOGIC;
  SIGNAL mux_2094_nl : STD_LOGIC;
  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL or_2258_nl : STD_LOGIC;
  SIGNAL mux_2153_nl : STD_LOGIC;
  SIGNAL mux_2152_nl : STD_LOGIC;
  SIGNAL mux_2151_nl : STD_LOGIC;
  SIGNAL mux_2150_nl : STD_LOGIC;
  SIGNAL mux_2149_nl : STD_LOGIC;
  SIGNAL or_2310_nl : STD_LOGIC;
  SIGNAL or_2309_nl : STD_LOGIC;
  SIGNAL mux_2148_nl : STD_LOGIC;
  SIGNAL mux_2147_nl : STD_LOGIC;
  SIGNAL mux_2146_nl : STD_LOGIC;
  SIGNAL or_2308_nl : STD_LOGIC;
  SIGNAL mux_2145_nl : STD_LOGIC;
  SIGNAL mux_2144_nl : STD_LOGIC;
  SIGNAL mux_2143_nl : STD_LOGIC;
  SIGNAL mux_2142_nl : STD_LOGIC;
  SIGNAL or_2305_nl : STD_LOGIC;
  SIGNAL mux_2141_nl : STD_LOGIC;
  SIGNAL nand_392_nl : STD_LOGIC;
  SIGNAL or_2304_nl : STD_LOGIC;
  SIGNAL mux_2140_nl : STD_LOGIC;
  SIGNAL mux_2139_nl : STD_LOGIC;
  SIGNAL mux_2138_nl : STD_LOGIC;
  SIGNAL mux_2137_nl : STD_LOGIC;
  SIGNAL mux_2136_nl : STD_LOGIC;
  SIGNAL or_2303_nl : STD_LOGIC;
  SIGNAL mux_2130_nl : STD_LOGIC;
  SIGNAL mux_2129_nl : STD_LOGIC;
  SIGNAL mux_2128_nl : STD_LOGIC;
  SIGNAL mux_2127_nl : STD_LOGIC;
  SIGNAL mux_2126_nl : STD_LOGIC;
  SIGNAL or_2367_nl : STD_LOGIC;
  SIGNAL or_2292_nl : STD_LOGIC;
  SIGNAL or_nl : STD_LOGIC;
  SIGNAL mux_1740_nl : STD_LOGIC;
  SIGNAL or_1923_nl : STD_LOGIC;
  SIGNAL or_1922_nl : STD_LOGIC;
  SIGNAL mux_2156_nl : STD_LOGIC;
  SIGNAL or_2365_nl : STD_LOGIC;
  SIGNAL mux_2155_nl : STD_LOGIC;
  SIGNAL or_2316_nl : STD_LOGIC;
  SIGNAL mux_2154_nl : STD_LOGIC;
  SIGNAL or_2315_nl : STD_LOGIC;
  SIGNAL or_2313_nl : STD_LOGIC;
  SIGNAL or_2366_nl : STD_LOGIC;
  SIGNAL mux_1749_nl : STD_LOGIC;
  SIGNAL nor_269_nl : STD_LOGIC;
  SIGNAL mux_1748_nl : STD_LOGIC;
  SIGNAL mux_1747_nl : STD_LOGIC;
  SIGNAL mux_1754_nl : STD_LOGIC;
  SIGNAL mux_1753_nl : STD_LOGIC;
  SIGNAL mux_1752_nl : STD_LOGIC;
  SIGNAL or_1936_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_1_acc_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL mux_1842_nl : STD_LOGIC;
  SIGNAL mux_1841_nl : STD_LOGIC;
  SIGNAL mux_1840_nl : STD_LOGIC;
  SIGNAL mux_1839_nl : STD_LOGIC;
  SIGNAL mux_1838_nl : STD_LOGIC;
  SIGNAL mux_1836_nl : STD_LOGIC;
  SIGNAL mux_1835_nl : STD_LOGIC;
  SIGNAL or_2033_nl : STD_LOGIC;
  SIGNAL nand_146_nl : STD_LOGIC;
  SIGNAL mux_1845_nl : STD_LOGIC;
  SIGNAL nand_338_nl : STD_LOGIC;
  SIGNAL mux_1848_nl : STD_LOGIC;
  SIGNAL mux_67_nl : STD_LOGIC;
  SIGNAL mux_66_nl : STD_LOGIC;
  SIGNAL or_23_nl : STD_LOGIC;
  SIGNAL nand_145_nl : STD_LOGIC;
  SIGNAL mux_1858_nl : STD_LOGIC;
  SIGNAL mux_1857_nl : STD_LOGIC;
  SIGNAL mux_1856_nl : STD_LOGIC;
  SIGNAL mux_1855_nl : STD_LOGIC;
  SIGNAL mux_1853_nl : STD_LOGIC;
  SIGNAL mux_1851_nl : STD_LOGIC;
  SIGNAL mux_1849_nl : STD_LOGIC;
  SIGNAL mux_1862_nl : STD_LOGIC;
  SIGNAL mux_1861_nl : STD_LOGIC;
  SIGNAL mux_1866_nl : STD_LOGIC;
  SIGNAL or_2041_nl : STD_LOGIC;
  SIGNAL mux_1865_nl : STD_LOGIC;
  SIGNAL mux_1864_nl : STD_LOGIC;
  SIGNAL mux_1863_nl : STD_LOGIC;
  SIGNAL mux_1869_nl : STD_LOGIC;
  SIGNAL mux_1868_nl : STD_LOGIC;
  SIGNAL mux_1867_nl : STD_LOGIC;
  SIGNAL or_2043_nl : STD_LOGIC;
  SIGNAL mux_1872_nl : STD_LOGIC;
  SIGNAL mux_1871_nl : STD_LOGIC;
  SIGNAL mux_1870_nl : STD_LOGIC;
  SIGNAL or_2175_nl : STD_LOGIC;
  SIGNAL mux_1874_nl : STD_LOGIC;
  SIGNAL mux_1873_nl : STD_LOGIC;
  SIGNAL and_248_nl : STD_LOGIC;
  SIGNAL mux_1875_nl : STD_LOGIC;
  SIGNAL and_213_nl : STD_LOGIC;
  SIGNAL mux_1877_nl : STD_LOGIC;
  SIGNAL or_2047_nl : STD_LOGIC;
  SIGNAL mux_1876_nl : STD_LOGIC;
  SIGNAL mux_1880_nl : STD_LOGIC;
  SIGNAL mux_1879_nl : STD_LOGIC;
  SIGNAL mux_1885_nl : STD_LOGIC;
  SIGNAL mux_1884_nl : STD_LOGIC;
  SIGNAL mux_1883_nl : STD_LOGIC;
  SIGNAL mux_1882_nl : STD_LOGIC;
  SIGNAL or_110_nl : STD_LOGIC;
  SIGNAL mux_1888_nl : STD_LOGIC;
  SIGNAL mux_1887_nl : STD_LOGIC;
  SIGNAL and_245_nl : STD_LOGIC;
  SIGNAL mux_459_nl : STD_LOGIC;
  SIGNAL mux_1896_nl : STD_LOGIC;
  SIGNAL mux_1895_nl : STD_LOGIC;
  SIGNAL mux_1894_nl : STD_LOGIC;
  SIGNAL mux_1893_nl : STD_LOGIC;
  SIGNAL mux_1892_nl : STD_LOGIC;
  SIGNAL mux_1891_nl : STD_LOGIC;
  SIGNAL nor_nl : STD_LOGIC;
  SIGNAL and_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_nor_11_nl : STD_LOGIC;
  SIGNAL mux_1904_nl : STD_LOGIC;
  SIGNAL nor_758_nl : STD_LOGIC;
  SIGNAL and_256_nl : STD_LOGIC;
  SIGNAL mux_1910_nl : STD_LOGIC;
  SIGNAL mux_1907_nl : STD_LOGIC;
  SIGNAL and_445_nl : STD_LOGIC;
  SIGNAL mux_1800_nl : STD_LOGIC;
  SIGNAL mux_1905_nl : STD_LOGIC;
  SIGNAL and_446_nl : STD_LOGIC;
  SIGNAL mux_1901_nl : STD_LOGIC;
  SIGNAL mux_1794_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_6_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_7_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_8_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_9_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_10_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_11_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_12_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_13_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_14_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_15_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_16_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_17_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_18_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_19_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_20_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_21_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_and_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_186_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL mux_1955_nl : STD_LOGIC;
  SIGNAL mux_1954_nl : STD_LOGIC;
  SIGNAL mux_1953_nl : STD_LOGIC;
  SIGNAL mux_1952_nl : STD_LOGIC;
  SIGNAL mux_1951_nl : STD_LOGIC;
  SIGNAL mux_1950_nl : STD_LOGIC;
  SIGNAL mux_1948_nl : STD_LOGIC;
  SIGNAL mux_1947_nl : STD_LOGIC;
  SIGNAL mux_1946_nl : STD_LOGIC;
  SIGNAL mux_1945_nl : STD_LOGIC;
  SIGNAL mux_1944_nl : STD_LOGIC;
  SIGNAL mux_1943_nl : STD_LOGIC;
  SIGNAL mux_1941_nl : STD_LOGIC;
  SIGNAL mux_1940_nl : STD_LOGIC;
  SIGNAL mux_1937_nl : STD_LOGIC;
  SIGNAL mux_1936_nl : STD_LOGIC;
  SIGNAL mux_1935_nl : STD_LOGIC;
  SIGNAL mux_1932_nl : STD_LOGIC;
  SIGNAL mux_1931_nl : STD_LOGIC;
  SIGNAL mux_1930_nl : STD_LOGIC;
  SIGNAL mux_1929_nl : STD_LOGIC;
  SIGNAL mux_1924_nl : STD_LOGIC;
  SIGNAL mux_1919_nl : STD_LOGIC;
  SIGNAL mux_1918_nl : STD_LOGIC;
  SIGNAL mux_1916_nl : STD_LOGIC;
  SIGNAL mux_1915_nl : STD_LOGIC;
  SIGNAL mux_1913_nl : STD_LOGIC;
  SIGNAL not_4628_nl : STD_LOGIC;
  SIGNAL not_nl : STD_LOGIC;
  SIGNAL mux_2196_nl : STD_LOGIC;
  SIGNAL mux_2195_nl : STD_LOGIC;
  SIGNAL mux_2194_nl : STD_LOGIC;
  SIGNAL mux_2193_nl : STD_LOGIC;
  SIGNAL mux_2192_nl : STD_LOGIC;
  SIGNAL mux_2191_nl : STD_LOGIC;
  SIGNAL mux_2190_nl : STD_LOGIC;
  SIGNAL mux_2189_nl : STD_LOGIC;
  SIGNAL mux_2187_nl : STD_LOGIC;
  SIGNAL mux_2186_nl : STD_LOGIC;
  SIGNAL mux_2185_nl : STD_LOGIC;
  SIGNAL mux_2184_nl : STD_LOGIC;
  SIGNAL mux_2183_nl : STD_LOGIC;
  SIGNAL mux_2182_nl : STD_LOGIC;
  SIGNAL mux_2181_nl : STD_LOGIC;
  SIGNAL mux_2177_nl : STD_LOGIC;
  SIGNAL mux_2174_nl : STD_LOGIC;
  SIGNAL mux_2173_nl : STD_LOGIC;
  SIGNAL mux_2172_nl : STD_LOGIC;
  SIGNAL mux_2165_nl : STD_LOGIC;
  SIGNAL mux_2161_nl : STD_LOGIC;
  SIGNAL mux_2157_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_k_COMP_LOOP_k_mux_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL mux_2243_nl : STD_LOGIC;
  SIGNAL mux_2242_nl : STD_LOGIC;
  SIGNAL mux_2241_nl : STD_LOGIC;
  SIGNAL mux_2240_nl : STD_LOGIC;
  SIGNAL mux_2239_nl : STD_LOGIC;
  SIGNAL mux_2238_nl : STD_LOGIC;
  SIGNAL mux_2237_nl : STD_LOGIC;
  SIGNAL or_2347_nl : STD_LOGIC;
  SIGNAL mux_2236_nl : STD_LOGIC;
  SIGNAL mux_2235_nl : STD_LOGIC;
  SIGNAL mux_2234_nl : STD_LOGIC;
  SIGNAL mux_2233_nl : STD_LOGIC;
  SIGNAL mux_2230_nl : STD_LOGIC;
  SIGNAL mux_2228_nl : STD_LOGIC;
  SIGNAL mux_2227_nl : STD_LOGIC;
  SIGNAL mux_2226_nl : STD_LOGIC;
  SIGNAL mux_2225_nl : STD_LOGIC;
  SIGNAL mux_2224_nl : STD_LOGIC;
  SIGNAL mux_2223_nl : STD_LOGIC;
  SIGNAL mux_2218_nl : STD_LOGIC;
  SIGNAL mux_2213_nl : STD_LOGIC;
  SIGNAL mux_2212_nl : STD_LOGIC;
  SIGNAL mux_2210_nl : STD_LOGIC;
  SIGNAL mux_2209_nl : STD_LOGIC;
  SIGNAL mux_2207_nl : STD_LOGIC;
  SIGNAL mux_2204_nl : STD_LOGIC;
  SIGNAL mux_2203_nl : STD_LOGIC;
  SIGNAL mux_2201_nl : STD_LOGIC;
  SIGNAL mux_2200_nl : STD_LOGIC;
  SIGNAL mux_2198_nl : STD_LOGIC;
  SIGNAL mux_2262_nl : STD_LOGIC;
  SIGNAL nor_797_nl : STD_LOGIC;
  SIGNAL mux_2261_nl : STD_LOGIC;
  SIGNAL mux_2260_nl : STD_LOGIC;
  SIGNAL nand_396_nl : STD_LOGIC;
  SIGNAL mux_2259_nl : STD_LOGIC;
  SIGNAL or_2362_nl : STD_LOGIC;
  SIGNAL mux_2258_nl : STD_LOGIC;
  SIGNAL mux_2257_nl : STD_LOGIC;
  SIGNAL nand_397_nl : STD_LOGIC;
  SIGNAL mux_2255_nl : STD_LOGIC;
  SIGNAL and_700_nl : STD_LOGIC;
  SIGNAL mux_2254_nl : STD_LOGIC;
  SIGNAL nor_798_nl : STD_LOGIC;
  SIGNAL mux_2253_nl : STD_LOGIC;
  SIGNAL nor_799_nl : STD_LOGIC;
  SIGNAL nor_800_nl : STD_LOGIC;
  SIGNAL mux_2252_nl : STD_LOGIC;
  SIGNAL or_2356_nl : STD_LOGIC;
  SIGNAL mux_2250_nl : STD_LOGIC;
  SIGNAL nand_394_nl : STD_LOGIC;
  SIGNAL mux_2247_nl : STD_LOGIC;
  SIGNAL nand_398_nl : STD_LOGIC;
  SIGNAL mux_2246_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_209_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_and_930_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_932_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_934_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_and_936_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_27_nl : STD_LOGIC;
  SIGNAL mux_51_nl : STD_LOGIC;
  SIGNAL nor_727_nl : STD_LOGIC;
  SIGNAL or_2152_nl : STD_LOGIC;
  SIGNAL nand_314_nl : STD_LOGIC;
  SIGNAL mux_514_nl : STD_LOGIC;
  SIGNAL or_265_nl : STD_LOGIC;
  SIGNAL mux_520_nl : STD_LOGIC;
  SIGNAL mux_1520_nl : STD_LOGIC;
  SIGNAL mux_1548_nl : STD_LOGIC;
  SIGNAL mux_1564_nl : STD_LOGIC;
  SIGNAL mux_1584_nl : STD_LOGIC;
  SIGNAL mux_1587_nl : STD_LOGIC;
  SIGNAL mux_1601_nl : STD_LOGIC;
  SIGNAL nor_275_nl : STD_LOGIC;
  SIGNAL mux_1611_nl : STD_LOGIC;
  SIGNAL and_272_nl : STD_LOGIC;
  SIGNAL mux_1610_nl : STD_LOGIC;
  SIGNAL nor_272_nl : STD_LOGIC;
  SIGNAL mux_1606_nl : STD_LOGIC;
  SIGNAL mux_1605_nl : STD_LOGIC;
  SIGNAL nor_273_nl : STD_LOGIC;
  SIGNAL and_273_nl : STD_LOGIC;
  SIGNAL mux_1603_nl : STD_LOGIC;
  SIGNAL nor_274_nl : STD_LOGIC;
  SIGNAL or_1849_nl : STD_LOGIC;
  SIGNAL or_1863_nl : STD_LOGIC;
  SIGNAL mux_1671_nl : STD_LOGIC;
  SIGNAL nand_111_nl : STD_LOGIC;
  SIGNAL mux_1670_nl : STD_LOGIC;
  SIGNAL nand_110_nl : STD_LOGIC;
  SIGNAL mux_1679_nl : STD_LOGIC;
  SIGNAL nand_151_nl : STD_LOGIC;
  SIGNAL nand_342_nl : STD_LOGIC;
  SIGNAL or_2000_nl : STD_LOGIC;
  SIGNAL mux_1779_nl : STD_LOGIC;
  SIGNAL and_261_nl : STD_LOGIC;
  SIGNAL mux_1804_nl : STD_LOGIC;
  SIGNAL mux_1803_nl : STD_LOGIC;
  SIGNAL or_1996_nl : STD_LOGIC;
  SIGNAL mux_1774_nl : STD_LOGIC;
  SIGNAL mux_1770_nl : STD_LOGIC;
  SIGNAL and_263_nl : STD_LOGIC;
  SIGNAL mux_1769_nl : STD_LOGIC;
  SIGNAL mux_1831_nl : STD_LOGIC;
  SIGNAL mux_1830_nl : STD_LOGIC;
  SIGNAL mux_1829_nl : STD_LOGIC;
  SIGNAL mux_1828_nl : STD_LOGIC;
  SIGNAL mux_1827_nl : STD_LOGIC;
  SIGNAL nor_248_nl : STD_LOGIC;
  SIGNAL mux_1843_nl : STD_LOGIC;
  SIGNAL nor_244_nl : STD_LOGIC;
  SIGNAL and_368_nl : STD_LOGIC;
  SIGNAL or_2091_nl : STD_LOGIC;
  SIGNAL and_42_nl : STD_LOGIC;
  SIGNAL and_52_nl : STD_LOGIC;
  SIGNAL and_57_nl : STD_LOGIC;
  SIGNAL and_67_nl : STD_LOGIC;
  SIGNAL and_73_nl : STD_LOGIC;
  SIGNAL and_80_nl : STD_LOGIC;
  SIGNAL and_87_nl : STD_LOGIC;
  SIGNAL and_93_nl : STD_LOGIC;
  SIGNAL and_99_nl : STD_LOGIC;
  SIGNAL and_103_nl : STD_LOGIC;
  SIGNAL and_107_nl : STD_LOGIC;
  SIGNAL and_111_nl : STD_LOGIC;
  SIGNAL and_116_nl : STD_LOGIC;
  SIGNAL and_120_nl : STD_LOGIC;
  SIGNAL and_124_nl : STD_LOGIC;
  SIGNAL and_129_nl : STD_LOGIC;
  SIGNAL and_131_nl : STD_LOGIC;
  SIGNAL mux_526_nl : STD_LOGIC;
  SIGNAL mux_525_nl : STD_LOGIC;
  SIGNAL or_280_nl : STD_LOGIC;
  SIGNAL mux_524_nl : STD_LOGIC;
  SIGNAL mux_523_nl : STD_LOGIC;
  SIGNAL mux_522_nl : STD_LOGIC;
  SIGNAL mux_521_nl : STD_LOGIC;
  SIGNAL or_275_nl : STD_LOGIC;
  SIGNAL mux_519_nl : STD_LOGIC;
  SIGNAL or_274_nl : STD_LOGIC;
  SIGNAL mux_518_nl : STD_LOGIC;
  SIGNAL mux_517_nl : STD_LOGIC;
  SIGNAL or_272_nl : STD_LOGIC;
  SIGNAL mux_516_nl : STD_LOGIC;
  SIGNAL or_271_nl : STD_LOGIC;
  SIGNAL or_269_nl : STD_LOGIC;
  SIGNAL mux_515_nl : STD_LOGIC;
  SIGNAL and_132_nl : STD_LOGIC;
  SIGNAL and_134_nl : STD_LOGIC;
  SIGNAL and_135_nl : STD_LOGIC;
  SIGNAL and_136_nl : STD_LOGIC;
  SIGNAL and_137_nl : STD_LOGIC;
  SIGNAL and_138_nl : STD_LOGIC;
  SIGNAL and_139_nl : STD_LOGIC;
  SIGNAL and_140_nl : STD_LOGIC;
  SIGNAL and_142_nl : STD_LOGIC;
  SIGNAL and_144_nl : STD_LOGIC;
  SIGNAL and_145_nl : STD_LOGIC;
  SIGNAL and_146_nl : STD_LOGIC;
  SIGNAL and_148_nl : STD_LOGIC;
  SIGNAL and_150_nl : STD_LOGIC;
  SIGNAL and_152_nl : STD_LOGIC;
  SIGNAL mux_556_nl : STD_LOGIC;
  SIGNAL mux_555_nl : STD_LOGIC;
  SIGNAL nor_689_nl : STD_LOGIC;
  SIGNAL mux_554_nl : STD_LOGIC;
  SIGNAL nand_10_nl : STD_LOGIC;
  SIGNAL mux_553_nl : STD_LOGIC;
  SIGNAL mux_552_nl : STD_LOGIC;
  SIGNAL or_319_nl : STD_LOGIC;
  SIGNAL mux_551_nl : STD_LOGIC;
  SIGNAL or_318_nl : STD_LOGIC;
  SIGNAL or_317_nl : STD_LOGIC;
  SIGNAL mux_550_nl : STD_LOGIC;
  SIGNAL nor_690_nl : STD_LOGIC;
  SIGNAL nor_691_nl : STD_LOGIC;
  SIGNAL mux_549_nl : STD_LOGIC;
  SIGNAL or_313_nl : STD_LOGIC;
  SIGNAL mux_548_nl : STD_LOGIC;
  SIGNAL and_344_nl : STD_LOGIC;
  SIGNAL mux_547_nl : STD_LOGIC;
  SIGNAL or_310_nl : STD_LOGIC;
  SIGNAL mux_546_nl : STD_LOGIC;
  SIGNAL mux_545_nl : STD_LOGIC;
  SIGNAL mux_544_nl : STD_LOGIC;
  SIGNAL or_308_nl : STD_LOGIC;
  SIGNAL mux_543_nl : STD_LOGIC;
  SIGNAL or_306_nl : STD_LOGIC;
  SIGNAL or_305_nl : STD_LOGIC;
  SIGNAL mux_542_nl : STD_LOGIC;
  SIGNAL or_304_nl : STD_LOGIC;
  SIGNAL nor_692_nl : STD_LOGIC;
  SIGNAL mux_541_nl : STD_LOGIC;
  SIGNAL nor_693_nl : STD_LOGIC;
  SIGNAL mux_540_nl : STD_LOGIC;
  SIGNAL mux_539_nl : STD_LOGIC;
  SIGNAL or_301_nl : STD_LOGIC;
  SIGNAL mux_538_nl : STD_LOGIC;
  SIGNAL mux_537_nl : STD_LOGIC;
  SIGNAL or_299_nl : STD_LOGIC;
  SIGNAL mux_536_nl : STD_LOGIC;
  SIGNAL or_297_nl : STD_LOGIC;
  SIGNAL mux_535_nl : STD_LOGIC;
  SIGNAL or_296_nl : STD_LOGIC;
  SIGNAL mux_534_nl : STD_LOGIC;
  SIGNAL or_295_nl : STD_LOGIC;
  SIGNAL nor_694_nl : STD_LOGIC;
  SIGNAL mux_533_nl : STD_LOGIC;
  SIGNAL nand_8_nl : STD_LOGIC;
  SIGNAL mux_532_nl : STD_LOGIC;
  SIGNAL or_292_nl : STD_LOGIC;
  SIGNAL mux_531_nl : STD_LOGIC;
  SIGNAL mux_530_nl : STD_LOGIC;
  SIGNAL or_290_nl : STD_LOGIC;
  SIGNAL mux_529_nl : STD_LOGIC;
  SIGNAL or_286_nl : STD_LOGIC;
  SIGNAL or_285_nl : STD_LOGIC;
  SIGNAL mux_528_nl : STD_LOGIC;
  SIGNAL or_284_nl : STD_LOGIC;
  SIGNAL mux_527_nl : STD_LOGIC;
  SIGNAL or_283_nl : STD_LOGIC;
  SIGNAL mux_587_nl : STD_LOGIC;
  SIGNAL mux_586_nl : STD_LOGIC;
  SIGNAL nor_669_nl : STD_LOGIC;
  SIGNAL mux_585_nl : STD_LOGIC;
  SIGNAL mux_584_nl : STD_LOGIC;
  SIGNAL or_372_nl : STD_LOGIC;
  SIGNAL mux_583_nl : STD_LOGIC;
  SIGNAL or_371_nl : STD_LOGIC;
  SIGNAL mux_582_nl : STD_LOGIC;
  SIGNAL mux_581_nl : STD_LOGIC;
  SIGNAL or_366_nl : STD_LOGIC;
  SIGNAL mux_580_nl : STD_LOGIC;
  SIGNAL or_365_nl : STD_LOGIC;
  SIGNAL or_363_nl : STD_LOGIC;
  SIGNAL mux_579_nl : STD_LOGIC;
  SIGNAL nor_670_nl : STD_LOGIC;
  SIGNAL mux_578_nl : STD_LOGIC;
  SIGNAL mux_577_nl : STD_LOGIC;
  SIGNAL or_361_nl : STD_LOGIC;
  SIGNAL or_359_nl : STD_LOGIC;
  SIGNAL or_358_nl : STD_LOGIC;
  SIGNAL nor_671_nl : STD_LOGIC;
  SIGNAL mux_576_nl : STD_LOGIC;
  SIGNAL mux_575_nl : STD_LOGIC;
  SIGNAL nor_672_nl : STD_LOGIC;
  SIGNAL and_342_nl : STD_LOGIC;
  SIGNAL mux_574_nl : STD_LOGIC;
  SIGNAL nor_673_nl : STD_LOGIC;
  SIGNAL mux_573_nl : STD_LOGIC;
  SIGNAL nor_674_nl : STD_LOGIC;
  SIGNAL nor_675_nl : STD_LOGIC;
  SIGNAL and_343_nl : STD_LOGIC;
  SIGNAL mux_572_nl : STD_LOGIC;
  SIGNAL mux_571_nl : STD_LOGIC;
  SIGNAL mux_570_nl : STD_LOGIC;
  SIGNAL nor_676_nl : STD_LOGIC;
  SIGNAL nor_677_nl : STD_LOGIC;
  SIGNAL mux_569_nl : STD_LOGIC;
  SIGNAL nor_679_nl : STD_LOGIC;
  SIGNAL mux_568_nl : STD_LOGIC;
  SIGNAL mux_567_nl : STD_LOGIC;
  SIGNAL nor_680_nl : STD_LOGIC;
  SIGNAL nor_681_nl : STD_LOGIC;
  SIGNAL nor_682_nl : STD_LOGIC;
  SIGNAL nor_683_nl : STD_LOGIC;
  SIGNAL mux_566_nl : STD_LOGIC;
  SIGNAL nand_11_nl : STD_LOGIC;
  SIGNAL mux_565_nl : STD_LOGIC;
  SIGNAL mux_564_nl : STD_LOGIC;
  SIGNAL mux_563_nl : STD_LOGIC;
  SIGNAL nor_685_nl : STD_LOGIC;
  SIGNAL mux_562_nl : STD_LOGIC;
  SIGNAL nor_686_nl : STD_LOGIC;
  SIGNAL nor_687_nl : STD_LOGIC;
  SIGNAL nor_688_nl : STD_LOGIC;
  SIGNAL or_329_nl : STD_LOGIC;
  SIGNAL mux_561_nl : STD_LOGIC;
  SIGNAL or_328_nl : STD_LOGIC;
  SIGNAL mux_560_nl : STD_LOGIC;
  SIGNAL mux_559_nl : STD_LOGIC;
  SIGNAL or_326_nl : STD_LOGIC;
  SIGNAL mux_558_nl : STD_LOGIC;
  SIGNAL or_322_nl : STD_LOGIC;
  SIGNAL mux_618_nl : STD_LOGIC;
  SIGNAL mux_617_nl : STD_LOGIC;
  SIGNAL mux_616_nl : STD_LOGIC;
  SIGNAL nor_661_nl : STD_LOGIC;
  SIGNAL mux_615_nl : STD_LOGIC;
  SIGNAL mux_614_nl : STD_LOGIC;
  SIGNAL or_413_nl : STD_LOGIC;
  SIGNAL mux_613_nl : STD_LOGIC;
  SIGNAL or_412_nl : STD_LOGIC;
  SIGNAL and_341_nl : STD_LOGIC;
  SIGNAL mux_612_nl : STD_LOGIC;
  SIGNAL or_410_nl : STD_LOGIC;
  SIGNAL mux_611_nl : STD_LOGIC;
  SIGNAL mux_610_nl : STD_LOGIC;
  SIGNAL or_409_nl : STD_LOGIC;
  SIGNAL mux_609_nl : STD_LOGIC;
  SIGNAL or_408_nl : STD_LOGIC;
  SIGNAL nor_662_nl : STD_LOGIC;
  SIGNAL mux_608_nl : STD_LOGIC;
  SIGNAL or_405_nl : STD_LOGIC;
  SIGNAL nor_663_nl : STD_LOGIC;
  SIGNAL mux_607_nl : STD_LOGIC;
  SIGNAL mux_606_nl : STD_LOGIC;
  SIGNAL or_402_nl : STD_LOGIC;
  SIGNAL or_401_nl : STD_LOGIC;
  SIGNAL nand_14_nl : STD_LOGIC;
  SIGNAL mux_605_nl : STD_LOGIC;
  SIGNAL or_400_nl : STD_LOGIC;
  SIGNAL mux_604_nl : STD_LOGIC;
  SIGNAL or_399_nl : STD_LOGIC;
  SIGNAL mux_603_nl : STD_LOGIC;
  SIGNAL mux_602_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL mux_601_nl : STD_LOGIC;
  SIGNAL nor_665_nl : STD_LOGIC;
  SIGNAL nor_666_nl : STD_LOGIC;
  SIGNAL mux_600_nl : STD_LOGIC;
  SIGNAL or_394_nl : STD_LOGIC;
  SIGNAL mux_599_nl : STD_LOGIC;
  SIGNAL or_393_nl : STD_LOGIC;
  SIGNAL mux_598_nl : STD_LOGIC;
  SIGNAL nor_667_nl : STD_LOGIC;
  SIGNAL mux_597_nl : STD_LOGIC;
  SIGNAL or_389_nl : STD_LOGIC;
  SIGNAL mux_596_nl : STD_LOGIC;
  SIGNAL mux_595_nl : STD_LOGIC;
  SIGNAL or_388_nl : STD_LOGIC;
  SIGNAL mux_594_nl : STD_LOGIC;
  SIGNAL or_387_nl : STD_LOGIC;
  SIGNAL nor_668_nl : STD_LOGIC;
  SIGNAL mux_593_nl : STD_LOGIC;
  SIGNAL mux_592_nl : STD_LOGIC;
  SIGNAL mux_591_nl : STD_LOGIC;
  SIGNAL or_383_nl : STD_LOGIC;
  SIGNAL mux_590_nl : STD_LOGIC;
  SIGNAL or_380_nl : STD_LOGIC;
  SIGNAL or_378_nl : STD_LOGIC;
  SIGNAL mux_589_nl : STD_LOGIC;
  SIGNAL or_377_nl : STD_LOGIC;
  SIGNAL mux_649_nl : STD_LOGIC;
  SIGNAL mux_648_nl : STD_LOGIC;
  SIGNAL nor_641_nl : STD_LOGIC;
  SIGNAL mux_647_nl : STD_LOGIC;
  SIGNAL mux_646_nl : STD_LOGIC;
  SIGNAL or_465_nl : STD_LOGIC;
  SIGNAL mux_645_nl : STD_LOGIC;
  SIGNAL or_464_nl : STD_LOGIC;
  SIGNAL mux_644_nl : STD_LOGIC;
  SIGNAL mux_643_nl : STD_LOGIC;
  SIGNAL or_461_nl : STD_LOGIC;
  SIGNAL or_459_nl : STD_LOGIC;
  SIGNAL mux_642_nl : STD_LOGIC;
  SIGNAL or_458_nl : STD_LOGIC;
  SIGNAL or_456_nl : STD_LOGIC;
  SIGNAL mux_641_nl : STD_LOGIC;
  SIGNAL nor_642_nl : STD_LOGIC;
  SIGNAL mux_640_nl : STD_LOGIC;
  SIGNAL mux_639_nl : STD_LOGIC;
  SIGNAL or_454_nl : STD_LOGIC;
  SIGNAL or_452_nl : STD_LOGIC;
  SIGNAL or_451_nl : STD_LOGIC;
  SIGNAL nor_643_nl : STD_LOGIC;
  SIGNAL mux_638_nl : STD_LOGIC;
  SIGNAL mux_637_nl : STD_LOGIC;
  SIGNAL nor_644_nl : STD_LOGIC;
  SIGNAL and_339_nl : STD_LOGIC;
  SIGNAL mux_636_nl : STD_LOGIC;
  SIGNAL nor_645_nl : STD_LOGIC;
  SIGNAL mux_635_nl : STD_LOGIC;
  SIGNAL nor_646_nl : STD_LOGIC;
  SIGNAL nor_647_nl : STD_LOGIC;
  SIGNAL and_340_nl : STD_LOGIC;
  SIGNAL mux_634_nl : STD_LOGIC;
  SIGNAL mux_633_nl : STD_LOGIC;
  SIGNAL mux_632_nl : STD_LOGIC;
  SIGNAL nor_648_nl : STD_LOGIC;
  SIGNAL nor_649_nl : STD_LOGIC;
  SIGNAL mux_631_nl : STD_LOGIC;
  SIGNAL nor_651_nl : STD_LOGIC;
  SIGNAL mux_630_nl : STD_LOGIC;
  SIGNAL mux_629_nl : STD_LOGIC;
  SIGNAL nor_652_nl : STD_LOGIC;
  SIGNAL nor_653_nl : STD_LOGIC;
  SIGNAL nor_654_nl : STD_LOGIC;
  SIGNAL nor_655_nl : STD_LOGIC;
  SIGNAL mux_628_nl : STD_LOGIC;
  SIGNAL nand_17_nl : STD_LOGIC;
  SIGNAL mux_627_nl : STD_LOGIC;
  SIGNAL mux_626_nl : STD_LOGIC;
  SIGNAL mux_625_nl : STD_LOGIC;
  SIGNAL nor_657_nl : STD_LOGIC;
  SIGNAL mux_624_nl : STD_LOGIC;
  SIGNAL nor_658_nl : STD_LOGIC;
  SIGNAL nor_659_nl : STD_LOGIC;
  SIGNAL nor_660_nl : STD_LOGIC;
  SIGNAL or_422_nl : STD_LOGIC;
  SIGNAL mux_623_nl : STD_LOGIC;
  SIGNAL or_421_nl : STD_LOGIC;
  SIGNAL mux_622_nl : STD_LOGIC;
  SIGNAL mux_621_nl : STD_LOGIC;
  SIGNAL or_419_nl : STD_LOGIC;
  SIGNAL or_418_nl : STD_LOGIC;
  SIGNAL mux_620_nl : STD_LOGIC;
  SIGNAL or_415_nl : STD_LOGIC;
  SIGNAL mux_680_nl : STD_LOGIC;
  SIGNAL mux_679_nl : STD_LOGIC;
  SIGNAL nor_635_nl : STD_LOGIC;
  SIGNAL mux_678_nl : STD_LOGIC;
  SIGNAL nand_22_nl : STD_LOGIC;
  SIGNAL mux_677_nl : STD_LOGIC;
  SIGNAL mux_676_nl : STD_LOGIC;
  SIGNAL or_505_nl : STD_LOGIC;
  SIGNAL mux_675_nl : STD_LOGIC;
  SIGNAL or_504_nl : STD_LOGIC;
  SIGNAL or_503_nl : STD_LOGIC;
  SIGNAL mux_674_nl : STD_LOGIC;
  SIGNAL nor_636_nl : STD_LOGIC;
  SIGNAL nor_637_nl : STD_LOGIC;
  SIGNAL mux_673_nl : STD_LOGIC;
  SIGNAL or_499_nl : STD_LOGIC;
  SIGNAL mux_672_nl : STD_LOGIC;
  SIGNAL and_338_nl : STD_LOGIC;
  SIGNAL mux_671_nl : STD_LOGIC;
  SIGNAL or_496_nl : STD_LOGIC;
  SIGNAL mux_670_nl : STD_LOGIC;
  SIGNAL mux_669_nl : STD_LOGIC;
  SIGNAL mux_668_nl : STD_LOGIC;
  SIGNAL or_494_nl : STD_LOGIC;
  SIGNAL mux_667_nl : STD_LOGIC;
  SIGNAL or_492_nl : STD_LOGIC;
  SIGNAL or_491_nl : STD_LOGIC;
  SIGNAL mux_666_nl : STD_LOGIC;
  SIGNAL or_490_nl : STD_LOGIC;
  SIGNAL nor_638_nl : STD_LOGIC;
  SIGNAL mux_665_nl : STD_LOGIC;
  SIGNAL nor_639_nl : STD_LOGIC;
  SIGNAL mux_664_nl : STD_LOGIC;
  SIGNAL mux_663_nl : STD_LOGIC;
  SIGNAL or_487_nl : STD_LOGIC;
  SIGNAL mux_662_nl : STD_LOGIC;
  SIGNAL mux_661_nl : STD_LOGIC;
  SIGNAL or_485_nl : STD_LOGIC;
  SIGNAL mux_660_nl : STD_LOGIC;
  SIGNAL or_483_nl : STD_LOGIC;
  SIGNAL mux_659_nl : STD_LOGIC;
  SIGNAL or_482_nl : STD_LOGIC;
  SIGNAL mux_658_nl : STD_LOGIC;
  SIGNAL or_481_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL mux_657_nl : STD_LOGIC;
  SIGNAL nand_20_nl : STD_LOGIC;
  SIGNAL mux_656_nl : STD_LOGIC;
  SIGNAL or_478_nl : STD_LOGIC;
  SIGNAL mux_655_nl : STD_LOGIC;
  SIGNAL mux_654_nl : STD_LOGIC;
  SIGNAL or_476_nl : STD_LOGIC;
  SIGNAL mux_653_nl : STD_LOGIC;
  SIGNAL or_472_nl : STD_LOGIC;
  SIGNAL or_471_nl : STD_LOGIC;
  SIGNAL mux_652_nl : STD_LOGIC;
  SIGNAL or_470_nl : STD_LOGIC;
  SIGNAL mux_651_nl : STD_LOGIC;
  SIGNAL or_469_nl : STD_LOGIC;
  SIGNAL mux_711_nl : STD_LOGIC;
  SIGNAL mux_710_nl : STD_LOGIC;
  SIGNAL nor_615_nl : STD_LOGIC;
  SIGNAL mux_709_nl : STD_LOGIC;
  SIGNAL mux_708_nl : STD_LOGIC;
  SIGNAL or_558_nl : STD_LOGIC;
  SIGNAL mux_707_nl : STD_LOGIC;
  SIGNAL or_557_nl : STD_LOGIC;
  SIGNAL mux_706_nl : STD_LOGIC;
  SIGNAL mux_705_nl : STD_LOGIC;
  SIGNAL or_552_nl : STD_LOGIC;
  SIGNAL mux_704_nl : STD_LOGIC;
  SIGNAL or_551_nl : STD_LOGIC;
  SIGNAL or_549_nl : STD_LOGIC;
  SIGNAL mux_703_nl : STD_LOGIC;
  SIGNAL nor_616_nl : STD_LOGIC;
  SIGNAL mux_702_nl : STD_LOGIC;
  SIGNAL mux_701_nl : STD_LOGIC;
  SIGNAL or_547_nl : STD_LOGIC;
  SIGNAL or_545_nl : STD_LOGIC;
  SIGNAL or_544_nl : STD_LOGIC;
  SIGNAL nor_617_nl : STD_LOGIC;
  SIGNAL mux_700_nl : STD_LOGIC;
  SIGNAL mux_699_nl : STD_LOGIC;
  SIGNAL nor_618_nl : STD_LOGIC;
  SIGNAL and_336_nl : STD_LOGIC;
  SIGNAL mux_698_nl : STD_LOGIC;
  SIGNAL nor_619_nl : STD_LOGIC;
  SIGNAL mux_697_nl : STD_LOGIC;
  SIGNAL nor_620_nl : STD_LOGIC;
  SIGNAL nor_621_nl : STD_LOGIC;
  SIGNAL and_337_nl : STD_LOGIC;
  SIGNAL mux_696_nl : STD_LOGIC;
  SIGNAL mux_695_nl : STD_LOGIC;
  SIGNAL mux_694_nl : STD_LOGIC;
  SIGNAL nor_622_nl : STD_LOGIC;
  SIGNAL nor_623_nl : STD_LOGIC;
  SIGNAL mux_693_nl : STD_LOGIC;
  SIGNAL nor_625_nl : STD_LOGIC;
  SIGNAL mux_692_nl : STD_LOGIC;
  SIGNAL mux_691_nl : STD_LOGIC;
  SIGNAL nor_626_nl : STD_LOGIC;
  SIGNAL nor_627_nl : STD_LOGIC;
  SIGNAL nor_628_nl : STD_LOGIC;
  SIGNAL nor_629_nl : STD_LOGIC;
  SIGNAL mux_690_nl : STD_LOGIC;
  SIGNAL nand_23_nl : STD_LOGIC;
  SIGNAL mux_689_nl : STD_LOGIC;
  SIGNAL mux_688_nl : STD_LOGIC;
  SIGNAL mux_687_nl : STD_LOGIC;
  SIGNAL nor_631_nl : STD_LOGIC;
  SIGNAL mux_686_nl : STD_LOGIC;
  SIGNAL nor_632_nl : STD_LOGIC;
  SIGNAL nor_633_nl : STD_LOGIC;
  SIGNAL nor_634_nl : STD_LOGIC;
  SIGNAL or_515_nl : STD_LOGIC;
  SIGNAL mux_685_nl : STD_LOGIC;
  SIGNAL or_514_nl : STD_LOGIC;
  SIGNAL mux_684_nl : STD_LOGIC;
  SIGNAL mux_683_nl : STD_LOGIC;
  SIGNAL or_512_nl : STD_LOGIC;
  SIGNAL mux_682_nl : STD_LOGIC;
  SIGNAL or_508_nl : STD_LOGIC;
  SIGNAL mux_742_nl : STD_LOGIC;
  SIGNAL mux_741_nl : STD_LOGIC;
  SIGNAL nor_609_nl : STD_LOGIC;
  SIGNAL mux_740_nl : STD_LOGIC;
  SIGNAL nand_28_nl : STD_LOGIC;
  SIGNAL mux_739_nl : STD_LOGIC;
  SIGNAL mux_738_nl : STD_LOGIC;
  SIGNAL or_598_nl : STD_LOGIC;
  SIGNAL mux_737_nl : STD_LOGIC;
  SIGNAL or_597_nl : STD_LOGIC;
  SIGNAL or_596_nl : STD_LOGIC;
  SIGNAL mux_736_nl : STD_LOGIC;
  SIGNAL and_439_nl : STD_LOGIC;
  SIGNAL nor_611_nl : STD_LOGIC;
  SIGNAL mux_735_nl : STD_LOGIC;
  SIGNAL or_592_nl : STD_LOGIC;
  SIGNAL mux_734_nl : STD_LOGIC;
  SIGNAL and_335_nl : STD_LOGIC;
  SIGNAL mux_733_nl : STD_LOGIC;
  SIGNAL or_589_nl : STD_LOGIC;
  SIGNAL mux_732_nl : STD_LOGIC;
  SIGNAL mux_731_nl : STD_LOGIC;
  SIGNAL mux_730_nl : STD_LOGIC;
  SIGNAL or_587_nl : STD_LOGIC;
  SIGNAL mux_729_nl : STD_LOGIC;
  SIGNAL or_585_nl : STD_LOGIC;
  SIGNAL or_584_nl : STD_LOGIC;
  SIGNAL mux_728_nl : STD_LOGIC;
  SIGNAL or_583_nl : STD_LOGIC;
  SIGNAL nor_612_nl : STD_LOGIC;
  SIGNAL mux_727_nl : STD_LOGIC;
  SIGNAL nor_613_nl : STD_LOGIC;
  SIGNAL mux_726_nl : STD_LOGIC;
  SIGNAL mux_725_nl : STD_LOGIC;
  SIGNAL or_580_nl : STD_LOGIC;
  SIGNAL mux_724_nl : STD_LOGIC;
  SIGNAL mux_723_nl : STD_LOGIC;
  SIGNAL or_578_nl : STD_LOGIC;
  SIGNAL mux_722_nl : STD_LOGIC;
  SIGNAL or_576_nl : STD_LOGIC;
  SIGNAL mux_721_nl : STD_LOGIC;
  SIGNAL or_575_nl : STD_LOGIC;
  SIGNAL mux_720_nl : STD_LOGIC;
  SIGNAL or_574_nl : STD_LOGIC;
  SIGNAL nor_614_nl : STD_LOGIC;
  SIGNAL mux_719_nl : STD_LOGIC;
  SIGNAL nand_26_nl : STD_LOGIC;
  SIGNAL mux_718_nl : STD_LOGIC;
  SIGNAL or_571_nl : STD_LOGIC;
  SIGNAL mux_717_nl : STD_LOGIC;
  SIGNAL mux_716_nl : STD_LOGIC;
  SIGNAL or_569_nl : STD_LOGIC;
  SIGNAL mux_715_nl : STD_LOGIC;
  SIGNAL or_565_nl : STD_LOGIC;
  SIGNAL or_564_nl : STD_LOGIC;
  SIGNAL mux_714_nl : STD_LOGIC;
  SIGNAL or_563_nl : STD_LOGIC;
  SIGNAL mux_713_nl : STD_LOGIC;
  SIGNAL or_562_nl : STD_LOGIC;
  SIGNAL mux_773_nl : STD_LOGIC;
  SIGNAL mux_772_nl : STD_LOGIC;
  SIGNAL nor_589_nl : STD_LOGIC;
  SIGNAL mux_771_nl : STD_LOGIC;
  SIGNAL mux_770_nl : STD_LOGIC;
  SIGNAL or_651_nl : STD_LOGIC;
  SIGNAL mux_769_nl : STD_LOGIC;
  SIGNAL or_650_nl : STD_LOGIC;
  SIGNAL mux_768_nl : STD_LOGIC;
  SIGNAL mux_767_nl : STD_LOGIC;
  SIGNAL or_647_nl : STD_LOGIC;
  SIGNAL or_645_nl : STD_LOGIC;
  SIGNAL mux_766_nl : STD_LOGIC;
  SIGNAL or_644_nl : STD_LOGIC;
  SIGNAL or_642_nl : STD_LOGIC;
  SIGNAL mux_765_nl : STD_LOGIC;
  SIGNAL nor_590_nl : STD_LOGIC;
  SIGNAL mux_764_nl : STD_LOGIC;
  SIGNAL mux_763_nl : STD_LOGIC;
  SIGNAL or_640_nl : STD_LOGIC;
  SIGNAL or_638_nl : STD_LOGIC;
  SIGNAL or_637_nl : STD_LOGIC;
  SIGNAL nor_591_nl : STD_LOGIC;
  SIGNAL mux_762_nl : STD_LOGIC;
  SIGNAL mux_761_nl : STD_LOGIC;
  SIGNAL nor_592_nl : STD_LOGIC;
  SIGNAL and_333_nl : STD_LOGIC;
  SIGNAL mux_760_nl : STD_LOGIC;
  SIGNAL nor_593_nl : STD_LOGIC;
  SIGNAL mux_759_nl : STD_LOGIC;
  SIGNAL nor_594_nl : STD_LOGIC;
  SIGNAL nor_595_nl : STD_LOGIC;
  SIGNAL and_334_nl : STD_LOGIC;
  SIGNAL mux_758_nl : STD_LOGIC;
  SIGNAL mux_757_nl : STD_LOGIC;
  SIGNAL mux_756_nl : STD_LOGIC;
  SIGNAL nor_596_nl : STD_LOGIC;
  SIGNAL nor_597_nl : STD_LOGIC;
  SIGNAL mux_755_nl : STD_LOGIC;
  SIGNAL nor_599_nl : STD_LOGIC;
  SIGNAL mux_754_nl : STD_LOGIC;
  SIGNAL mux_753_nl : STD_LOGIC;
  SIGNAL nor_600_nl : STD_LOGIC;
  SIGNAL nor_601_nl : STD_LOGIC;
  SIGNAL nor_602_nl : STD_LOGIC;
  SIGNAL nor_603_nl : STD_LOGIC;
  SIGNAL mux_752_nl : STD_LOGIC;
  SIGNAL nand_29_nl : STD_LOGIC;
  SIGNAL mux_751_nl : STD_LOGIC;
  SIGNAL mux_750_nl : STD_LOGIC;
  SIGNAL mux_749_nl : STD_LOGIC;
  SIGNAL nor_605_nl : STD_LOGIC;
  SIGNAL mux_748_nl : STD_LOGIC;
  SIGNAL nor_606_nl : STD_LOGIC;
  SIGNAL nor_607_nl : STD_LOGIC;
  SIGNAL nor_608_nl : STD_LOGIC;
  SIGNAL or_608_nl : STD_LOGIC;
  SIGNAL mux_747_nl : STD_LOGIC;
  SIGNAL or_607_nl : STD_LOGIC;
  SIGNAL mux_746_nl : STD_LOGIC;
  SIGNAL mux_745_nl : STD_LOGIC;
  SIGNAL or_605_nl : STD_LOGIC;
  SIGNAL or_604_nl : STD_LOGIC;
  SIGNAL mux_744_nl : STD_LOGIC;
  SIGNAL or_601_nl : STD_LOGIC;
  SIGNAL mux_804_nl : STD_LOGIC;
  SIGNAL mux_803_nl : STD_LOGIC;
  SIGNAL nor_583_nl : STD_LOGIC;
  SIGNAL mux_802_nl : STD_LOGIC;
  SIGNAL nand_34_nl : STD_LOGIC;
  SIGNAL mux_801_nl : STD_LOGIC;
  SIGNAL mux_800_nl : STD_LOGIC;
  SIGNAL or_691_nl : STD_LOGIC;
  SIGNAL mux_799_nl : STD_LOGIC;
  SIGNAL or_690_nl : STD_LOGIC;
  SIGNAL or_689_nl : STD_LOGIC;
  SIGNAL mux_798_nl : STD_LOGIC;
  SIGNAL nor_584_nl : STD_LOGIC;
  SIGNAL nor_585_nl : STD_LOGIC;
  SIGNAL mux_797_nl : STD_LOGIC;
  SIGNAL or_685_nl : STD_LOGIC;
  SIGNAL mux_796_nl : STD_LOGIC;
  SIGNAL and_332_nl : STD_LOGIC;
  SIGNAL mux_795_nl : STD_LOGIC;
  SIGNAL or_682_nl : STD_LOGIC;
  SIGNAL mux_794_nl : STD_LOGIC;
  SIGNAL mux_793_nl : STD_LOGIC;
  SIGNAL mux_792_nl : STD_LOGIC;
  SIGNAL or_680_nl : STD_LOGIC;
  SIGNAL mux_791_nl : STD_LOGIC;
  SIGNAL or_678_nl : STD_LOGIC;
  SIGNAL or_677_nl : STD_LOGIC;
  SIGNAL mux_790_nl : STD_LOGIC;
  SIGNAL or_676_nl : STD_LOGIC;
  SIGNAL nor_586_nl : STD_LOGIC;
  SIGNAL mux_789_nl : STD_LOGIC;
  SIGNAL nor_587_nl : STD_LOGIC;
  SIGNAL mux_788_nl : STD_LOGIC;
  SIGNAL mux_787_nl : STD_LOGIC;
  SIGNAL or_673_nl : STD_LOGIC;
  SIGNAL mux_786_nl : STD_LOGIC;
  SIGNAL mux_785_nl : STD_LOGIC;
  SIGNAL or_671_nl : STD_LOGIC;
  SIGNAL mux_784_nl : STD_LOGIC;
  SIGNAL or_669_nl : STD_LOGIC;
  SIGNAL mux_783_nl : STD_LOGIC;
  SIGNAL or_668_nl : STD_LOGIC;
  SIGNAL mux_782_nl : STD_LOGIC;
  SIGNAL or_667_nl : STD_LOGIC;
  SIGNAL nor_588_nl : STD_LOGIC;
  SIGNAL mux_781_nl : STD_LOGIC;
  SIGNAL nand_32_nl : STD_LOGIC;
  SIGNAL mux_780_nl : STD_LOGIC;
  SIGNAL or_664_nl : STD_LOGIC;
  SIGNAL mux_779_nl : STD_LOGIC;
  SIGNAL mux_778_nl : STD_LOGIC;
  SIGNAL or_662_nl : STD_LOGIC;
  SIGNAL mux_777_nl : STD_LOGIC;
  SIGNAL or_658_nl : STD_LOGIC;
  SIGNAL or_657_nl : STD_LOGIC;
  SIGNAL mux_776_nl : STD_LOGIC;
  SIGNAL or_656_nl : STD_LOGIC;
  SIGNAL mux_775_nl : STD_LOGIC;
  SIGNAL or_655_nl : STD_LOGIC;
  SIGNAL mux_835_nl : STD_LOGIC;
  SIGNAL mux_834_nl : STD_LOGIC;
  SIGNAL nor_563_nl : STD_LOGIC;
  SIGNAL mux_833_nl : STD_LOGIC;
  SIGNAL mux_832_nl : STD_LOGIC;
  SIGNAL or_744_nl : STD_LOGIC;
  SIGNAL mux_831_nl : STD_LOGIC;
  SIGNAL or_743_nl : STD_LOGIC;
  SIGNAL mux_830_nl : STD_LOGIC;
  SIGNAL mux_829_nl : STD_LOGIC;
  SIGNAL or_738_nl : STD_LOGIC;
  SIGNAL mux_828_nl : STD_LOGIC;
  SIGNAL or_737_nl : STD_LOGIC;
  SIGNAL or_735_nl : STD_LOGIC;
  SIGNAL mux_827_nl : STD_LOGIC;
  SIGNAL nor_564_nl : STD_LOGIC;
  SIGNAL mux_826_nl : STD_LOGIC;
  SIGNAL mux_825_nl : STD_LOGIC;
  SIGNAL or_733_nl : STD_LOGIC;
  SIGNAL or_731_nl : STD_LOGIC;
  SIGNAL or_730_nl : STD_LOGIC;
  SIGNAL nor_565_nl : STD_LOGIC;
  SIGNAL mux_824_nl : STD_LOGIC;
  SIGNAL mux_823_nl : STD_LOGIC;
  SIGNAL nor_566_nl : STD_LOGIC;
  SIGNAL and_330_nl : STD_LOGIC;
  SIGNAL mux_822_nl : STD_LOGIC;
  SIGNAL nor_567_nl : STD_LOGIC;
  SIGNAL mux_821_nl : STD_LOGIC;
  SIGNAL nor_568_nl : STD_LOGIC;
  SIGNAL nor_569_nl : STD_LOGIC;
  SIGNAL and_331_nl : STD_LOGIC;
  SIGNAL mux_820_nl : STD_LOGIC;
  SIGNAL mux_819_nl : STD_LOGIC;
  SIGNAL mux_818_nl : STD_LOGIC;
  SIGNAL nor_570_nl : STD_LOGIC;
  SIGNAL nor_571_nl : STD_LOGIC;
  SIGNAL mux_817_nl : STD_LOGIC;
  SIGNAL nor_573_nl : STD_LOGIC;
  SIGNAL mux_816_nl : STD_LOGIC;
  SIGNAL mux_815_nl : STD_LOGIC;
  SIGNAL nor_574_nl : STD_LOGIC;
  SIGNAL nor_575_nl : STD_LOGIC;
  SIGNAL nor_576_nl : STD_LOGIC;
  SIGNAL nor_577_nl : STD_LOGIC;
  SIGNAL mux_814_nl : STD_LOGIC;
  SIGNAL nand_35_nl : STD_LOGIC;
  SIGNAL mux_813_nl : STD_LOGIC;
  SIGNAL mux_812_nl : STD_LOGIC;
  SIGNAL mux_811_nl : STD_LOGIC;
  SIGNAL nor_579_nl : STD_LOGIC;
  SIGNAL mux_810_nl : STD_LOGIC;
  SIGNAL nor_580_nl : STD_LOGIC;
  SIGNAL nor_581_nl : STD_LOGIC;
  SIGNAL nor_582_nl : STD_LOGIC;
  SIGNAL or_701_nl : STD_LOGIC;
  SIGNAL mux_809_nl : STD_LOGIC;
  SIGNAL or_700_nl : STD_LOGIC;
  SIGNAL mux_808_nl : STD_LOGIC;
  SIGNAL mux_807_nl : STD_LOGIC;
  SIGNAL or_698_nl : STD_LOGIC;
  SIGNAL mux_806_nl : STD_LOGIC;
  SIGNAL or_694_nl : STD_LOGIC;
  SIGNAL mux_866_nl : STD_LOGIC;
  SIGNAL mux_865_nl : STD_LOGIC;
  SIGNAL mux_864_nl : STD_LOGIC;
  SIGNAL nor_555_nl : STD_LOGIC;
  SIGNAL mux_863_nl : STD_LOGIC;
  SIGNAL mux_862_nl : STD_LOGIC;
  SIGNAL or_785_nl : STD_LOGIC;
  SIGNAL mux_861_nl : STD_LOGIC;
  SIGNAL or_784_nl : STD_LOGIC;
  SIGNAL and_329_nl : STD_LOGIC;
  SIGNAL mux_860_nl : STD_LOGIC;
  SIGNAL or_782_nl : STD_LOGIC;
  SIGNAL mux_859_nl : STD_LOGIC;
  SIGNAL mux_858_nl : STD_LOGIC;
  SIGNAL or_781_nl : STD_LOGIC;
  SIGNAL mux_857_nl : STD_LOGIC;
  SIGNAL or_780_nl : STD_LOGIC;
  SIGNAL nor_556_nl : STD_LOGIC;
  SIGNAL mux_856_nl : STD_LOGIC;
  SIGNAL or_777_nl : STD_LOGIC;
  SIGNAL nor_557_nl : STD_LOGIC;
  SIGNAL mux_855_nl : STD_LOGIC;
  SIGNAL mux_854_nl : STD_LOGIC;
  SIGNAL or_774_nl : STD_LOGIC;
  SIGNAL or_773_nl : STD_LOGIC;
  SIGNAL nand_38_nl : STD_LOGIC;
  SIGNAL mux_853_nl : STD_LOGIC;
  SIGNAL or_772_nl : STD_LOGIC;
  SIGNAL mux_852_nl : STD_LOGIC;
  SIGNAL or_771_nl : STD_LOGIC;
  SIGNAL mux_851_nl : STD_LOGIC;
  SIGNAL mux_850_nl : STD_LOGIC;
  SIGNAL nor_558_nl : STD_LOGIC;
  SIGNAL mux_849_nl : STD_LOGIC;
  SIGNAL nor_559_nl : STD_LOGIC;
  SIGNAL nor_560_nl : STD_LOGIC;
  SIGNAL mux_848_nl : STD_LOGIC;
  SIGNAL or_766_nl : STD_LOGIC;
  SIGNAL mux_847_nl : STD_LOGIC;
  SIGNAL or_765_nl : STD_LOGIC;
  SIGNAL mux_846_nl : STD_LOGIC;
  SIGNAL nor_561_nl : STD_LOGIC;
  SIGNAL mux_845_nl : STD_LOGIC;
  SIGNAL or_761_nl : STD_LOGIC;
  SIGNAL mux_844_nl : STD_LOGIC;
  SIGNAL mux_843_nl : STD_LOGIC;
  SIGNAL or_760_nl : STD_LOGIC;
  SIGNAL mux_842_nl : STD_LOGIC;
  SIGNAL or_759_nl : STD_LOGIC;
  SIGNAL nor_562_nl : STD_LOGIC;
  SIGNAL mux_841_nl : STD_LOGIC;
  SIGNAL mux_840_nl : STD_LOGIC;
  SIGNAL mux_839_nl : STD_LOGIC;
  SIGNAL or_755_nl : STD_LOGIC;
  SIGNAL mux_838_nl : STD_LOGIC;
  SIGNAL or_752_nl : STD_LOGIC;
  SIGNAL or_750_nl : STD_LOGIC;
  SIGNAL mux_837_nl : STD_LOGIC;
  SIGNAL or_749_nl : STD_LOGIC;
  SIGNAL mux_897_nl : STD_LOGIC;
  SIGNAL mux_896_nl : STD_LOGIC;
  SIGNAL nor_535_nl : STD_LOGIC;
  SIGNAL mux_895_nl : STD_LOGIC;
  SIGNAL mux_894_nl : STD_LOGIC;
  SIGNAL or_837_nl : STD_LOGIC;
  SIGNAL mux_893_nl : STD_LOGIC;
  SIGNAL or_836_nl : STD_LOGIC;
  SIGNAL mux_892_nl : STD_LOGIC;
  SIGNAL mux_891_nl : STD_LOGIC;
  SIGNAL or_833_nl : STD_LOGIC;
  SIGNAL or_831_nl : STD_LOGIC;
  SIGNAL mux_890_nl : STD_LOGIC;
  SIGNAL or_830_nl : STD_LOGIC;
  SIGNAL or_828_nl : STD_LOGIC;
  SIGNAL mux_889_nl : STD_LOGIC;
  SIGNAL nor_536_nl : STD_LOGIC;
  SIGNAL mux_888_nl : STD_LOGIC;
  SIGNAL mux_887_nl : STD_LOGIC;
  SIGNAL or_826_nl : STD_LOGIC;
  SIGNAL or_824_nl : STD_LOGIC;
  SIGNAL or_823_nl : STD_LOGIC;
  SIGNAL nor_537_nl : STD_LOGIC;
  SIGNAL mux_886_nl : STD_LOGIC;
  SIGNAL mux_885_nl : STD_LOGIC;
  SIGNAL nor_538_nl : STD_LOGIC;
  SIGNAL and_327_nl : STD_LOGIC;
  SIGNAL mux_884_nl : STD_LOGIC;
  SIGNAL nor_539_nl : STD_LOGIC;
  SIGNAL mux_883_nl : STD_LOGIC;
  SIGNAL nor_540_nl : STD_LOGIC;
  SIGNAL nor_541_nl : STD_LOGIC;
  SIGNAL and_328_nl : STD_LOGIC;
  SIGNAL mux_882_nl : STD_LOGIC;
  SIGNAL mux_881_nl : STD_LOGIC;
  SIGNAL mux_880_nl : STD_LOGIC;
  SIGNAL nor_542_nl : STD_LOGIC;
  SIGNAL nor_543_nl : STD_LOGIC;
  SIGNAL mux_879_nl : STD_LOGIC;
  SIGNAL nor_545_nl : STD_LOGIC;
  SIGNAL mux_878_nl : STD_LOGIC;
  SIGNAL mux_877_nl : STD_LOGIC;
  SIGNAL nor_546_nl : STD_LOGIC;
  SIGNAL nor_547_nl : STD_LOGIC;
  SIGNAL nor_548_nl : STD_LOGIC;
  SIGNAL nor_549_nl : STD_LOGIC;
  SIGNAL mux_876_nl : STD_LOGIC;
  SIGNAL nand_41_nl : STD_LOGIC;
  SIGNAL mux_875_nl : STD_LOGIC;
  SIGNAL mux_874_nl : STD_LOGIC;
  SIGNAL mux_873_nl : STD_LOGIC;
  SIGNAL nor_551_nl : STD_LOGIC;
  SIGNAL mux_872_nl : STD_LOGIC;
  SIGNAL nor_552_nl : STD_LOGIC;
  SIGNAL nor_553_nl : STD_LOGIC;
  SIGNAL nor_554_nl : STD_LOGIC;
  SIGNAL or_794_nl : STD_LOGIC;
  SIGNAL mux_871_nl : STD_LOGIC;
  SIGNAL or_793_nl : STD_LOGIC;
  SIGNAL mux_870_nl : STD_LOGIC;
  SIGNAL mux_869_nl : STD_LOGIC;
  SIGNAL or_791_nl : STD_LOGIC;
  SIGNAL or_790_nl : STD_LOGIC;
  SIGNAL mux_868_nl : STD_LOGIC;
  SIGNAL or_787_nl : STD_LOGIC;
  SIGNAL mux_928_nl : STD_LOGIC;
  SIGNAL mux_927_nl : STD_LOGIC;
  SIGNAL nor_529_nl : STD_LOGIC;
  SIGNAL mux_926_nl : STD_LOGIC;
  SIGNAL nand_46_nl : STD_LOGIC;
  SIGNAL mux_925_nl : STD_LOGIC;
  SIGNAL mux_924_nl : STD_LOGIC;
  SIGNAL or_877_nl : STD_LOGIC;
  SIGNAL mux_923_nl : STD_LOGIC;
  SIGNAL or_876_nl : STD_LOGIC;
  SIGNAL or_875_nl : STD_LOGIC;
  SIGNAL mux_922_nl : STD_LOGIC;
  SIGNAL and_438_nl : STD_LOGIC;
  SIGNAL nor_531_nl : STD_LOGIC;
  SIGNAL mux_921_nl : STD_LOGIC;
  SIGNAL or_871_nl : STD_LOGIC;
  SIGNAL mux_920_nl : STD_LOGIC;
  SIGNAL and_326_nl : STD_LOGIC;
  SIGNAL mux_919_nl : STD_LOGIC;
  SIGNAL or_868_nl : STD_LOGIC;
  SIGNAL mux_918_nl : STD_LOGIC;
  SIGNAL mux_917_nl : STD_LOGIC;
  SIGNAL mux_916_nl : STD_LOGIC;
  SIGNAL or_866_nl : STD_LOGIC;
  SIGNAL mux_915_nl : STD_LOGIC;
  SIGNAL or_864_nl : STD_LOGIC;
  SIGNAL or_863_nl : STD_LOGIC;
  SIGNAL mux_914_nl : STD_LOGIC;
  SIGNAL or_862_nl : STD_LOGIC;
  SIGNAL nor_532_nl : STD_LOGIC;
  SIGNAL mux_913_nl : STD_LOGIC;
  SIGNAL nor_533_nl : STD_LOGIC;
  SIGNAL mux_912_nl : STD_LOGIC;
  SIGNAL mux_911_nl : STD_LOGIC;
  SIGNAL or_859_nl : STD_LOGIC;
  SIGNAL mux_910_nl : STD_LOGIC;
  SIGNAL mux_909_nl : STD_LOGIC;
  SIGNAL or_857_nl : STD_LOGIC;
  SIGNAL mux_908_nl : STD_LOGIC;
  SIGNAL or_855_nl : STD_LOGIC;
  SIGNAL mux_907_nl : STD_LOGIC;
  SIGNAL or_854_nl : STD_LOGIC;
  SIGNAL mux_906_nl : STD_LOGIC;
  SIGNAL or_853_nl : STD_LOGIC;
  SIGNAL nor_534_nl : STD_LOGIC;
  SIGNAL mux_905_nl : STD_LOGIC;
  SIGNAL nand_44_nl : STD_LOGIC;
  SIGNAL mux_904_nl : STD_LOGIC;
  SIGNAL or_850_nl : STD_LOGIC;
  SIGNAL mux_903_nl : STD_LOGIC;
  SIGNAL mux_902_nl : STD_LOGIC;
  SIGNAL or_848_nl : STD_LOGIC;
  SIGNAL mux_901_nl : STD_LOGIC;
  SIGNAL or_844_nl : STD_LOGIC;
  SIGNAL or_843_nl : STD_LOGIC;
  SIGNAL mux_900_nl : STD_LOGIC;
  SIGNAL or_842_nl : STD_LOGIC;
  SIGNAL mux_899_nl : STD_LOGIC;
  SIGNAL or_841_nl : STD_LOGIC;
  SIGNAL mux_959_nl : STD_LOGIC;
  SIGNAL mux_958_nl : STD_LOGIC;
  SIGNAL nor_509_nl : STD_LOGIC;
  SIGNAL mux_957_nl : STD_LOGIC;
  SIGNAL mux_956_nl : STD_LOGIC;
  SIGNAL or_930_nl : STD_LOGIC;
  SIGNAL mux_955_nl : STD_LOGIC;
  SIGNAL or_929_nl : STD_LOGIC;
  SIGNAL mux_954_nl : STD_LOGIC;
  SIGNAL mux_953_nl : STD_LOGIC;
  SIGNAL or_924_nl : STD_LOGIC;
  SIGNAL mux_952_nl : STD_LOGIC;
  SIGNAL or_923_nl : STD_LOGIC;
  SIGNAL or_921_nl : STD_LOGIC;
  SIGNAL mux_951_nl : STD_LOGIC;
  SIGNAL nor_510_nl : STD_LOGIC;
  SIGNAL mux_950_nl : STD_LOGIC;
  SIGNAL mux_949_nl : STD_LOGIC;
  SIGNAL or_919_nl : STD_LOGIC;
  SIGNAL or_917_nl : STD_LOGIC;
  SIGNAL or_916_nl : STD_LOGIC;
  SIGNAL nor_511_nl : STD_LOGIC;
  SIGNAL mux_948_nl : STD_LOGIC;
  SIGNAL mux_947_nl : STD_LOGIC;
  SIGNAL nor_512_nl : STD_LOGIC;
  SIGNAL and_324_nl : STD_LOGIC;
  SIGNAL mux_946_nl : STD_LOGIC;
  SIGNAL nor_513_nl : STD_LOGIC;
  SIGNAL mux_945_nl : STD_LOGIC;
  SIGNAL nor_514_nl : STD_LOGIC;
  SIGNAL nor_515_nl : STD_LOGIC;
  SIGNAL and_325_nl : STD_LOGIC;
  SIGNAL mux_944_nl : STD_LOGIC;
  SIGNAL mux_943_nl : STD_LOGIC;
  SIGNAL mux_942_nl : STD_LOGIC;
  SIGNAL nor_516_nl : STD_LOGIC;
  SIGNAL nor_517_nl : STD_LOGIC;
  SIGNAL mux_941_nl : STD_LOGIC;
  SIGNAL nor_519_nl : STD_LOGIC;
  SIGNAL mux_940_nl : STD_LOGIC;
  SIGNAL mux_939_nl : STD_LOGIC;
  SIGNAL nor_520_nl : STD_LOGIC;
  SIGNAL nor_521_nl : STD_LOGIC;
  SIGNAL nor_522_nl : STD_LOGIC;
  SIGNAL nor_523_nl : STD_LOGIC;
  SIGNAL mux_938_nl : STD_LOGIC;
  SIGNAL nand_47_nl : STD_LOGIC;
  SIGNAL mux_937_nl : STD_LOGIC;
  SIGNAL mux_936_nl : STD_LOGIC;
  SIGNAL mux_935_nl : STD_LOGIC;
  SIGNAL nor_525_nl : STD_LOGIC;
  SIGNAL mux_934_nl : STD_LOGIC;
  SIGNAL nor_526_nl : STD_LOGIC;
  SIGNAL nor_527_nl : STD_LOGIC;
  SIGNAL nor_528_nl : STD_LOGIC;
  SIGNAL or_887_nl : STD_LOGIC;
  SIGNAL mux_933_nl : STD_LOGIC;
  SIGNAL or_886_nl : STD_LOGIC;
  SIGNAL mux_932_nl : STD_LOGIC;
  SIGNAL mux_931_nl : STD_LOGIC;
  SIGNAL or_884_nl : STD_LOGIC;
  SIGNAL mux_930_nl : STD_LOGIC;
  SIGNAL or_880_nl : STD_LOGIC;
  SIGNAL mux_990_nl : STD_LOGIC;
  SIGNAL mux_989_nl : STD_LOGIC;
  SIGNAL nor_503_nl : STD_LOGIC;
  SIGNAL mux_988_nl : STD_LOGIC;
  SIGNAL nand_52_nl : STD_LOGIC;
  SIGNAL mux_987_nl : STD_LOGIC;
  SIGNAL mux_986_nl : STD_LOGIC;
  SIGNAL or_970_nl : STD_LOGIC;
  SIGNAL mux_985_nl : STD_LOGIC;
  SIGNAL or_969_nl : STD_LOGIC;
  SIGNAL or_968_nl : STD_LOGIC;
  SIGNAL mux_984_nl : STD_LOGIC;
  SIGNAL and_437_nl : STD_LOGIC;
  SIGNAL nor_505_nl : STD_LOGIC;
  SIGNAL mux_983_nl : STD_LOGIC;
  SIGNAL or_964_nl : STD_LOGIC;
  SIGNAL mux_982_nl : STD_LOGIC;
  SIGNAL and_323_nl : STD_LOGIC;
  SIGNAL mux_981_nl : STD_LOGIC;
  SIGNAL nand_376_nl : STD_LOGIC;
  SIGNAL mux_980_nl : STD_LOGIC;
  SIGNAL mux_979_nl : STD_LOGIC;
  SIGNAL mux_978_nl : STD_LOGIC;
  SIGNAL or_959_nl : STD_LOGIC;
  SIGNAL mux_977_nl : STD_LOGIC;
  SIGNAL or_957_nl : STD_LOGIC;
  SIGNAL or_956_nl : STD_LOGIC;
  SIGNAL mux_976_nl : STD_LOGIC;
  SIGNAL or_955_nl : STD_LOGIC;
  SIGNAL nor_506_nl : STD_LOGIC;
  SIGNAL mux_975_nl : STD_LOGIC;
  SIGNAL nor_507_nl : STD_LOGIC;
  SIGNAL mux_974_nl : STD_LOGIC;
  SIGNAL mux_973_nl : STD_LOGIC;
  SIGNAL nand_371_nl : STD_LOGIC;
  SIGNAL mux_972_nl : STD_LOGIC;
  SIGNAL mux_971_nl : STD_LOGIC;
  SIGNAL or_950_nl : STD_LOGIC;
  SIGNAL mux_970_nl : STD_LOGIC;
  SIGNAL or_948_nl : STD_LOGIC;
  SIGNAL mux_969_nl : STD_LOGIC;
  SIGNAL or_947_nl : STD_LOGIC;
  SIGNAL mux_968_nl : STD_LOGIC;
  SIGNAL or_946_nl : STD_LOGIC;
  SIGNAL nor_508_nl : STD_LOGIC;
  SIGNAL mux_967_nl : STD_LOGIC;
  SIGNAL nand_50_nl : STD_LOGIC;
  SIGNAL mux_966_nl : STD_LOGIC;
  SIGNAL nand_360_nl : STD_LOGIC;
  SIGNAL mux_965_nl : STD_LOGIC;
  SIGNAL mux_964_nl : STD_LOGIC;
  SIGNAL or_941_nl : STD_LOGIC;
  SIGNAL mux_963_nl : STD_LOGIC;
  SIGNAL or_937_nl : STD_LOGIC;
  SIGNAL or_936_nl : STD_LOGIC;
  SIGNAL mux_962_nl : STD_LOGIC;
  SIGNAL or_935_nl : STD_LOGIC;
  SIGNAL mux_961_nl : STD_LOGIC;
  SIGNAL or_934_nl : STD_LOGIC;
  SIGNAL mux_1021_nl : STD_LOGIC;
  SIGNAL mux_1020_nl : STD_LOGIC;
  SIGNAL nor_484_nl : STD_LOGIC;
  SIGNAL mux_1019_nl : STD_LOGIC;
  SIGNAL mux_1018_nl : STD_LOGIC;
  SIGNAL nand_274_nl : STD_LOGIC;
  SIGNAL mux_1017_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL mux_1016_nl : STD_LOGIC;
  SIGNAL mux_1015_nl : STD_LOGIC;
  SIGNAL or_1019_nl : STD_LOGIC;
  SIGNAL or_1017_nl : STD_LOGIC;
  SIGNAL mux_1014_nl : STD_LOGIC;
  SIGNAL nand_370_nl : STD_LOGIC;
  SIGNAL or_1014_nl : STD_LOGIC;
  SIGNAL mux_1013_nl : STD_LOGIC;
  SIGNAL nor_485_nl : STD_LOGIC;
  SIGNAL mux_1012_nl : STD_LOGIC;
  SIGNAL mux_1011_nl : STD_LOGIC;
  SIGNAL or_1012_nl : STD_LOGIC;
  SIGNAL or_1010_nl : STD_LOGIC;
  SIGNAL or_1009_nl : STD_LOGIC;
  SIGNAL nor_486_nl : STD_LOGIC;
  SIGNAL mux_1010_nl : STD_LOGIC;
  SIGNAL mux_1009_nl : STD_LOGIC;
  SIGNAL nor_487_nl : STD_LOGIC;
  SIGNAL and_320_nl : STD_LOGIC;
  SIGNAL mux_1008_nl : STD_LOGIC;
  SIGNAL nor_488_nl : STD_LOGIC;
  SIGNAL mux_1007_nl : STD_LOGIC;
  SIGNAL and_321_nl : STD_LOGIC;
  SIGNAL nor_489_nl : STD_LOGIC;
  SIGNAL and_322_nl : STD_LOGIC;
  SIGNAL mux_1006_nl : STD_LOGIC;
  SIGNAL mux_1005_nl : STD_LOGIC;
  SIGNAL mux_1004_nl : STD_LOGIC;
  SIGNAL nor_490_nl : STD_LOGIC;
  SIGNAL nor_491_nl : STD_LOGIC;
  SIGNAL mux_1003_nl : STD_LOGIC;
  SIGNAL nor_493_nl : STD_LOGIC;
  SIGNAL mux_1002_nl : STD_LOGIC;
  SIGNAL mux_1001_nl : STD_LOGIC;
  SIGNAL nor_494_nl : STD_LOGIC;
  SIGNAL and_432_nl : STD_LOGIC;
  SIGNAL nor_496_nl : STD_LOGIC;
  SIGNAL nor_497_nl : STD_LOGIC;
  SIGNAL mux_1000_nl : STD_LOGIC;
  SIGNAL nand_53_nl : STD_LOGIC;
  SIGNAL mux_999_nl : STD_LOGIC;
  SIGNAL mux_998_nl : STD_LOGIC;
  SIGNAL mux_997_nl : STD_LOGIC;
  SIGNAL nor_499_nl : STD_LOGIC;
  SIGNAL mux_996_nl : STD_LOGIC;
  SIGNAL nor_500_nl : STD_LOGIC;
  SIGNAL nor_501_nl : STD_LOGIC;
  SIGNAL nor_502_nl : STD_LOGIC;
  SIGNAL or_980_nl : STD_LOGIC;
  SIGNAL mux_995_nl : STD_LOGIC;
  SIGNAL or_979_nl : STD_LOGIC;
  SIGNAL mux_994_nl : STD_LOGIC;
  SIGNAL mux_993_nl : STD_LOGIC;
  SIGNAL nand_282_nl : STD_LOGIC;
  SIGNAL or_976_nl : STD_LOGIC;
  SIGNAL mux_992_nl : STD_LOGIC;
  SIGNAL nand_354_nl : STD_LOGIC;
  SIGNAL mux_1052_nl : STD_LOGIC;
  SIGNAL mux_1051_nl : STD_LOGIC;
  SIGNAL nor_478_nl : STD_LOGIC;
  SIGNAL mux_1050_nl : STD_LOGIC;
  SIGNAL nand_58_nl : STD_LOGIC;
  SIGNAL mux_1049_nl : STD_LOGIC;
  SIGNAL mux_1048_nl : STD_LOGIC;
  SIGNAL or_1069_nl : STD_LOGIC;
  SIGNAL mux_1047_nl : STD_LOGIC;
  SIGNAL or_1068_nl : STD_LOGIC;
  SIGNAL or_1067_nl : STD_LOGIC;
  SIGNAL mux_1046_nl : STD_LOGIC;
  SIGNAL nor_479_nl : STD_LOGIC;
  SIGNAL nor_480_nl : STD_LOGIC;
  SIGNAL mux_1045_nl : STD_LOGIC;
  SIGNAL or_1062_nl : STD_LOGIC;
  SIGNAL mux_1044_nl : STD_LOGIC;
  SIGNAL and_319_nl : STD_LOGIC;
  SIGNAL mux_1043_nl : STD_LOGIC;
  SIGNAL or_1059_nl : STD_LOGIC;
  SIGNAL mux_1042_nl : STD_LOGIC;
  SIGNAL mux_1041_nl : STD_LOGIC;
  SIGNAL mux_1040_nl : STD_LOGIC;
  SIGNAL or_1057_nl : STD_LOGIC;
  SIGNAL mux_1039_nl : STD_LOGIC;
  SIGNAL or_1055_nl : STD_LOGIC;
  SIGNAL or_1054_nl : STD_LOGIC;
  SIGNAL mux_1038_nl : STD_LOGIC;
  SIGNAL or_1053_nl : STD_LOGIC;
  SIGNAL nor_481_nl : STD_LOGIC;
  SIGNAL mux_1037_nl : STD_LOGIC;
  SIGNAL nor_482_nl : STD_LOGIC;
  SIGNAL mux_1036_nl : STD_LOGIC;
  SIGNAL mux_1035_nl : STD_LOGIC;
  SIGNAL or_1049_nl : STD_LOGIC;
  SIGNAL mux_1034_nl : STD_LOGIC;
  SIGNAL mux_1033_nl : STD_LOGIC;
  SIGNAL or_1047_nl : STD_LOGIC;
  SIGNAL mux_1032_nl : STD_LOGIC;
  SIGNAL or_1045_nl : STD_LOGIC;
  SIGNAL mux_1031_nl : STD_LOGIC;
  SIGNAL or_1044_nl : STD_LOGIC;
  SIGNAL mux_1030_nl : STD_LOGIC;
  SIGNAL or_1043_nl : STD_LOGIC;
  SIGNAL nor_483_nl : STD_LOGIC;
  SIGNAL mux_1029_nl : STD_LOGIC;
  SIGNAL nand_56_nl : STD_LOGIC;
  SIGNAL mux_1028_nl : STD_LOGIC;
  SIGNAL or_1040_nl : STD_LOGIC;
  SIGNAL mux_1027_nl : STD_LOGIC;
  SIGNAL mux_1026_nl : STD_LOGIC;
  SIGNAL or_1038_nl : STD_LOGIC;
  SIGNAL mux_1025_nl : STD_LOGIC;
  SIGNAL or_1032_nl : STD_LOGIC;
  SIGNAL or_1031_nl : STD_LOGIC;
  SIGNAL mux_1024_nl : STD_LOGIC;
  SIGNAL or_1030_nl : STD_LOGIC;
  SIGNAL mux_1023_nl : STD_LOGIC;
  SIGNAL or_1029_nl : STD_LOGIC;
  SIGNAL mux_1083_nl : STD_LOGIC;
  SIGNAL mux_1082_nl : STD_LOGIC;
  SIGNAL nor_458_nl : STD_LOGIC;
  SIGNAL mux_1081_nl : STD_LOGIC;
  SIGNAL mux_1080_nl : STD_LOGIC;
  SIGNAL or_1122_nl : STD_LOGIC;
  SIGNAL mux_1079_nl : STD_LOGIC;
  SIGNAL or_1121_nl : STD_LOGIC;
  SIGNAL mux_1078_nl : STD_LOGIC;
  SIGNAL mux_1077_nl : STD_LOGIC;
  SIGNAL or_1118_nl : STD_LOGIC;
  SIGNAL or_1116_nl : STD_LOGIC;
  SIGNAL mux_1076_nl : STD_LOGIC;
  SIGNAL or_1115_nl : STD_LOGIC;
  SIGNAL or_1113_nl : STD_LOGIC;
  SIGNAL mux_1075_nl : STD_LOGIC;
  SIGNAL nor_459_nl : STD_LOGIC;
  SIGNAL mux_1074_nl : STD_LOGIC;
  SIGNAL mux_1073_nl : STD_LOGIC;
  SIGNAL or_1111_nl : STD_LOGIC;
  SIGNAL or_1109_nl : STD_LOGIC;
  SIGNAL or_1108_nl : STD_LOGIC;
  SIGNAL nor_460_nl : STD_LOGIC;
  SIGNAL mux_1072_nl : STD_LOGIC;
  SIGNAL mux_1071_nl : STD_LOGIC;
  SIGNAL nor_461_nl : STD_LOGIC;
  SIGNAL and_317_nl : STD_LOGIC;
  SIGNAL mux_1070_nl : STD_LOGIC;
  SIGNAL nor_462_nl : STD_LOGIC;
  SIGNAL mux_1069_nl : STD_LOGIC;
  SIGNAL nor_463_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL and_318_nl : STD_LOGIC;
  SIGNAL mux_1068_nl : STD_LOGIC;
  SIGNAL mux_1067_nl : STD_LOGIC;
  SIGNAL mux_1066_nl : STD_LOGIC;
  SIGNAL nor_465_nl : STD_LOGIC;
  SIGNAL nor_466_nl : STD_LOGIC;
  SIGNAL mux_1065_nl : STD_LOGIC;
  SIGNAL nor_468_nl : STD_LOGIC;
  SIGNAL mux_1064_nl : STD_LOGIC;
  SIGNAL mux_1063_nl : STD_LOGIC;
  SIGNAL nor_469_nl : STD_LOGIC;
  SIGNAL nor_470_nl : STD_LOGIC;
  SIGNAL nor_471_nl : STD_LOGIC;
  SIGNAL nor_472_nl : STD_LOGIC;
  SIGNAL mux_1062_nl : STD_LOGIC;
  SIGNAL nand_59_nl : STD_LOGIC;
  SIGNAL mux_1061_nl : STD_LOGIC;
  SIGNAL mux_1060_nl : STD_LOGIC;
  SIGNAL mux_1059_nl : STD_LOGIC;
  SIGNAL nor_474_nl : STD_LOGIC;
  SIGNAL mux_1058_nl : STD_LOGIC;
  SIGNAL nor_475_nl : STD_LOGIC;
  SIGNAL nor_476_nl : STD_LOGIC;
  SIGNAL nor_477_nl : STD_LOGIC;
  SIGNAL or_1079_nl : STD_LOGIC;
  SIGNAL mux_1057_nl : STD_LOGIC;
  SIGNAL or_1078_nl : STD_LOGIC;
  SIGNAL mux_1056_nl : STD_LOGIC;
  SIGNAL mux_1055_nl : STD_LOGIC;
  SIGNAL or_1076_nl : STD_LOGIC;
  SIGNAL or_1075_nl : STD_LOGIC;
  SIGNAL mux_1054_nl : STD_LOGIC;
  SIGNAL or_1072_nl : STD_LOGIC;
  SIGNAL mux_1114_nl : STD_LOGIC;
  SIGNAL mux_1113_nl : STD_LOGIC;
  SIGNAL mux_1112_nl : STD_LOGIC;
  SIGNAL nor_450_nl : STD_LOGIC;
  SIGNAL mux_1111_nl : STD_LOGIC;
  SIGNAL mux_1110_nl : STD_LOGIC;
  SIGNAL or_1169_nl : STD_LOGIC;
  SIGNAL mux_1109_nl : STD_LOGIC;
  SIGNAL or_1168_nl : STD_LOGIC;
  SIGNAL and_316_nl : STD_LOGIC;
  SIGNAL mux_1108_nl : STD_LOGIC;
  SIGNAL or_1166_nl : STD_LOGIC;
  SIGNAL mux_1107_nl : STD_LOGIC;
  SIGNAL mux_1106_nl : STD_LOGIC;
  SIGNAL or_1165_nl : STD_LOGIC;
  SIGNAL mux_1105_nl : STD_LOGIC;
  SIGNAL or_1164_nl : STD_LOGIC;
  SIGNAL nor_451_nl : STD_LOGIC;
  SIGNAL mux_1104_nl : STD_LOGIC;
  SIGNAL or_1161_nl : STD_LOGIC;
  SIGNAL nor_452_nl : STD_LOGIC;
  SIGNAL mux_1103_nl : STD_LOGIC;
  SIGNAL mux_1102_nl : STD_LOGIC;
  SIGNAL or_1158_nl : STD_LOGIC;
  SIGNAL or_1156_nl : STD_LOGIC;
  SIGNAL nand_62_nl : STD_LOGIC;
  SIGNAL mux_1101_nl : STD_LOGIC;
  SIGNAL or_1155_nl : STD_LOGIC;
  SIGNAL mux_1100_nl : STD_LOGIC;
  SIGNAL or_1154_nl : STD_LOGIC;
  SIGNAL mux_1099_nl : STD_LOGIC;
  SIGNAL mux_1098_nl : STD_LOGIC;
  SIGNAL nor_453_nl : STD_LOGIC;
  SIGNAL mux_1097_nl : STD_LOGIC;
  SIGNAL nor_454_nl : STD_LOGIC;
  SIGNAL nor_455_nl : STD_LOGIC;
  SIGNAL mux_1096_nl : STD_LOGIC;
  SIGNAL or_1148_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL or_1147_nl : STD_LOGIC;
  SIGNAL mux_1094_nl : STD_LOGIC;
  SIGNAL nor_456_nl : STD_LOGIC;
  SIGNAL mux_1093_nl : STD_LOGIC;
  SIGNAL or_1142_nl : STD_LOGIC;
  SIGNAL mux_1092_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL or_1141_nl : STD_LOGIC;
  SIGNAL mux_1090_nl : STD_LOGIC;
  SIGNAL or_1140_nl : STD_LOGIC;
  SIGNAL nor_457_nl : STD_LOGIC;
  SIGNAL mux_1089_nl : STD_LOGIC;
  SIGNAL mux_1088_nl : STD_LOGIC;
  SIGNAL mux_1087_nl : STD_LOGIC;
  SIGNAL or_1136_nl : STD_LOGIC;
  SIGNAL mux_1086_nl : STD_LOGIC;
  SIGNAL or_1131_nl : STD_LOGIC;
  SIGNAL or_1129_nl : STD_LOGIC;
  SIGNAL mux_1085_nl : STD_LOGIC;
  SIGNAL or_1128_nl : STD_LOGIC;
  SIGNAL mux_1145_nl : STD_LOGIC;
  SIGNAL mux_1144_nl : STD_LOGIC;
  SIGNAL nor_430_nl : STD_LOGIC;
  SIGNAL mux_1143_nl : STD_LOGIC;
  SIGNAL mux_1142_nl : STD_LOGIC;
  SIGNAL or_1221_nl : STD_LOGIC;
  SIGNAL mux_1141_nl : STD_LOGIC;
  SIGNAL or_1220_nl : STD_LOGIC;
  SIGNAL mux_1140_nl : STD_LOGIC;
  SIGNAL mux_1139_nl : STD_LOGIC;
  SIGNAL or_1217_nl : STD_LOGIC;
  SIGNAL or_1215_nl : STD_LOGIC;
  SIGNAL mux_1138_nl : STD_LOGIC;
  SIGNAL or_1214_nl : STD_LOGIC;
  SIGNAL or_1212_nl : STD_LOGIC;
  SIGNAL mux_1137_nl : STD_LOGIC;
  SIGNAL nor_431_nl : STD_LOGIC;
  SIGNAL mux_1136_nl : STD_LOGIC;
  SIGNAL mux_1135_nl : STD_LOGIC;
  SIGNAL or_1210_nl : STD_LOGIC;
  SIGNAL or_1208_nl : STD_LOGIC;
  SIGNAL or_1207_nl : STD_LOGIC;
  SIGNAL nor_432_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL nor_433_nl : STD_LOGIC;
  SIGNAL and_314_nl : STD_LOGIC;
  SIGNAL mux_1132_nl : STD_LOGIC;
  SIGNAL nor_434_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL nor_435_nl : STD_LOGIC;
  SIGNAL nor_436_nl : STD_LOGIC;
  SIGNAL and_315_nl : STD_LOGIC;
  SIGNAL mux_1130_nl : STD_LOGIC;
  SIGNAL mux_1129_nl : STD_LOGIC;
  SIGNAL mux_1128_nl : STD_LOGIC;
  SIGNAL nor_437_nl : STD_LOGIC;
  SIGNAL nor_438_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL nor_440_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL mux_1125_nl : STD_LOGIC;
  SIGNAL nor_441_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL nor_443_nl : STD_LOGIC;
  SIGNAL nor_444_nl : STD_LOGIC;
  SIGNAL mux_1124_nl : STD_LOGIC;
  SIGNAL nand_65_nl : STD_LOGIC;
  SIGNAL mux_1123_nl : STD_LOGIC;
  SIGNAL mux_1122_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL nor_446_nl : STD_LOGIC;
  SIGNAL mux_1120_nl : STD_LOGIC;
  SIGNAL nor_447_nl : STD_LOGIC;
  SIGNAL nor_448_nl : STD_LOGIC;
  SIGNAL nor_449_nl : STD_LOGIC;
  SIGNAL or_1178_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL or_1177_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL or_1175_nl : STD_LOGIC;
  SIGNAL or_1174_nl : STD_LOGIC;
  SIGNAL mux_1116_nl : STD_LOGIC;
  SIGNAL or_1171_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL mux_1175_nl : STD_LOGIC;
  SIGNAL nor_424_nl : STD_LOGIC;
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL nand_70_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL mux_1172_nl : STD_LOGIC;
  SIGNAL or_1267_nl : STD_LOGIC;
  SIGNAL mux_1171_nl : STD_LOGIC;
  SIGNAL or_1266_nl : STD_LOGIC;
  SIGNAL or_1265_nl : STD_LOGIC;
  SIGNAL mux_1170_nl : STD_LOGIC;
  SIGNAL and_442_nl : STD_LOGIC;
  SIGNAL nor_426_nl : STD_LOGIC;
  SIGNAL mux_1169_nl : STD_LOGIC;
  SIGNAL or_1260_nl : STD_LOGIC;
  SIGNAL mux_1168_nl : STD_LOGIC;
  SIGNAL and_313_nl : STD_LOGIC;
  SIGNAL mux_1167_nl : STD_LOGIC;
  SIGNAL or_1257_nl : STD_LOGIC;
  SIGNAL mux_1166_nl : STD_LOGIC;
  SIGNAL mux_1165_nl : STD_LOGIC;
  SIGNAL mux_1164_nl : STD_LOGIC;
  SIGNAL or_1255_nl : STD_LOGIC;
  SIGNAL mux_1163_nl : STD_LOGIC;
  SIGNAL or_1253_nl : STD_LOGIC;
  SIGNAL or_1252_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL or_1251_nl : STD_LOGIC;
  SIGNAL nor_427_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL nor_428_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL mux_1159_nl : STD_LOGIC;
  SIGNAL or_1247_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL mux_1157_nl : STD_LOGIC;
  SIGNAL or_1245_nl : STD_LOGIC;
  SIGNAL mux_1156_nl : STD_LOGIC;
  SIGNAL or_1243_nl : STD_LOGIC;
  SIGNAL mux_1155_nl : STD_LOGIC;
  SIGNAL or_1242_nl : STD_LOGIC;
  SIGNAL mux_1154_nl : STD_LOGIC;
  SIGNAL or_1241_nl : STD_LOGIC;
  SIGNAL nor_429_nl : STD_LOGIC;
  SIGNAL mux_1153_nl : STD_LOGIC;
  SIGNAL nand_68_nl : STD_LOGIC;
  SIGNAL mux_1152_nl : STD_LOGIC;
  SIGNAL or_1238_nl : STD_LOGIC;
  SIGNAL mux_1151_nl : STD_LOGIC;
  SIGNAL mux_1150_nl : STD_LOGIC;
  SIGNAL or_1236_nl : STD_LOGIC;
  SIGNAL mux_1149_nl : STD_LOGIC;
  SIGNAL or_1230_nl : STD_LOGIC;
  SIGNAL or_1229_nl : STD_LOGIC;
  SIGNAL mux_1148_nl : STD_LOGIC;
  SIGNAL or_1228_nl : STD_LOGIC;
  SIGNAL mux_1147_nl : STD_LOGIC;
  SIGNAL or_1227_nl : STD_LOGIC;
  SIGNAL mux_1207_nl : STD_LOGIC;
  SIGNAL mux_1206_nl : STD_LOGIC;
  SIGNAL nor_404_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL or_1320_nl : STD_LOGIC;
  SIGNAL mux_1203_nl : STD_LOGIC;
  SIGNAL or_1319_nl : STD_LOGIC;
  SIGNAL mux_1202_nl : STD_LOGIC;
  SIGNAL mux_1201_nl : STD_LOGIC;
  SIGNAL or_1316_nl : STD_LOGIC;
  SIGNAL or_1314_nl : STD_LOGIC;
  SIGNAL mux_1200_nl : STD_LOGIC;
  SIGNAL or_1313_nl : STD_LOGIC;
  SIGNAL or_1311_nl : STD_LOGIC;
  SIGNAL mux_1199_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL mux_1197_nl : STD_LOGIC;
  SIGNAL or_1309_nl : STD_LOGIC;
  SIGNAL or_1307_nl : STD_LOGIC;
  SIGNAL or_1306_nl : STD_LOGIC;
  SIGNAL nor_406_nl : STD_LOGIC;
  SIGNAL mux_1196_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL nor_407_nl : STD_LOGIC;
  SIGNAL and_311_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL nor_408_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL nor_409_nl : STD_LOGIC;
  SIGNAL nor_410_nl : STD_LOGIC;
  SIGNAL and_312_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL nor_411_nl : STD_LOGIC;
  SIGNAL nor_412_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL nor_414_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL nor_415_nl : STD_LOGIC;
  SIGNAL nor_416_nl : STD_LOGIC;
  SIGNAL nor_417_nl : STD_LOGIC;
  SIGNAL nor_418_nl : STD_LOGIC;
  SIGNAL mux_1186_nl : STD_LOGIC;
  SIGNAL nand_71_nl : STD_LOGIC;
  SIGNAL mux_1185_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL mux_1183_nl : STD_LOGIC;
  SIGNAL nor_420_nl : STD_LOGIC;
  SIGNAL mux_1182_nl : STD_LOGIC;
  SIGNAL nor_421_nl : STD_LOGIC;
  SIGNAL nor_422_nl : STD_LOGIC;
  SIGNAL nor_423_nl : STD_LOGIC;
  SIGNAL or_1277_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL or_1276_nl : STD_LOGIC;
  SIGNAL mux_1180_nl : STD_LOGIC;
  SIGNAL mux_1179_nl : STD_LOGIC;
  SIGNAL or_1274_nl : STD_LOGIC;
  SIGNAL or_1273_nl : STD_LOGIC;
  SIGNAL mux_1178_nl : STD_LOGIC;
  SIGNAL or_1270_nl : STD_LOGIC;
  SIGNAL mux_1238_nl : STD_LOGIC;
  SIGNAL mux_1237_nl : STD_LOGIC;
  SIGNAL nor_398_nl : STD_LOGIC;
  SIGNAL mux_1236_nl : STD_LOGIC;
  SIGNAL nand_76_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL or_1366_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL or_1365_nl : STD_LOGIC;
  SIGNAL or_1364_nl : STD_LOGIC;
  SIGNAL mux_1232_nl : STD_LOGIC;
  SIGNAL and_441_nl : STD_LOGIC;
  SIGNAL nor_400_nl : STD_LOGIC;
  SIGNAL mux_1231_nl : STD_LOGIC;
  SIGNAL or_1359_nl : STD_LOGIC;
  SIGNAL mux_1230_nl : STD_LOGIC;
  SIGNAL and_310_nl : STD_LOGIC;
  SIGNAL mux_1229_nl : STD_LOGIC;
  SIGNAL nand_378_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL mux_1226_nl : STD_LOGIC;
  SIGNAL or_1354_nl : STD_LOGIC;
  SIGNAL mux_1225_nl : STD_LOGIC;
  SIGNAL or_1352_nl : STD_LOGIC;
  SIGNAL or_1351_nl : STD_LOGIC;
  SIGNAL mux_1224_nl : STD_LOGIC;
  SIGNAL or_1350_nl : STD_LOGIC;
  SIGNAL nor_401_nl : STD_LOGIC;
  SIGNAL mux_1223_nl : STD_LOGIC;
  SIGNAL nor_402_nl : STD_LOGIC;
  SIGNAL mux_1222_nl : STD_LOGIC;
  SIGNAL mux_1221_nl : STD_LOGIC;
  SIGNAL nand_373_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL mux_1219_nl : STD_LOGIC;
  SIGNAL or_1344_nl : STD_LOGIC;
  SIGNAL mux_1218_nl : STD_LOGIC;
  SIGNAL or_1342_nl : STD_LOGIC;
  SIGNAL mux_1217_nl : STD_LOGIC;
  SIGNAL or_1341_nl : STD_LOGIC;
  SIGNAL mux_1216_nl : STD_LOGIC;
  SIGNAL or_1340_nl : STD_LOGIC;
  SIGNAL nor_403_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL nand_74_nl : STD_LOGIC;
  SIGNAL mux_1214_nl : STD_LOGIC;
  SIGNAL nand_363_nl : STD_LOGIC;
  SIGNAL mux_1213_nl : STD_LOGIC;
  SIGNAL mux_1212_nl : STD_LOGIC;
  SIGNAL or_1335_nl : STD_LOGIC;
  SIGNAL mux_1211_nl : STD_LOGIC;
  SIGNAL or_1329_nl : STD_LOGIC;
  SIGNAL or_1328_nl : STD_LOGIC;
  SIGNAL mux_1210_nl : STD_LOGIC;
  SIGNAL or_1327_nl : STD_LOGIC;
  SIGNAL mux_1209_nl : STD_LOGIC;
  SIGNAL or_1326_nl : STD_LOGIC;
  SIGNAL mux_1269_nl : STD_LOGIC;
  SIGNAL mux_1268_nl : STD_LOGIC;
  SIGNAL nor_379_nl : STD_LOGIC;
  SIGNAL mux_1267_nl : STD_LOGIC;
  SIGNAL mux_1266_nl : STD_LOGIC;
  SIGNAL nand_240_nl : STD_LOGIC;
  SIGNAL mux_1265_nl : STD_LOGIC;
  SIGNAL or_1418_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL or_1415_nl : STD_LOGIC;
  SIGNAL or_1413_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL nand_369_nl : STD_LOGIC;
  SIGNAL or_1410_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL nor_380_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL mux_1259_nl : STD_LOGIC;
  SIGNAL or_1408_nl : STD_LOGIC;
  SIGNAL or_1406_nl : STD_LOGIC;
  SIGNAL or_1405_nl : STD_LOGIC;
  SIGNAL nor_381_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL nor_382_nl : STD_LOGIC;
  SIGNAL and_307_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL nor_383_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL and_308_nl : STD_LOGIC;
  SIGNAL nor_384_nl : STD_LOGIC;
  SIGNAL and_309_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL nor_385_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL mux_1251_nl : STD_LOGIC;
  SIGNAL nor_388_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL nor_389_nl : STD_LOGIC;
  SIGNAL and_431_nl : STD_LOGIC;
  SIGNAL nor_391_nl : STD_LOGIC;
  SIGNAL nor_392_nl : STD_LOGIC;
  SIGNAL mux_1248_nl : STD_LOGIC;
  SIGNAL nand_77_nl : STD_LOGIC;
  SIGNAL mux_1247_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL mux_1245_nl : STD_LOGIC;
  SIGNAL nor_394_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL nor_395_nl : STD_LOGIC;
  SIGNAL nor_396_nl : STD_LOGIC;
  SIGNAL nor_397_nl : STD_LOGIC;
  SIGNAL or_1376_nl : STD_LOGIC;
  SIGNAL mux_1243_nl : STD_LOGIC;
  SIGNAL or_1375_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL nand_248_nl : STD_LOGIC;
  SIGNAL or_1372_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL nand_352_nl : STD_LOGIC;
  SIGNAL mux_1300_nl : STD_LOGIC;
  SIGNAL mux_1299_nl : STD_LOGIC;
  SIGNAL nor_373_nl : STD_LOGIC;
  SIGNAL mux_1298_nl : STD_LOGIC;
  SIGNAL nand_82_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL mux_1296_nl : STD_LOGIC;
  SIGNAL or_1465_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL or_1464_nl : STD_LOGIC;
  SIGNAL or_1463_nl : STD_LOGIC;
  SIGNAL mux_1294_nl : STD_LOGIC;
  SIGNAL and_436_nl : STD_LOGIC;
  SIGNAL nor_375_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL or_1458_nl : STD_LOGIC;
  SIGNAL mux_1292_nl : STD_LOGIC;
  SIGNAL and_306_nl : STD_LOGIC;
  SIGNAL mux_1291_nl : STD_LOGIC;
  SIGNAL or_1455_nl : STD_LOGIC;
  SIGNAL mux_1290_nl : STD_LOGIC;
  SIGNAL mux_1289_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL or_1453_nl : STD_LOGIC;
  SIGNAL mux_1287_nl : STD_LOGIC;
  SIGNAL or_1451_nl : STD_LOGIC;
  SIGNAL or_1450_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL or_1449_nl : STD_LOGIC;
  SIGNAL nor_376_nl : STD_LOGIC;
  SIGNAL mux_1285_nl : STD_LOGIC;
  SIGNAL nor_377_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL mux_1283_nl : STD_LOGIC;
  SIGNAL or_1445_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL mux_1281_nl : STD_LOGIC;
  SIGNAL or_1443_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL or_1441_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL or_1440_nl : STD_LOGIC;
  SIGNAL mux_1278_nl : STD_LOGIC;
  SIGNAL or_1439_nl : STD_LOGIC;
  SIGNAL nor_378_nl : STD_LOGIC;
  SIGNAL mux_1277_nl : STD_LOGIC;
  SIGNAL nand_80_nl : STD_LOGIC;
  SIGNAL mux_1276_nl : STD_LOGIC;
  SIGNAL or_1436_nl : STD_LOGIC;
  SIGNAL mux_1275_nl : STD_LOGIC;
  SIGNAL mux_1274_nl : STD_LOGIC;
  SIGNAL or_1434_nl : STD_LOGIC;
  SIGNAL mux_1273_nl : STD_LOGIC;
  SIGNAL or_1428_nl : STD_LOGIC;
  SIGNAL or_1427_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL or_1426_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL or_1425_nl : STD_LOGIC;
  SIGNAL mux_1331_nl : STD_LOGIC;
  SIGNAL mux_1330_nl : STD_LOGIC;
  SIGNAL nor_353_nl : STD_LOGIC;
  SIGNAL mux_1329_nl : STD_LOGIC;
  SIGNAL mux_1328_nl : STD_LOGIC;
  SIGNAL or_1518_nl : STD_LOGIC;
  SIGNAL mux_1327_nl : STD_LOGIC;
  SIGNAL or_1517_nl : STD_LOGIC;
  SIGNAL mux_1326_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL or_1514_nl : STD_LOGIC;
  SIGNAL or_1512_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL or_1511_nl : STD_LOGIC;
  SIGNAL or_1509_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL nor_354_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL or_1507_nl : STD_LOGIC;
  SIGNAL or_1505_nl : STD_LOGIC;
  SIGNAL or_1504_nl : STD_LOGIC;
  SIGNAL nor_355_nl : STD_LOGIC;
  SIGNAL mux_1320_nl : STD_LOGIC;
  SIGNAL mux_1319_nl : STD_LOGIC;
  SIGNAL nor_356_nl : STD_LOGIC;
  SIGNAL and_304_nl : STD_LOGIC;
  SIGNAL mux_1318_nl : STD_LOGIC;
  SIGNAL nor_357_nl : STD_LOGIC;
  SIGNAL mux_1317_nl : STD_LOGIC;
  SIGNAL nor_358_nl : STD_LOGIC;
  SIGNAL nor_359_nl : STD_LOGIC;
  SIGNAL and_305_nl : STD_LOGIC;
  SIGNAL mux_1316_nl : STD_LOGIC;
  SIGNAL mux_1315_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL nor_360_nl : STD_LOGIC;
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL nor_363_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL nor_364_nl : STD_LOGIC;
  SIGNAL nor_365_nl : STD_LOGIC;
  SIGNAL nor_366_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL nand_83_nl : STD_LOGIC;
  SIGNAL mux_1309_nl : STD_LOGIC;
  SIGNAL mux_1308_nl : STD_LOGIC;
  SIGNAL mux_1307_nl : STD_LOGIC;
  SIGNAL nor_369_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL nor_370_nl : STD_LOGIC;
  SIGNAL nor_371_nl : STD_LOGIC;
  SIGNAL nor_372_nl : STD_LOGIC;
  SIGNAL or_1475_nl : STD_LOGIC;
  SIGNAL mux_1305_nl : STD_LOGIC;
  SIGNAL or_1474_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL mux_1303_nl : STD_LOGIC;
  SIGNAL or_1472_nl : STD_LOGIC;
  SIGNAL or_1471_nl : STD_LOGIC;
  SIGNAL mux_1302_nl : STD_LOGIC;
  SIGNAL or_1468_nl : STD_LOGIC;
  SIGNAL mux_1362_nl : STD_LOGIC;
  SIGNAL mux_1361_nl : STD_LOGIC;
  SIGNAL mux_1360_nl : STD_LOGIC;
  SIGNAL nor_346_nl : STD_LOGIC;
  SIGNAL mux_1359_nl : STD_LOGIC;
  SIGNAL mux_1358_nl : STD_LOGIC;
  SIGNAL or_1565_nl : STD_LOGIC;
  SIGNAL mux_1357_nl : STD_LOGIC;
  SIGNAL or_1564_nl : STD_LOGIC;
  SIGNAL and_302_nl : STD_LOGIC;
  SIGNAL mux_1356_nl : STD_LOGIC;
  SIGNAL nand_230_nl : STD_LOGIC;
  SIGNAL mux_1355_nl : STD_LOGIC;
  SIGNAL mux_1354_nl : STD_LOGIC;
  SIGNAL or_1561_nl : STD_LOGIC;
  SIGNAL mux_1353_nl : STD_LOGIC;
  SIGNAL or_1560_nl : STD_LOGIC;
  SIGNAL nor_347_nl : STD_LOGIC;
  SIGNAL mux_1352_nl : STD_LOGIC;
  SIGNAL or_1557_nl : STD_LOGIC;
  SIGNAL nor_348_nl : STD_LOGIC;
  SIGNAL mux_1351_nl : STD_LOGIC;
  SIGNAL mux_1350_nl : STD_LOGIC;
  SIGNAL or_1554_nl : STD_LOGIC;
  SIGNAL nand_231_nl : STD_LOGIC;
  SIGNAL nand_86_nl : STD_LOGIC;
  SIGNAL mux_1349_nl : STD_LOGIC;
  SIGNAL or_1551_nl : STD_LOGIC;
  SIGNAL mux_1348_nl : STD_LOGIC;
  SIGNAL or_1550_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL nor_349_nl : STD_LOGIC;
  SIGNAL mux_1345_nl : STD_LOGIC;
  SIGNAL and_303_nl : STD_LOGIC;
  SIGNAL nor_350_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL or_1544_nl : STD_LOGIC;
  SIGNAL mux_1343_nl : STD_LOGIC;
  SIGNAL or_1543_nl : STD_LOGIC;
  SIGNAL mux_1342_nl : STD_LOGIC;
  SIGNAL nor_351_nl : STD_LOGIC;
  SIGNAL mux_1341_nl : STD_LOGIC;
  SIGNAL nand_232_nl : STD_LOGIC;
  SIGNAL mux_1340_nl : STD_LOGIC;
  SIGNAL mux_1339_nl : STD_LOGIC;
  SIGNAL or_1537_nl : STD_LOGIC;
  SIGNAL mux_1338_nl : STD_LOGIC;
  SIGNAL or_1536_nl : STD_LOGIC;
  SIGNAL nor_352_nl : STD_LOGIC;
  SIGNAL mux_1337_nl : STD_LOGIC;
  SIGNAL mux_1336_nl : STD_LOGIC;
  SIGNAL mux_1335_nl : STD_LOGIC;
  SIGNAL or_1532_nl : STD_LOGIC;
  SIGNAL mux_1334_nl : STD_LOGIC;
  SIGNAL or_1527_nl : STD_LOGIC;
  SIGNAL or_1525_nl : STD_LOGIC;
  SIGNAL mux_1333_nl : STD_LOGIC;
  SIGNAL or_1524_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL nor_327_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL nand_216_nl : STD_LOGIC;
  SIGNAL mux_1389_nl : STD_LOGIC;
  SIGNAL or_1615_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL mux_1387_nl : STD_LOGIC;
  SIGNAL or_1612_nl : STD_LOGIC;
  SIGNAL or_1611_nl : STD_LOGIC;
  SIGNAL mux_1386_nl : STD_LOGIC;
  SIGNAL nand_368_nl : STD_LOGIC;
  SIGNAL or_1608_nl : STD_LOGIC;
  SIGNAL mux_1385_nl : STD_LOGIC;
  SIGNAL nor_328_nl : STD_LOGIC;
  SIGNAL mux_1384_nl : STD_LOGIC;
  SIGNAL mux_1383_nl : STD_LOGIC;
  SIGNAL or_1606_nl : STD_LOGIC;
  SIGNAL or_1604_nl : STD_LOGIC;
  SIGNAL or_1603_nl : STD_LOGIC;
  SIGNAL nor_329_nl : STD_LOGIC;
  SIGNAL mux_1382_nl : STD_LOGIC;
  SIGNAL mux_1381_nl : STD_LOGIC;
  SIGNAL nor_330_nl : STD_LOGIC;
  SIGNAL and_299_nl : STD_LOGIC;
  SIGNAL mux_1380_nl : STD_LOGIC;
  SIGNAL nor_331_nl : STD_LOGIC;
  SIGNAL mux_1379_nl : STD_LOGIC;
  SIGNAL and_300_nl : STD_LOGIC;
  SIGNAL nor_332_nl : STD_LOGIC;
  SIGNAL and_301_nl : STD_LOGIC;
  SIGNAL mux_1378_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL mux_1376_nl : STD_LOGIC;
  SIGNAL nor_333_nl : STD_LOGIC;
  SIGNAL nor_334_nl : STD_LOGIC;
  SIGNAL mux_1375_nl : STD_LOGIC;
  SIGNAL nor_336_nl : STD_LOGIC;
  SIGNAL mux_1374_nl : STD_LOGIC;
  SIGNAL mux_1373_nl : STD_LOGIC;
  SIGNAL nor_337_nl : STD_LOGIC;
  SIGNAL and_430_nl : STD_LOGIC;
  SIGNAL nor_339_nl : STD_LOGIC;
  SIGNAL nor_340_nl : STD_LOGIC;
  SIGNAL mux_1372_nl : STD_LOGIC;
  SIGNAL nand_89_nl : STD_LOGIC;
  SIGNAL mux_1371_nl : STD_LOGIC;
  SIGNAL mux_1370_nl : STD_LOGIC;
  SIGNAL mux_1369_nl : STD_LOGIC;
  SIGNAL nor_342_nl : STD_LOGIC;
  SIGNAL mux_1368_nl : STD_LOGIC;
  SIGNAL nor_343_nl : STD_LOGIC;
  SIGNAL nor_344_nl : STD_LOGIC;
  SIGNAL nor_345_nl : STD_LOGIC;
  SIGNAL or_1574_nl : STD_LOGIC;
  SIGNAL mux_1367_nl : STD_LOGIC;
  SIGNAL or_1573_nl : STD_LOGIC;
  SIGNAL mux_1366_nl : STD_LOGIC;
  SIGNAL mux_1365_nl : STD_LOGIC;
  SIGNAL nand_224_nl : STD_LOGIC;
  SIGNAL or_1570_nl : STD_LOGIC;
  SIGNAL mux_1364_nl : STD_LOGIC;
  SIGNAL nand_351_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL nor_321_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL nand_94_nl : STD_LOGIC;
  SIGNAL mux_1421_nl : STD_LOGIC;
  SIGNAL mux_1420_nl : STD_LOGIC;
  SIGNAL or_1662_nl : STD_LOGIC;
  SIGNAL mux_1419_nl : STD_LOGIC;
  SIGNAL or_1661_nl : STD_LOGIC;
  SIGNAL or_1660_nl : STD_LOGIC;
  SIGNAL mux_1418_nl : STD_LOGIC;
  SIGNAL and_435_nl : STD_LOGIC;
  SIGNAL nor_323_nl : STD_LOGIC;
  SIGNAL mux_1417_nl : STD_LOGIC;
  SIGNAL or_1655_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL and_298_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL nand_375_nl : STD_LOGIC;
  SIGNAL mux_1414_nl : STD_LOGIC;
  SIGNAL mux_1413_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL or_1650_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL or_1648_nl : STD_LOGIC;
  SIGNAL or_1647_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL or_1646_nl : STD_LOGIC;
  SIGNAL nor_324_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL nor_325_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL nand_367_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL or_1640_nl : STD_LOGIC;
  SIGNAL mux_1404_nl : STD_LOGIC;
  SIGNAL or_1638_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL or_1637_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL or_1636_nl : STD_LOGIC;
  SIGNAL nor_326_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL nand_92_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL nand_359_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL or_1631_nl : STD_LOGIC;
  SIGNAL mux_1397_nl : STD_LOGIC;
  SIGNAL or_1625_nl : STD_LOGIC;
  SIGNAL or_1624_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL or_1623_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL or_1622_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL mux_1454_nl : STD_LOGIC;
  SIGNAL nor_302_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL nand_196_nl : STD_LOGIC;
  SIGNAL mux_1451_nl : STD_LOGIC;
  SIGNAL or_1712_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL or_1709_nl : STD_LOGIC;
  SIGNAL or_1707_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL nand_366_nl : STD_LOGIC;
  SIGNAL or_1704_nl : STD_LOGIC;
  SIGNAL mux_1447_nl : STD_LOGIC;
  SIGNAL nor_303_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL or_1702_nl : STD_LOGIC;
  SIGNAL or_1700_nl : STD_LOGIC;
  SIGNAL or_1699_nl : STD_LOGIC;
  SIGNAL nor_304_nl : STD_LOGIC;
  SIGNAL mux_1444_nl : STD_LOGIC;
  SIGNAL mux_1443_nl : STD_LOGIC;
  SIGNAL nor_305_nl : STD_LOGIC;
  SIGNAL and_295_nl : STD_LOGIC;
  SIGNAL mux_1442_nl : STD_LOGIC;
  SIGNAL nor_306_nl : STD_LOGIC;
  SIGNAL mux_1441_nl : STD_LOGIC;
  SIGNAL and_296_nl : STD_LOGIC;
  SIGNAL nor_307_nl : STD_LOGIC;
  SIGNAL and_297_nl : STD_LOGIC;
  SIGNAL mux_1440_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL nor_308_nl : STD_LOGIC;
  SIGNAL nor_309_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL nor_311_nl : STD_LOGIC;
  SIGNAL mux_1436_nl : STD_LOGIC;
  SIGNAL mux_1435_nl : STD_LOGIC;
  SIGNAL nor_312_nl : STD_LOGIC;
  SIGNAL and_429_nl : STD_LOGIC;
  SIGNAL nor_314_nl : STD_LOGIC;
  SIGNAL nor_315_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL nand_95_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL nor_317_nl : STD_LOGIC;
  SIGNAL mux_1430_nl : STD_LOGIC;
  SIGNAL nor_318_nl : STD_LOGIC;
  SIGNAL nor_319_nl : STD_LOGIC;
  SIGNAL nor_320_nl : STD_LOGIC;
  SIGNAL or_1671_nl : STD_LOGIC;
  SIGNAL mux_1429_nl : STD_LOGIC;
  SIGNAL or_1670_nl : STD_LOGIC;
  SIGNAL mux_1428_nl : STD_LOGIC;
  SIGNAL mux_1427_nl : STD_LOGIC;
  SIGNAL nand_204_nl : STD_LOGIC;
  SIGNAL or_1667_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL nand_350_nl : STD_LOGIC;
  SIGNAL mux_1486_nl : STD_LOGIC;
  SIGNAL mux_1485_nl : STD_LOGIC;
  SIGNAL nor_296_nl : STD_LOGIC;
  SIGNAL mux_1484_nl : STD_LOGIC;
  SIGNAL nand_100_nl : STD_LOGIC;
  SIGNAL mux_1483_nl : STD_LOGIC;
  SIGNAL mux_1482_nl : STD_LOGIC;
  SIGNAL or_1756_nl : STD_LOGIC;
  SIGNAL mux_1481_nl : STD_LOGIC;
  SIGNAL nand_178_nl : STD_LOGIC;
  SIGNAL or_1754_nl : STD_LOGIC;
  SIGNAL mux_1480_nl : STD_LOGIC;
  SIGNAL and_434_nl : STD_LOGIC;
  SIGNAL nor_298_nl : STD_LOGIC;
  SIGNAL mux_1479_nl : STD_LOGIC;
  SIGNAL nand_377_nl : STD_LOGIC;
  SIGNAL mux_1478_nl : STD_LOGIC;
  SIGNAL and_294_nl : STD_LOGIC;
  SIGNAL mux_1477_nl : STD_LOGIC;
  SIGNAL nand_374_nl : STD_LOGIC;
  SIGNAL mux_1476_nl : STD_LOGIC;
  SIGNAL mux_1475_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL nand_372_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL nand_183_nl : STD_LOGIC;
  SIGNAL or_1741_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL nand_184_nl : STD_LOGIC;
  SIGNAL nor_299_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL nor_300_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL mux_1469_nl : STD_LOGIC;
  SIGNAL nand_365_nl : STD_LOGIC;
  SIGNAL mux_1468_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL nand_362_nl : STD_LOGIC;
  SIGNAL mux_1466_nl : STD_LOGIC;
  SIGNAL nand_187_nl : STD_LOGIC;
  SIGNAL mux_1465_nl : STD_LOGIC;
  SIGNAL or_1731_nl : STD_LOGIC;
  SIGNAL mux_1464_nl : STD_LOGIC;
  SIGNAL nand_188_nl : STD_LOGIC;
  SIGNAL nor_301_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL nand_98_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL nand_358_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL mux_1460_nl : STD_LOGIC;
  SIGNAL nand_349_nl : STD_LOGIC;
  SIGNAL mux_1459_nl : STD_LOGIC;
  SIGNAL nand_191_nl : STD_LOGIC;
  SIGNAL or_1721_nl : STD_LOGIC;
  SIGNAL mux_1458_nl : STD_LOGIC;
  SIGNAL or_1720_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL nand_192_nl : STD_LOGIC;
  SIGNAL mux_1517_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL nor_282_nl : STD_LOGIC;
  SIGNAL mux_1515_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL nand_158_nl : STD_LOGIC;
  SIGNAL mux_1513_nl : STD_LOGIC;
  SIGNAL or_1802_nl : STD_LOGIC;
  SIGNAL mux_1512_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL nand_162_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL nand_364_nl : STD_LOGIC;
  SIGNAL or_1796_nl : STD_LOGIC;
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL nor_283_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL nand_361_nl : STD_LOGIC;
  SIGNAL nand_164_nl : STD_LOGIC;
  SIGNAL or_1791_nl : STD_LOGIC;
  SIGNAL nor_284_nl : STD_LOGIC;
  SIGNAL mux_1506_nl : STD_LOGIC;
  SIGNAL mux_1505_nl : STD_LOGIC;
  SIGNAL nor_285_nl : STD_LOGIC;
  SIGNAL and_286_nl : STD_LOGIC;
  SIGNAL mux_1504_nl : STD_LOGIC;
  SIGNAL nor_286_nl : STD_LOGIC;
  SIGNAL mux_1503_nl : STD_LOGIC;
  SIGNAL and_287_nl : STD_LOGIC;
  SIGNAL and_288_nl : STD_LOGIC;
  SIGNAL and_289_nl : STD_LOGIC;
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL mux_1500_nl : STD_LOGIC;
  SIGNAL and_290_nl : STD_LOGIC;
  SIGNAL nor_287_nl : STD_LOGIC;
  SIGNAL mux_1499_nl : STD_LOGIC;
  SIGNAL and_427_nl : STD_LOGIC;
  SIGNAL mux_1498_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL and_292_nl : STD_LOGIC;
  SIGNAL and_428_nl : STD_LOGIC;
  SIGNAL nor_290_nl : STD_LOGIC;
  SIGNAL nor_291_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL nand_101_nl : STD_LOGIC;
  SIGNAL mux_1495_nl : STD_LOGIC;
  SIGNAL mux_1494_nl : STD_LOGIC;
  SIGNAL mux_1493_nl : STD_LOGIC;
  SIGNAL and_433_nl : STD_LOGIC;
  SIGNAL mux_1492_nl : STD_LOGIC;
  SIGNAL nor_293_nl : STD_LOGIC;
  SIGNAL and_440_nl : STD_LOGIC;
  SIGNAL nor_295_nl : STD_LOGIC;
  SIGNAL or_1764_nl : STD_LOGIC;
  SIGNAL mux_1491_nl : STD_LOGIC;
  SIGNAL or_1763_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL mux_1489_nl : STD_LOGIC;
  SIGNAL nand_172_nl : STD_LOGIC;
  SIGNAL mux_1488_nl : STD_LOGIC;
  SIGNAL nand_348_nl : STD_LOGIC;
  SIGNAL or_2213_nl : STD_LOGIC;
  SIGNAL mux_2057_nl : STD_LOGIC;
  SIGNAL mux_2065_nl : STD_LOGIC;
  SIGNAL mux_2064_nl : STD_LOGIC;
  SIGNAL or_2219_nl : STD_LOGIC;
  SIGNAL mux_2063_nl : STD_LOGIC;
  SIGNAL or_2218_nl : STD_LOGIC;
  SIGNAL mux_2062_nl : STD_LOGIC;
  SIGNAL mux_2061_nl : STD_LOGIC;
  SIGNAL or_2214_nl : STD_LOGIC;
  SIGNAL mux_2060_nl : STD_LOGIC;
  SIGNAL mux_2059_nl : STD_LOGIC;
  SIGNAL or_2209_nl : STD_LOGIC;
  SIGNAL or_2208_nl : STD_LOGIC;
  SIGNAL mux_2056_nl : STD_LOGIC;
  SIGNAL or_2207_nl : STD_LOGIC;
  SIGNAL mux_2055_nl : STD_LOGIC;
  SIGNAL or_2261_nl : STD_LOGIC;
  SIGNAL or_2267_nl : STD_LOGIC;
  SIGNAL or_2266_nl : STD_LOGIC;
  SIGNAL mux_2097_nl : STD_LOGIC;
  SIGNAL or_2271_nl : STD_LOGIC;
  SIGNAL or_2270_nl : STD_LOGIC;
  SIGNAL nand_388_nl : STD_LOGIC;
  SIGNAL mux_2103_nl : STD_LOGIC;
  SIGNAL nand_389_nl : STD_LOGIC;
  SIGNAL mux_2102_nl : STD_LOGIC;
  SIGNAL mux_2101_nl : STD_LOGIC;
  SIGNAL or_2272_nl : STD_LOGIC;
  SIGNAL or_2282_nl : STD_LOGIC;
  SIGNAL mux_2123_nl : STD_LOGIC;
  SIGNAL or_2302_nl : STD_LOGIC;
  SIGNAL mux_2134_nl : STD_LOGIC;
  SIGNAL mux_2132_nl : STD_LOGIC;
  SIGNAL mux_2131_nl : STD_LOGIC;
  SIGNAL mux_2163_nl : STD_LOGIC;
  SIGNAL mux_2170_nl : STD_LOGIC;
  SIGNAL mux_2169_nl : STD_LOGIC;
  SIGNAL mux_2167_nl : STD_LOGIC;
  SIGNAL mux_2166_nl : STD_LOGIC;
  SIGNAL mux_2175_nl : STD_LOGIC;
  SIGNAL mux_2179_nl : STD_LOGIC;
  SIGNAL or_2346_nl : STD_LOGIC;
  SIGNAL mux_2215_nl : STD_LOGIC;
  SIGNAL mux_2220_nl : STD_LOGIC;
  SIGNAL or_2350_nl : STD_LOGIC;
  SIGNAL nand_399_nl : STD_LOGIC;
  SIGNAL or_2360_nl : STD_LOGIC;
  SIGNAL acc_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_3_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_15_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_or_52_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_53_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_mux1h_271_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_or_54_nl : STD_LOGIC;
  SIGNAL acc_1_nl : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_or_4_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_mux_16_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_or_55_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_or_56_nl : STD_LOGIC;
  SIGNAL COMP_LOOP_COMP_LOOP_or_5_nl : STD_LOGIC;
  SIGNAL operator_64_false_1_mux_1_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL acc_3_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_35_nl : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nand_1_nl : STD_LOGIC;
  SIGNAL acc_4_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL COMP_LOOP_mux_36_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL COMP_LOOP_or_57_nl : STD_LOGIC;
  SIGNAL acc_5_nl : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL COMP_LOOP_or_58_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_COMP_LOOP_nor_63_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL COMP_LOOP_mux1h_272_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_706_nl : STD_LOGIC;
  SIGNAL and_707_nl : STD_LOGIC;
  SIGNAL and_708_nl : STD_LOGIC;
  SIGNAL and_709_nl : STD_LOGIC;
  SIGNAL and_710_nl : STD_LOGIC;
  SIGNAL and_711_nl : STD_LOGIC;
  SIGNAL and_712_nl : STD_LOGIC;
  SIGNAL and_713_nl : STD_LOGIC;
  SIGNAL and_714_nl : STD_LOGIC;
  SIGNAL and_715_nl : STD_LOGIC;
  SIGNAL and_716_nl : STD_LOGIC;
  SIGNAL and_717_nl : STD_LOGIC;
  SIGNAL and_718_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_STAGE_LOOP_or_1_nl : STD_LOGIC;
  SIGNAL STAGE_LOOP_STAGE_LOOP_mux_2_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL STAGE_LOOP_or_2_nl : STD_LOGIC;
  SIGNAL operator_64_false_acc_nl : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_64_false_operator_64_false_operator_64_false_nor_1_nl : STD_LOGIC_VECTOR
      (60 DOWNTO 0);
  SIGNAL operator_64_false_mux_1_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_64_false_mux1h_1_nl : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL and_719_nl : STD_LOGIC;
  SIGNAL and_720_nl : STD_LOGIC;
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL r_rsci_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL r_rsci_idat_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);

  COMPONENT modulo_dev
    PORT (
      base_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      m_rsc_dat : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      return_rsc_z : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      ccs_ccore_start_rsc_dat : IN STD_LOGIC;
      ccs_ccore_clk : IN STD_LOGIC;
      ccs_ccore_srst : IN STD_LOGIC;
      ccs_ccore_en : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL modulo_dev_cmp_base_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_cmp_m_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_cmp_return_rsc_z_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL modulo_dev_cmp_ccs_ccore_start_rsc_dat : STD_LOGIC;

  SIGNAL operator_66_true_div_cmp_a_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_b : STD_LOGIC_VECTOR (10 DOWNTO 0);
  SIGNAL operator_66_true_div_cmp_z_1 : STD_LOGIC_VECTOR (64 DOWNTO 0);

  SIGNAL STAGE_LOOP_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL STAGE_LOOP_lshift_rg_z : STD_LOGIC_VECTOR (9 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_core_wait_dp
    PORT(
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      modulo_dev_cmp_ccs_ccore_en : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_wait_dp_inst_ensig_cgo_iro : STD_LOGIC;

  COMPONENT inPlaceNTT_DIT_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      STAGE_LOOP_C_3_tr0 : IN STD_LOGIC;
      modExp_dev_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_1_tr0 : IN STD_LOGIC;
      COMP_LOOP_1_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_32_tr0 : IN STD_LOGIC;
      COMP_LOOP_2_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_64_tr0 : IN STD_LOGIC;
      COMP_LOOP_3_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_96_tr0 : IN STD_LOGIC;
      COMP_LOOP_4_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_128_tr0 : IN STD_LOGIC;
      COMP_LOOP_5_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_160_tr0 : IN STD_LOGIC;
      COMP_LOOP_6_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_192_tr0 : IN STD_LOGIC;
      COMP_LOOP_7_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_224_tr0 : IN STD_LOGIC;
      COMP_LOOP_8_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_256_tr0 : IN STD_LOGIC;
      COMP_LOOP_9_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_288_tr0 : IN STD_LOGIC;
      COMP_LOOP_10_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_320_tr0 : IN STD_LOGIC;
      COMP_LOOP_11_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_352_tr0 : IN STD_LOGIC;
      COMP_LOOP_12_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_384_tr0 : IN STD_LOGIC;
      COMP_LOOP_13_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_416_tr0 : IN STD_LOGIC;
      COMP_LOOP_14_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_448_tr0 : IN STD_LOGIC;
      COMP_LOOP_15_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_480_tr0 : IN STD_LOGIC;
      COMP_LOOP_16_modExp_dev_1_while_C_14_tr0 : IN STD_LOGIC;
      COMP_LOOP_C_512_tr0 : IN STD_LOGIC;
      VEC_LOOP_C_0_tr0 : IN STD_LOGIC;
      STAGE_LOOP_C_4_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (9 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_3_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_32_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_96_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_160_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_224_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_288_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_352_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_416_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_480_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_4_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_11_2(input_10 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_14_2(input_13 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(13 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_16_2(input_15 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_16_2(input_15 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(15 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_3_2(input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_64_4_2(input_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_17_2(input_16 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(16 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_55_2_2(input_0 : STD_LOGIC_VECTOR(54 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(54 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(54 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_61_2_2(input_0 : STD_LOGIC_VECTOR(60 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(60 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(60 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_64_2_2(input_0 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(63 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_65_2_2(input_0 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(64 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(64 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_6_2_2(input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_9_2_2(input_0 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(8 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 5,
      width => 64
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  r_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 6,
      width => 64
      )
    PORT MAP(
      dat => r_rsci_dat,
      idat => r_rsci_idat_1
    );
  r_rsci_dat <= r_rsc_dat;
  r_rsci_idat <= r_rsci_idat_1;

  vec_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_15_lz
    );
  vec_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_14_lz
    );
  vec_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_13_lz
    );
  vec_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_12_lz
    );
  vec_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_11_lz
    );
  vec_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_10_lz
    );
  vec_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_9_lz
    );
  vec_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_8_lz
    );
  vec_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_7_lz
    );
  vec_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_6_lz
    );
  vec_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_5_lz
    );
  vec_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_4_lz
    );
  vec_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_3_lz
    );
  vec_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_2_lz
    );
  vec_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_1_lz
    );
  vec_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => vec_rsc_triosy_0_0_lz
    );
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => p_rsc_triosy_lz
    );
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_vec_rsc_triosy_0_15_obj_ld_cse,
      lz => r_rsc_triosy_lz
    );
  modulo_dev_cmp : modulo_dev
    PORT MAP(
      base_rsc_dat => modulo_dev_cmp_base_rsc_dat,
      m_rsc_dat => modulo_dev_cmp_m_rsc_dat,
      return_rsc_z => modulo_dev_cmp_return_rsc_z_1,
      ccs_ccore_start_rsc_dat => modulo_dev_cmp_ccs_ccore_start_rsc_dat,
      ccs_ccore_clk => clk,
      ccs_ccore_srst => rst,
      ccs_ccore_en => modulo_dev_cmp_ccs_ccore_en
    );
  modulo_dev_cmp_base_rsc_dat <= MUX1HOT_v_64_3_2(operator_64_false_acc_mut_63_0,
      COMP_LOOP_1_mul_itm, STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_4_dfm)
      + SIGNED(modulo_dev_cmp_return_rsc_z), 64)), STD_LOGIC_VECTOR'( (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(((fsm_output(4))
      AND (NOT (MUX_s_1_2_2(or_tmp_1799, (MUX_s_1_2_2(or_tmp_1794, or_tmp_1793, fsm_output(6))),
      fsm_output(2))))), (NOT((fsm_output(4)) OR (MUX_s_1_2_2(or_2306_cse, (MUX_s_1_2_2(or_tmp_1788,
      or_tmp_1796, fsm_output(6))), fsm_output(2))))), fsm_output(5))), (MUX_s_1_2_2((NOT((fsm_output(4))
      OR mux_tmp_1537)), ((fsm_output(4)) AND (NOT mux_tmp_1534)), fsm_output(5))),
      fsm_output(1))), (MUX_s_1_2_2(((fsm_output(5)) AND (NOT (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_1799,
      or_tmp_1794, fsm_output(6))), or_tmp_1793, fsm_output(2))), mux_tmp_1537, fsm_output(4))))),
      (NOT((fsm_output(5)) OR (MUX_s_1_2_2(mux_tmp_1534, (MUX_s_1_2_2(or_tmp_1788,
      ((fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR
      (fsm_output(8))), fsm_output(2))), fsm_output(4))))), fsm_output(1))), fsm_output(0)))
      & ((and_dcpl_35 AND and_dcpl_122) OR (and_dcpl_30 AND and_dcpl_65) OR (and_dcpl_51
      AND and_dcpl_28) OR (and_dcpl_57 AND and_dcpl_28) OR (and_dcpl_55 AND and_dcpl_39)
      OR (and_dcpl_30 AND and_dcpl_91) OR (and_dcpl_40 AND and_dcpl_130) OR (and_dcpl_45
      AND and_dcpl_130) OR (and_dcpl_89 AND and_dcpl_73) OR (and_dcpl_87 AND and_dcpl_83)
      OR (and_dcpl_68 AND and_dcpl_79) OR (and_dcpl_75 AND and_dcpl_136) OR (and_dcpl_81
      AND and_dcpl_138) OR (and_dcpl_87 AND and_dcpl_101) OR (and_dcpl_68 AND and_dcpl_99)
      OR (and_dcpl_95 AND and_dcpl_103)) & not_tmp_370));
  modulo_dev_cmp_m_rsc_dat <= p_sva;
  modulo_dev_cmp_return_rsc_z <= modulo_dev_cmp_return_rsc_z_1;
  modulo_dev_cmp_ccs_ccore_start_rsc_dat <= NOT (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(mux_tmp_1563,
      ((NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (fsm_output(5)) OR (fsm_output(9))
      OR (fsm_output(8))), fsm_output(7))), (MUX_s_1_2_2(mux_tmp_1562, (MUX_s_1_2_2(or_tmp_1835,
      or_tmp_1825, fsm_output(1))), fsm_output(7))), fsm_output(4))), (MUX_s_1_2_2(mux_tmp_1566,
      (MUX_s_1_2_2((NOT((fsm_output(1)) AND (fsm_output(5)) AND (fsm_output(9)) AND
      (NOT (fsm_output(8))))), ((fsm_output(1)) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR (fsm_output(8))), fsm_output(7))), fsm_output(4))), fsm_output(3))), (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(mux_tmp_1579,
      (MUX_s_1_2_2(or_tmp_1841, or_tmp_1827, fsm_output(1))), fsm_output(7))), (MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_1841,
      or_tmp_1838, fsm_output(1))), (MUX_s_1_2_2(or_tmp_1841, or_tmp_1824, fsm_output(1))),
      fsm_output(7))), fsm_output(4))), (MUX_s_1_2_2((MUX_s_1_2_2(mux_tmp_1573, (MUX_s_1_2_2(or_tmp_1840,
      or_tmp_1830, fsm_output(1))), fsm_output(7))), (MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_1823,
      or_tmp_1818, fsm_output(1))), (MUX_s_1_2_2(or_tmp_1830, or_tmp_1840, fsm_output(1))),
      fsm_output(7))), fsm_output(4))), fsm_output(3))), fsm_output(2))), (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_1830,
      or_tmp_1835, fsm_output(1))), (MUX_s_1_2_2(or_tmp_1838, or_tmp_1835, fsm_output(1))),
      fsm_output(7))), (MUX_s_1_2_2(((fsm_output(1)) OR (fsm_output(6)) OR (NOT (fsm_output(5)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8)))), mux_tmp_1579, fsm_output(7))),
      fsm_output(4))), (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_1824, ((fsm_output(5))
      OR (NOT (fsm_output(9))) OR (fsm_output(8))), fsm_output(1))), ((fsm_output(1))
      OR (fsm_output(6)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(9))) OR (fsm_output(8))),
      fsm_output(7))), (MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_1831, or_tmp_1827, fsm_output(1))),
      mux_tmp_1573, fsm_output(7))), fsm_output(4))), fsm_output(3))), (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(((NOT
      (fsm_output(1))) OR (fsm_output(6)) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (fsm_output(8))), (MUX_s_1_2_2(or_tmp_1825, or_tmp_1827, fsm_output(1))),
      fsm_output(7))), (MUX_s_1_2_2((MUX_s_1_2_2(((NOT (fsm_output(5))) OR (fsm_output(9))
      OR (fsm_output(8))), or_tmp_1825, fsm_output(1))), mux_tmp_1566, fsm_output(7))),
      fsm_output(4))), (MUX_s_1_2_2((MUX_s_1_2_2(((NOT (fsm_output(1))) OR (NOT (fsm_output(6)))
      OR (fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(8)))), mux_tmp_1563,
      fsm_output(7))), mux_tmp_1562, fsm_output(4))), fsm_output(3))), fsm_output(2))),
      fsm_output(0)));

  operator_66_true_div_cmp : work.mgc_comps.mgc_div
    GENERIC MAP(
      width_a => 65,
      width_b => 11,
      signd => 1
      )
    PORT MAP(
      a => operator_66_true_div_cmp_a_1,
      b => operator_66_true_div_cmp_b,
      z => operator_66_true_div_cmp_z_1
    );
  operator_66_true_div_cmp_a_1 <= operator_66_true_div_cmp_a;
  operator_66_true_div_cmp_b <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(operator_66_true_div_cmp_b_9_0));
  operator_66_true_div_cmp_z <= operator_66_true_div_cmp_z_1;

  STAGE_LOOP_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 0,
      width_s => 4,
      width_z => 10
      )
    PORT MAP(
      a => STAGE_LOOP_lshift_rg_a,
      s => STAGE_LOOP_lshift_rg_s,
      z => STAGE_LOOP_lshift_rg_z
    );
  STAGE_LOOP_lshift_rg_a(0) <= '1';
  STAGE_LOOP_lshift_rg_s <= STAGE_LOOP_i_3_0_sva;
  STAGE_LOOP_lshift_psp_sva_mx0w0 <= STAGE_LOOP_lshift_rg_z;

  inPlaceNTT_DIT_core_wait_dp_inst : inPlaceNTT_DIT_core_wait_dp
    PORT MAP(
      ensig_cgo_iro => inPlaceNTT_DIT_core_wait_dp_inst_ensig_cgo_iro,
      ensig_cgo => reg_ensig_cgo_cse,
      modulo_dev_cmp_ccs_ccore_en => modulo_dev_cmp_ccs_ccore_en
    );
  inPlaceNTT_DIT_core_wait_dp_inst_ensig_cgo_iro <= NOT mux_1581_itm;

  inPlaceNTT_DIT_core_core_fsm_inst : inPlaceNTT_DIT_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => inPlaceNTT_DIT_core_core_fsm_inst_fsm_output,
      STAGE_LOOP_C_3_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_3_tr0,
      modExp_dev_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_1_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_32_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_32_tr0,
      COMP_LOOP_2_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_64_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0,
      COMP_LOOP_3_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_96_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_96_tr0,
      COMP_LOOP_4_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_128_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0,
      COMP_LOOP_5_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_160_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_160_tr0,
      COMP_LOOP_6_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_192_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0,
      COMP_LOOP_7_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_224_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_224_tr0,
      COMP_LOOP_8_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_256_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0,
      COMP_LOOP_9_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_288_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_288_tr0,
      COMP_LOOP_10_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_320_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0,
      COMP_LOOP_11_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_352_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_352_tr0,
      COMP_LOOP_12_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_384_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0,
      COMP_LOOP_13_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_416_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_416_tr0,
      COMP_LOOP_14_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_448_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0,
      COMP_LOOP_15_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_480_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_480_tr0,
      COMP_LOOP_16_modExp_dev_1_while_C_14_tr0 => COMP_LOOP_COMP_LOOP_and_137_itm,
      COMP_LOOP_C_512_tr0 => COMP_LOOP_COMP_LOOP_and_10_itm,
      VEC_LOOP_C_0_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_4_tr0 => inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_4_tr0
    );
  fsm_output <= inPlaceNTT_DIT_core_core_fsm_inst_fsm_output;
  inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_3_tr0 <= NOT (z_out_8_64_2(62));
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 <= NOT COMP_LOOP_nor_11_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_32_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_96_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_160_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_224_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_288_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_352_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_416_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0 <= NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_480_tr0 <= NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 <= VEC_LOOP_acc_1_psp_1(10);
  inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_4_tr0 <= NOT (z_out_8_64_2(0));

  nand_308_cse <= NOT((z_out_6_10_1(0)) AND (fsm_output(5)) AND (fsm_output(7)) AND
      (fsm_output(4)));
  nand_270_cse_1 <= NOT((z_out_6_10_1(3)) AND (fsm_output(5)) AND (fsm_output(7))
      AND (fsm_output(4)));
  nand_264_cse <= NOT((z_out_6_10_1(3)) AND (z_out_6_10_1(0)) AND (fsm_output(5))
      AND (fsm_output(7)) AND (fsm_output(4)));
  nand_260_cse_1 <= NOT((z_out_6_10_1(1)) AND (z_out_6_10_1(3)) AND (fsm_output(5))
      AND (fsm_output(7)) AND (fsm_output(4)));
  or_2146_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"));
  and_357_cse <= (fsm_output(0)) AND (fsm_output(2)) AND (fsm_output(3));
  mux_1575_nl <= MUX_s_1_2_2((NOT (fsm_output(9))), nor_tmp_14, fsm_output(3));
  mux_1576_nl <= MUX_s_1_2_2(mux_1575_nl, mux_461_cse, fsm_output(2));
  mux_1574_nl <= MUX_s_1_2_2(mux_tmp_1514, mux_tmp_1488, fsm_output(0));
  mux_1577_nl <= MUX_s_1_2_2(mux_1576_nl, mux_1574_nl, fsm_output(6));
  mux_1578_nl <= MUX_s_1_2_2(mux_1577_nl, mux_tmp_1498, fsm_output(7));
  mux_1570_nl <= MUX_s_1_2_2(mux_424_cse, nor_tmp_14, or_214_cse);
  mux_1571_nl <= MUX_s_1_2_2(mux_1570_nl, mux_tmp_1496, fsm_output(0));
  and_278_nl <= (and_357_cse OR (fsm_output(9))) AND (fsm_output(8));
  mux_1572_nl <= MUX_s_1_2_2(mux_1571_nl, and_278_nl, fsm_output(6));
  mux_1569_nl <= MUX_s_1_2_2(mux_tmp_1503, mux_tmp_1501, fsm_output(6));
  mux_1573_nl <= MUX_s_1_2_2(mux_1572_nl, mux_1569_nl, fsm_output(7));
  mux_1579_nl <= MUX_s_1_2_2(mux_1578_nl, mux_1573_nl, fsm_output(5));
  mux_1566_nl <= MUX_s_1_2_2(mux_tmp_1514, mux_tmp_1496, fsm_output(6));
  mux_1567_nl <= MUX_s_1_2_2(mux_1566_nl, mux_tmp_1477, fsm_output(7));
  and_280_nl <= ((NOT((fsm_output(0)) OR (fsm_output(2)) OR (fsm_output(3)))) OR
      (fsm_output(9))) AND (fsm_output(8));
  mux_1562_nl <= MUX_s_1_2_2(and_280_nl, mux_tmp_1489, fsm_output(6));
  mux_1561_nl <= MUX_s_1_2_2(mux_tmp_1485, nor_tmp_190, fsm_output(6));
  mux_1563_nl <= MUX_s_1_2_2(mux_1562_nl, mux_1561_nl, fsm_output(7));
  mux_1568_nl <= MUX_s_1_2_2(mux_1567_nl, mux_1563_nl, fsm_output(5));
  mux_1580_nl <= MUX_s_1_2_2(mux_1579_nl, mux_1568_nl, fsm_output(4));
  mux_1555_nl <= MUX_s_1_2_2(nor_697_cse, nor_tmp_14, or_2146_cse);
  mux_1556_nl <= MUX_s_1_2_2(mux_1555_nl, mux_tmp_1482, fsm_output(0));
  mux_1557_nl <= MUX_s_1_2_2(mux_1556_nl, mux_tmp_1503, fsm_output(6));
  mux_1551_nl <= MUX_s_1_2_2(nor_tmp_14, mux_tmp_1470, fsm_output(0));
  mux_1553_nl <= MUX_s_1_2_2(mux_tmp_1501, mux_1551_nl, fsm_output(6));
  mux_1558_nl <= MUX_s_1_2_2(mux_1557_nl, mux_1553_nl, fsm_output(7));
  mux_1544_nl <= MUX_s_1_2_2(nor_tmp_186, mux_tmp_1471, fsm_output(2));
  mux_1545_nl <= MUX_s_1_2_2(mux_tmp_1473, mux_1544_nl, fsm_output(0));
  mux_1546_nl <= MUX_s_1_2_2(mux_tmp_1476, mux_1545_nl, fsm_output(6));
  mux_1550_nl <= MUX_s_1_2_2(mux_tmp_1498, mux_1546_nl, fsm_output(7));
  mux_1559_nl <= MUX_s_1_2_2(mux_1558_nl, mux_1550_nl, fsm_output(5));
  mux_1541_nl <= MUX_s_1_2_2(mux_tmp_1489, mux_tmp_1485, fsm_output(6));
  mux_1530_nl <= MUX_s_1_2_2((fsm_output(9)), nor_tmp_14, or_214_cse);
  mux_1531_nl <= MUX_s_1_2_2(mux_tmp_1476, mux_1530_nl, fsm_output(0));
  mux_1532_nl <= MUX_s_1_2_2(nor_tmp_190, mux_1531_nl, fsm_output(6));
  mux_1542_nl <= MUX_s_1_2_2(mux_1541_nl, mux_1532_nl, fsm_output(7));
  mux_1525_nl <= MUX_s_1_2_2(mux_tmp_1473, mux_tmp_1470, fsm_output(6));
  mux_1529_nl <= MUX_s_1_2_2(mux_tmp_1477, mux_1525_nl, fsm_output(7));
  mux_1543_nl <= MUX_s_1_2_2(mux_1542_nl, mux_1529_nl, fsm_output(5));
  mux_1560_nl <= MUX_s_1_2_2(mux_1559_nl, mux_1543_nl, fsm_output(4));
  mux_1581_itm <= MUX_s_1_2_2(mux_1580_nl, mux_1560_nl, fsm_output(1));
  or_1973_cse <= (fsm_output(6)) OR (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR (fsm_output(3)) OR (fsm_output(8));
  nor_256_cse <= NOT((fsm_output(4)) OR (fsm_output(6)) OR (fsm_output(2)) OR (NOT
      (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(8)));
  or_1916_cse <= (NOT (fsm_output(8))) OR (fsm_output(9)) OR (fsm_output(3));
  or_1982_cse <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (fsm_output(9)) OR (NOT (fsm_output(8)));
  or_1967_cse <= (NOT (fsm_output(6))) OR (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(9))
      OR (fsm_output(3)) OR (fsm_output(8));
  or_1977_cse <= (NOT (fsm_output(2))) OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(3))
      OR (fsm_output(8));
  or_1976_cse <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(3))
      OR (fsm_output(8));
  mux_1788_cse <= MUX_s_1_2_2(or_1977_cse, or_1976_cse, fsm_output(6));
  or_1995_cse <= (fsm_output(2)) OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9))
      OR (NOT (fsm_output(8)));
  mux_1802_cse <= MUX_s_1_2_2(or_1995_cse, or_1977_cse, fsm_output(6));
  mux_1797_cse <= MUX_s_1_2_2(nand_357_cse, or_279_cse, fsm_output(6));
  or_1980_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(9))
      OR nand_321_cse;
  mux_1789_cse <= MUX_s_1_2_2(or_1980_nl, or_279_cse, fsm_output(6));
  mux_1784_cse <= MUX_s_1_2_2(or_279_cse, nand_tmp_106, fsm_output(6));
  mux_1785_cse <= MUX_s_1_2_2(mux_1784_cse, or_1973_cse, fsm_output(4));
  and_259_cse <= (fsm_output(4)) AND (NOT mux_1602_cse);
  mux_1725_nl <= MUX_s_1_2_2(or_2306_cse, mux_tmp_1610, fsm_output(2));
  mux_1726_cse <= MUX_s_1_2_2(mux_1725_nl, mux_tmp_1623, fsm_output(1));
  modExp_dev_while_mux_2_nl <= MUX_v_64_2_2(operator_64_false_acc_mut_63_0, modExp_dev_result_sva,
      mux_2066_cse);
  modExp_dev_while_mux_3_nl <= MUX_v_64_2_2(modExp_dev_result_sva, r_sva, mux_2066_cse);
  mul_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(UNSIGNED'( UNSIGNED(modExp_dev_while_mux_2_nl)
      * UNSIGNED(modExp_dev_while_mux_3_nl)), 64));
  COMP_LOOP_1_acc_8_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_4_dfm) -
      SIGNED(modulo_dev_cmp_return_rsc_z), 64));
  modExp_dev_while_or_1_nl <= and_dcpl_183 OR not_tmp_402;
  and_258_nl <= (fsm_output(4)) AND (NOT mux_1789_cse);
  nor_255_nl <= NOT((fsm_output(4)) OR mux_1788_cse);
  mux_1790_nl <= MUX_s_1_2_2(and_258_nl, nor_255_nl, fsm_output(5));
  mux_1787_nl <= MUX_s_1_2_2(nor_256_cse, and_259_cse, fsm_output(5));
  mux_1791_nl <= MUX_s_1_2_2(mux_1790_nl, mux_1787_nl, fsm_output(1));
  and_260_nl <= (fsm_output(5)) AND (NOT mux_1785_cse);
  mux_1783_nl <= MUX_s_1_2_2(mux_1602_cse, or_1967_cse, fsm_output(4));
  nor_257_nl <= NOT((fsm_output(5)) OR mux_1783_nl);
  mux_1786_nl <= MUX_s_1_2_2(and_260_nl, nor_257_nl, fsm_output(1));
  mux_1792_nl <= MUX_s_1_2_2(mux_1791_nl, mux_1786_nl, fsm_output(0));
  modExp_dev_while_mux1h_nl <= MUX1HOT_v_64_4_2(STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(mul_nl),
      64)), STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
      modulo_dev_cmp_return_rsc_z, STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(COMP_LOOP_1_acc_8_nl),
      64)), STD_LOGIC_VECTOR'( modExp_dev_while_or_1_nl & mux_1911_cse & mux_1792_nl
      & not_tmp_370));
  mux_1693_nl <= MUX_s_1_2_2(or_1916_cse, or_tmp_1854, fsm_output(7));
  or_1896_nl <= (fsm_output(2)) OR mux_1693_nl;
  mux_1694_nl <= MUX_s_1_2_2(or_1896_nl, mux_tmp_1618, fsm_output(1));
  mux_1691_nl <= MUX_s_1_2_2(or_tmp_1799, mux_tmp_1610, fsm_output(2));
  mux_1692_nl <= MUX_s_1_2_2(mux_1691_nl, or_tmp_1855, fsm_output(1));
  mux_1695_nl <= MUX_s_1_2_2(mux_1694_nl, mux_1692_nl, fsm_output(5));
  mux_1696_nl <= MUX_s_1_2_2(mux_1695_nl, mux_tmp_1621, fsm_output(6));
  mux_1727_nl <= MUX_s_1_2_2(or_2306_cse, or_tmp_1793, fsm_output(2));
  mux_1688_nl <= MUX_s_1_2_2(mux_1727_nl, mux_tmp_1625, fsm_output(1));
  mux_1689_nl <= MUX_s_1_2_2(mux_1688_nl, mux_1726_cse, fsm_output(5));
  mux_1686_nl <= MUX_s_1_2_2(mux_tmp_1629, mux_tmp_1626, fsm_output(5));
  mux_1690_nl <= MUX_s_1_2_2(mux_1689_nl, mux_1686_nl, fsm_output(6));
  mux_1697_nl <= MUX_s_1_2_2(mux_1696_nl, mux_1690_nl, fsm_output(4));
  mux_1683_nl <= MUX_s_1_2_2(mux_1726_cse, mux_tmp_1629, fsm_output(5));
  mux_1713_nl <= MUX_s_1_2_2(mux_tmp_1623, or_1880_cse, fsm_output(1));
  mux_1678_nl <= MUX_s_1_2_2(mux_tmp_1626, mux_1713_nl, fsm_output(5));
  mux_1684_nl <= MUX_s_1_2_2(mux_1683_nl, mux_1678_nl, fsm_output(6));
  mux_1703_nl <= MUX_s_1_2_2(mux_tmp_1610, mux_1583_cse, fsm_output(2));
  mux_1667_nl <= MUX_s_1_2_2(or_tmp_1855, mux_1703_nl, fsm_output(1));
  mux_1664_nl <= MUX_s_1_2_2(mux_tmp_1612, or_1880_cse, fsm_output(1));
  mux_1668_nl <= MUX_s_1_2_2(mux_1667_nl, mux_1664_nl, fsm_output(5));
  mux_1673_nl <= MUX_s_1_2_2(mux_tmp_1621, mux_1668_nl, fsm_output(6));
  mux_1685_nl <= MUX_s_1_2_2(mux_1684_nl, mux_1673_nl, fsm_output(4));
  mux_1698_nl <= MUX_s_1_2_2(mux_1697_nl, mux_1685_nl, fsm_output(0));
  operator_64_false_operator_64_false_mux_rgt <= MUX_v_65_2_2(('0' & modExp_dev_while_mux1h_nl),
      z_out_9, mux_1698_nl);
  or_2306_cse <= (fsm_output(7)) OR (NOT (fsm_output(8))) OR (fsm_output(3)) OR (fsm_output(9));
  nor_810_cse <= NOT((NOT (fsm_output(0))) OR (fsm_output(4)));
  and_418_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_267_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_195_rgt <= and_dcpl_132 AND and_dcpl_48;
  or_2012_cse <= (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(8));
  modExp_dev_while_or_2_cse <= and_dcpl_36 OR and_dcpl_44 OR and_dcpl_52 OR and_dcpl_58
      OR and_dcpl_63 OR and_dcpl_72 OR and_dcpl_78 OR and_dcpl_84 OR and_dcpl_90
      OR and_dcpl_93 OR and_dcpl_97 OR and_dcpl_102 OR and_dcpl_106 OR and_dcpl_110
      OR and_dcpl_115 OR and_dcpl_119;
  or_2186_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  or_2040_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  or_103_cse <= (fsm_output(5)) OR (fsm_output(4)) OR (fsm_output(7));
  and_375_cse <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"));
  and_376_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"));
  and_247_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  mux_424_cse <= MUX_s_1_2_2((NOT (fsm_output(8))), (fsm_output(8)), fsm_output(9));
  or_214_cse <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01"));
  or_212_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"));
  mux_461_cse <= MUX_s_1_2_2(mux_424_cse, nor_tmp_14, fsm_output(3));
  mux_459_nl <= MUX_s_1_2_2(mux_424_cse, (fsm_output(9)), fsm_output(3));
  mux_460_cse <= MUX_s_1_2_2(mux_459_nl, nor_tmp_14, fsm_output(2));
  nor_697_cse <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00")));
  mux_1904_nl <= MUX_s_1_2_2(mux_1797_cse, mux_1788_cse, fsm_output(4));
  nor_760_cse <= NOT((fsm_output(5)) OR mux_1904_nl);
  nor_758_nl <= NOT((fsm_output(4)) OR mux_1802_cse);
  and_256_nl <= (fsm_output(4)) AND (NOT mux_1797_cse);
  mux_1909_cse <= MUX_s_1_2_2(nor_758_nl, and_256_nl, fsm_output(5));
  mux_1800_nl <= MUX_s_1_2_2(or_279_cse, nand_tmp, fsm_output(6));
  and_445_nl <= (fsm_output(4)) AND (NOT mux_1800_nl);
  mux_1907_nl <= MUX_s_1_2_2(and_445_nl, nor_256_cse, fsm_output(5));
  mux_1910_nl <= MUX_s_1_2_2(mux_1909_cse, mux_1907_nl, fsm_output(1));
  mux_1794_nl <= MUX_s_1_2_2(nand_tmp, or_1982_cse, fsm_output(6));
  mux_1901_nl <= MUX_s_1_2_2(mux_1794_nl, or_1967_cse, fsm_output(4));
  and_446_nl <= (fsm_output(5)) AND (NOT mux_1901_nl);
  mux_1905_nl <= MUX_s_1_2_2(nor_760_cse, and_446_nl, fsm_output(1));
  mux_1911_cse <= MUX_s_1_2_2(mux_1910_nl, mux_1905_nl, fsm_output(0));
  mux_1949_cse <= MUX_s_1_2_2((fsm_output(8)), or_tmp_2044, fsm_output(3));
  or_2336_cse <= (NOT((fsm_output(3)) OR (NOT (fsm_output(9))))) OR (fsm_output(8));
  COMP_LOOP_k_COMP_LOOP_k_mux_nl <= MUX_v_5_2_2(COMP_LOOP_k_9_4_sva_4_0, (z_out_9(8
      DOWNTO 4)), not_tmp_402);
  COMP_LOOP_mux1h_192_rgt <= MUX_v_10_2_2((STD_LOGIC_VECTOR'( "00000") & COMP_LOOP_k_COMP_LOOP_k_mux_nl),
      z_out_6_10_1, modExp_dev_while_or_2_cse);
  or_2348_cse <= (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(1));
  or_279_cse <= (fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(9))) OR (fsm_output(8))
      OR (NOT (fsm_output(3)));
  COMP_LOOP_acc_13_psp_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0(9
      DOWNTO 2)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 &
      STD_LOGIC_VECTOR'( "01")), 7), 8), 8));
  COMP_LOOP_acc_1_cse_2_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
      "0001")), 9), 10), 10));
  VEC_LOOP_acc_1_psp_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      10), 11), 11));
  nor_728_cse <= NOT((fsm_output(3)) OR (NOT (fsm_output(9))) OR (fsm_output(8)));
  nor_727_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(8))));
  mux_51_nl <= MUX_s_1_2_2(nor_727_nl, nor_728_cse, fsm_output(7));
  nand_tmp <= NOT((fsm_output(2)) AND mux_51_nl);
  nand_357_cse <= NOT((fsm_output(2)) AND (fsm_output(7)) AND (fsm_output(3)) AND
      (NOT (fsm_output(9))) AND (fsm_output(8)));
  or_tmp_20 <= (fsm_output(5)) OR and_375_cse;
  nor_tmp_14 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("11"));
  or_tmp_74 <= (fsm_output(5)) OR (fsm_output(7));
  nor_tmp_40 <= (fsm_output(5)) AND (fsm_output(7));
  nand_321_cse <= NOT((fsm_output(3)) AND (fsm_output(8)));
  and_dcpl_13 <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_14 <= and_dcpl_13 AND (NOT (fsm_output(6)));
  and_dcpl_15 <= and_dcpl_14 AND nor_697_cse;
  and_dcpl_16 <= NOT((fsm_output(4)) OR (fsm_output(0)));
  and_dcpl_17 <= NOT((fsm_output(5)) OR (fsm_output(7)));
  and_dcpl_18 <= and_dcpl_17 AND (NOT (fsm_output(3)));
  and_dcpl_19 <= and_dcpl_18 AND and_dcpl_16;
  and_dcpl_23 <= and_418_cse AND (NOT (fsm_output(6)));
  or_2152_nl <= (fsm_output(9)) OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(1))
      OR (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(7))
      OR (fsm_output(5));
  nand_314_nl <= NOT((fsm_output(9)) AND ((fsm_output(6)) OR and_247_cse OR (fsm_output(5))
      OR (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(7))));
  not_tmp_121 <= MUX_s_1_2_2(or_2152_nl, nand_314_nl, fsm_output(8));
  and_dcpl_26 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_27 <= and_dcpl_26 AND (NOT (fsm_output(6)));
  and_dcpl_28 <= and_dcpl_27 AND nor_697_cse;
  and_dcpl_29 <= (fsm_output(4)) AND (NOT (fsm_output(0)));
  and_dcpl_30 <= and_dcpl_18 AND and_dcpl_29;
  and_dcpl_32 <= (NOT (fsm_output(4))) AND (fsm_output(0));
  and_dcpl_33 <= (fsm_output(5)) AND (NOT (fsm_output(7)));
  and_dcpl_34 <= and_dcpl_33 AND (NOT (fsm_output(3)));
  and_dcpl_35 <= and_dcpl_34 AND and_dcpl_32;
  and_dcpl_36 <= and_dcpl_35 AND and_dcpl_28;
  and_dcpl_37 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_38 <= and_dcpl_37 AND (fsm_output(6));
  and_dcpl_39 <= and_dcpl_38 AND nor_697_cse;
  and_dcpl_40 <= and_dcpl_18 AND and_dcpl_32;
  and_dcpl_42 <= and_dcpl_26 AND (fsm_output(6));
  and_dcpl_43 <= and_dcpl_42 AND nor_697_cse;
  and_dcpl_44 <= and_dcpl_30 AND and_dcpl_43;
  and_dcpl_45 <= and_dcpl_34 AND and_dcpl_29;
  and_dcpl_47 <= and_dcpl_37 AND (NOT (fsm_output(6)));
  and_dcpl_48 <= and_dcpl_47 AND nor_697_cse;
  and_dcpl_49 <= (NOT (fsm_output(5))) AND (fsm_output(7));
  and_dcpl_50 <= and_dcpl_49 AND (NOT (fsm_output(3)));
  and_dcpl_51 <= and_dcpl_50 AND and_dcpl_32;
  and_dcpl_52 <= and_dcpl_51 AND and_dcpl_48;
  and_dcpl_54 <= nor_tmp_40 AND (NOT (fsm_output(3)));
  and_dcpl_55 <= and_dcpl_54 AND and_dcpl_32;
  and_dcpl_57 <= and_dcpl_54 AND and_dcpl_29;
  and_dcpl_58 <= and_dcpl_57 AND and_dcpl_48;
  and_dcpl_59 <= and_dcpl_13 AND (fsm_output(6));
  and_dcpl_60 <= and_dcpl_59 AND nor_697_cse;
  and_dcpl_61 <= and_dcpl_50 AND and_dcpl_29;
  and_dcpl_63 <= and_dcpl_55 AND and_dcpl_60;
  and_dcpl_64 <= and_418_cse AND (fsm_output(6));
  and_dcpl_65 <= and_dcpl_64 AND nor_697_cse;
  and_dcpl_66 <= (fsm_output(4)) AND (fsm_output(0));
  and_dcpl_67 <= nor_tmp_40 AND (fsm_output(3));
  and_dcpl_68 <= and_dcpl_67 AND and_dcpl_66;
  and_dcpl_70 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_71 <= and_dcpl_14 AND and_dcpl_70;
  and_dcpl_72 <= and_dcpl_30 AND and_dcpl_71;
  and_dcpl_73 <= and_dcpl_23 AND and_dcpl_70;
  and_dcpl_74 <= and_dcpl_33 AND (fsm_output(3));
  and_dcpl_75 <= and_dcpl_74 AND and_dcpl_16;
  and_dcpl_78 <= and_dcpl_74 AND and_dcpl_66 AND and_dcpl_73;
  and_dcpl_79 <= and_dcpl_42 AND and_dcpl_70;
  and_dcpl_80 <= and_dcpl_17 AND (fsm_output(3));
  and_dcpl_81 <= and_dcpl_80 AND and_dcpl_66;
  and_dcpl_83 <= and_dcpl_64 AND and_dcpl_70;
  and_dcpl_84 <= and_dcpl_75 AND and_dcpl_83;
  and_dcpl_85 <= and_dcpl_27 AND and_dcpl_70;
  and_dcpl_86 <= and_dcpl_49 AND (fsm_output(3));
  and_dcpl_87 <= and_dcpl_86 AND and_dcpl_16;
  and_dcpl_89 <= and_dcpl_86 AND and_dcpl_66;
  and_dcpl_90 <= and_dcpl_89 AND and_dcpl_85;
  and_dcpl_91 <= and_dcpl_47 AND and_dcpl_70;
  and_dcpl_93 <= and_dcpl_87 AND and_dcpl_79;
  and_dcpl_94 <= and_dcpl_38 AND and_dcpl_70;
  and_dcpl_95 <= and_dcpl_67 AND and_dcpl_16;
  and_dcpl_97 <= and_dcpl_68 AND and_dcpl_94;
  and_dcpl_98 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_99 <= and_dcpl_14 AND and_dcpl_98;
  and_dcpl_101 <= and_dcpl_47 AND and_dcpl_98;
  and_dcpl_102 <= and_dcpl_75 AND and_dcpl_101;
  and_dcpl_103 <= and_dcpl_59 AND and_dcpl_98;
  and_dcpl_106 <= and_dcpl_81 AND and_dcpl_103;
  and_dcpl_107 <= and_dcpl_64 AND and_dcpl_98;
  and_dcpl_108 <= and_dcpl_34 AND and_dcpl_66;
  and_dcpl_110 <= and_dcpl_87 AND and_dcpl_99;
  and_dcpl_111 <= and_dcpl_23 AND and_dcpl_98;
  and_dcpl_112 <= and_dcpl_54 AND and_dcpl_16;
  and_dcpl_115 <= and_dcpl_54 AND and_dcpl_66 AND and_dcpl_111;
  and_dcpl_116 <= and_dcpl_42 AND and_dcpl_98;
  and_dcpl_117 <= and_dcpl_50 AND and_dcpl_66;
  and_dcpl_119 <= and_dcpl_112 AND and_dcpl_107;
  or_tmp_237 <= (NOT (fsm_output(9))) OR (fsm_output(8)) OR (fsm_output(3));
  or_265_nl <= (fsm_output(9)) OR (fsm_output(8)) OR (NOT (fsm_output(3)));
  mux_514_nl <= MUX_s_1_2_2(or_tmp_237, or_265_nl, fsm_output(7));
  nand_tmp_6 <= NOT((fsm_output(2)) AND (NOT mux_514_nl));
  or_tmp_239 <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (fsm_output(9)) OR nand_321_cse;
  or_tmp_241 <= (fsm_output(9)) OR nand_321_cse;
  mux_520_nl <= MUX_s_1_2_2(or_tmp_241, or_tmp_237, fsm_output(7));
  nand_tmp_7 <= NOT((fsm_output(2)) AND (NOT mux_520_nl));
  and_dcpl_122 <= and_dcpl_23 AND nor_697_cse;
  and_dcpl_130 <= and_dcpl_59 AND and_dcpl_70;
  and_dcpl_132 <= and_dcpl_18 AND and_dcpl_66;
  and_dcpl_136 <= and_dcpl_27 AND and_dcpl_98;
  and_dcpl_138 <= and_dcpl_38 AND and_dcpl_98;
  or_tmp_252 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  or_tmp_253 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  or_tmp_258 <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  or_tmp_259 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  not_tmp_133 <= NOT((fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(4)));
  not_tmp_134 <= NOT((fsm_output(7)) AND (fsm_output(4)));
  or_tmp_346 <= (fsm_output(1)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"));
  or_tmp_352 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"));
  or_tmp_353 <= (NOT (fsm_output(1))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"));
  or_tmp_362 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"));
  or_tmp_438 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  or_tmp_439 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  or_tmp_444 <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  or_tmp_445 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  or_tmp_531 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"));
  or_tmp_532 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"));
  or_tmp_537 <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"));
  or_tmp_538 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"));
  or_tmp_624 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"));
  or_tmp_625 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"));
  or_tmp_630 <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"));
  or_tmp_631 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"));
  or_tmp_718 <= (fsm_output(1)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"));
  or_tmp_724 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"));
  or_tmp_725 <= (NOT (fsm_output(1))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"));
  or_tmp_734 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"));
  or_tmp_810 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"));
  or_tmp_811 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"));
  or_tmp_816 <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"));
  or_tmp_817 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"));
  or_tmp_903 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"));
  or_tmp_904 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"));
  or_tmp_909 <= NOT((fsm_output(5)) AND (fsm_output(1)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("0111")));
  or_tmp_910 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"));
  or_tmp_997 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  or_tmp_999 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  or_tmp_1005 <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  or_tmp_1007 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  or_tmp_1097 <= (fsm_output(1)) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"));
  or_tmp_1104 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"));
  or_tmp_1106 <= (NOT (fsm_output(1))) OR (fsm_output(5)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"));
  or_tmp_1116 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"));
  or_tmp_1195 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  or_tmp_1197 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  or_tmp_1203 <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  or_tmp_1205 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  or_tmp_1294 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"));
  or_tmp_1296 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"));
  or_tmp_1302 <= NOT((fsm_output(5)) AND (fsm_output(1)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1011")));
  or_tmp_1304 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"));
  not_tmp_289 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11")));
  or_tmp_1393 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_289;
  or_tmp_1395 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_289;
  or_tmp_1401 <= (NOT (fsm_output(5))) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_289;
  or_tmp_1403 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_289;
  not_tmp_304 <= NOT((COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(0)) AND (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(2))
      AND (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3)));
  or_tmp_1493 <= (fsm_output(1)) OR (NOT (fsm_output(5))) OR (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1))
      OR not_tmp_304;
  or_tmp_1500 <= (NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1))
      OR not_tmp_304;
  or_tmp_1502 <= (NOT (fsm_output(1))) OR (fsm_output(5)) OR (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1))
      OR not_tmp_304;
  or_tmp_1512 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))
      OR (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1)) OR not_tmp_304;
  or_tmp_1590 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_289;
  or_tmp_1592 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR not_tmp_289;
  or_tmp_1598 <= (NOT((fsm_output(5)) AND (fsm_output(1)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("10")))) OR not_tmp_289;
  or_tmp_1600 <= (fsm_output(5)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR not_tmp_289;
  not_tmp_335 <= NOT(CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")));
  or_tmp_1687 <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1))
      OR not_tmp_335;
  or_tmp_1689 <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR not_tmp_335;
  not_tmp_336 <= NOT((fsm_output(5)) AND (fsm_output(1)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111")));
  or_tmp_1694 <= (fsm_output(5)) OR (NOT((fsm_output(1)) AND CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))));
  or_2151_cse <= (fsm_output(3)) OR (fsm_output(9));
  nor_tmp_186 <= or_2151_cse AND (fsm_output(8));
  mux_1520_nl <= MUX_s_1_2_2(nor_tmp_14, mux_424_cse, fsm_output(3));
  mux_tmp_1470 <= MUX_s_1_2_2(nor_tmp_186, mux_1520_nl, fsm_output(2));
  mux_tmp_1471 <= MUX_s_1_2_2((fsm_output(9)), nor_tmp_14, fsm_output(3));
  mux_tmp_1472 <= MUX_s_1_2_2((NOT (fsm_output(8))), (fsm_output(8)), or_2151_cse);
  mux_tmp_1473 <= MUX_s_1_2_2(mux_tmp_1472, mux_tmp_1471, fsm_output(2));
  mux_tmp_1476 <= MUX_s_1_2_2(mux_461_cse, mux_tmp_1471, fsm_output(2));
  nor_tmp_188 <= (and_376_cse OR (fsm_output(9))) AND (fsm_output(8));
  mux_tmp_1477 <= MUX_s_1_2_2(nor_tmp_188, mux_tmp_1476, fsm_output(6));
  nor_tmp_190 <= ((NOT((fsm_output(0)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(3)))))
      OR (fsm_output(9))) AND (fsm_output(8));
  mux_tmp_1482 <= MUX_s_1_2_2(mux_461_cse, nor_tmp_186, fsm_output(2));
  mux_tmp_1483 <= MUX_s_1_2_2(nor_tmp_14, (fsm_output(9)), fsm_output(3));
  mux_tmp_1484 <= MUX_s_1_2_2(mux_tmp_1483, nor_tmp_186, fsm_output(2));
  mux_tmp_1485 <= MUX_s_1_2_2(mux_tmp_1484, mux_tmp_1482, fsm_output(0));
  mux_tmp_1488 <= MUX_s_1_2_2(mux_tmp_1483, mux_461_cse, fsm_output(2));
  mux_tmp_1489 <= MUX_s_1_2_2(mux_tmp_1488, mux_460_cse, fsm_output(0));
  mux_tmp_1496 <= MUX_s_1_2_2(mux_tmp_1483, mux_tmp_1472, fsm_output(2));
  mux_1548_nl <= MUX_s_1_2_2(mux_tmp_1496, mux_tmp_1484, fsm_output(0));
  mux_tmp_1498 <= MUX_s_1_2_2(mux_1548_nl, nor_tmp_188, fsm_output(6));
  mux_tmp_1501 <= MUX_s_1_2_2(mux_tmp_1482, mux_tmp_1473, fsm_output(0));
  mux_tmp_1503 <= MUX_s_1_2_2(mux_460_cse, mux_tmp_1476, fsm_output(0));
  mux_1564_nl <= MUX_s_1_2_2((fsm_output(8)), (fsm_output(9)), fsm_output(3));
  mux_tmp_1514 <= MUX_s_1_2_2(mux_1564_nl, mux_461_cse, fsm_output(2));
  or_tmp_1788 <= (NOT (fsm_output(7))) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(8));
  or_tmp_1793 <= NOT((fsm_output(7)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (fsm_output(8)));
  or_tmp_1794 <= (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(9)))
      OR (fsm_output(8));
  or_1820_cse <= (NOT (fsm_output(3))) OR (fsm_output(9)) OR (NOT (fsm_output(8)));
  mux_1583_cse <= MUX_s_1_2_2(or_1820_cse, or_tmp_237, fsm_output(7));
  mux_1584_nl <= MUX_s_1_2_2(or_tmp_1793, mux_1583_cse, fsm_output(6));
  mux_tmp_1534 <= MUX_s_1_2_2(or_tmp_1794, mux_1584_nl, fsm_output(2));
  or_tmp_1796 <= (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9)) OR (fsm_output(8));
  mux_1587_nl <= MUX_s_1_2_2(or_2306_cse, or_tmp_1788, fsm_output(6));
  mux_tmp_1537 <= MUX_s_1_2_2(mux_1587_nl, or_tmp_1796, fsm_output(2));
  or_tmp_1799 <= NOT((fsm_output(7)) AND (fsm_output(3)) AND (fsm_output(9)) AND
      (NOT (fsm_output(8))));
  nor_275_nl <= NOT((fsm_output(9)) OR nand_321_cse);
  mux_1601_nl <= MUX_s_1_2_2(nor_275_nl, nor_728_cse, fsm_output(7));
  nand_tmp_106 <= NOT((fsm_output(2)) AND mux_1601_nl);
  mux_1602_cse <= MUX_s_1_2_2(nand_tmp_106, or_tmp_239, fsm_output(6));
  mux_1610_nl <= MUX_s_1_2_2(mux_1789_cse, mux_1788_cse, fsm_output(4));
  and_272_nl <= (fsm_output(5)) AND (NOT mux_1610_nl);
  nor_272_nl <= NOT((fsm_output(5)) OR mux_1785_cse);
  mux_1611_nl <= MUX_s_1_2_2(and_272_nl, nor_272_nl, fsm_output(1));
  nor_273_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR
      (NOT (fsm_output(7))) OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(8)));
  and_273_nl <= (fsm_output(4)) AND (NOT mux_1784_cse);
  mux_1605_nl <= MUX_s_1_2_2(nor_273_nl, and_273_nl, fsm_output(5));
  nor_274_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR
      (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(3)) OR (fsm_output(8)));
  mux_1603_nl <= MUX_s_1_2_2(and_259_cse, nor_274_nl, fsm_output(5));
  mux_1606_nl <= MUX_s_1_2_2(mux_1605_nl, mux_1603_nl, fsm_output(1));
  not_tmp_370 <= MUX_s_1_2_2(mux_1611_nl, mux_1606_nl, fsm_output(0));
  or_tmp_1816 <= (fsm_output(6)) OR (fsm_output(5)) OR (fsm_output(9)) OR (NOT (fsm_output(8)));
  or_tmp_1818 <= NOT((fsm_output(6)) AND (fsm_output(5)) AND (NOT (fsm_output(9)))
      AND (fsm_output(8)));
  mux_tmp_1562 <= MUX_s_1_2_2(or_tmp_1818, or_tmp_1816, fsm_output(1));
  or_1849_nl <= (NOT (fsm_output(5))) OR (fsm_output(9)) OR (NOT (fsm_output(8)));
  mux_tmp_1563 <= MUX_s_1_2_2(or_1849_nl, or_tmp_1816, fsm_output(1));
  or_tmp_1823 <= (fsm_output(6)) OR (fsm_output(5)) OR (NOT (fsm_output(9))) OR (fsm_output(8));
  or_tmp_1824 <= NOT((fsm_output(6)) AND (fsm_output(5)) AND (fsm_output(9)) AND
      (NOT (fsm_output(8))));
  mux_tmp_1566 <= MUX_s_1_2_2(or_tmp_1824, or_tmp_1823, fsm_output(1));
  or_tmp_1825 <= (fsm_output(6)) OR (fsm_output(5)) OR (fsm_output(9)) OR (fsm_output(8));
  or_tmp_1827 <= (NOT (fsm_output(6))) OR (fsm_output(5)) OR (NOT (fsm_output(9)))
      OR (fsm_output(8));
  or_tmp_1830 <= (NOT (fsm_output(6))) OR (fsm_output(5)) OR (fsm_output(9)) OR (NOT
      (fsm_output(8)));
  or_tmp_1831 <= (fsm_output(6)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(9)))
      OR (fsm_output(8));
  mux_tmp_1573 <= MUX_s_1_2_2(or_tmp_1831, or_tmp_1830, fsm_output(1));
  or_tmp_1835 <= (NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (fsm_output(9))
      OR (fsm_output(8));
  or_1863_nl <= (fsm_output(5)) OR (fsm_output(9)) OR (fsm_output(8));
  mux_tmp_1579 <= MUX_s_1_2_2(or_tmp_1835, or_1863_nl, fsm_output(1));
  or_tmp_1838 <= (NOT (fsm_output(6))) OR (fsm_output(5)) OR (fsm_output(9)) OR (fsm_output(8));
  or_tmp_1840 <= (fsm_output(6)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (NOT
      (fsm_output(8)));
  or_tmp_1841 <= (fsm_output(6)) OR (NOT (fsm_output(5))) OR (fsm_output(9)) OR (fsm_output(8));
  and_dcpl_169 <= and_dcpl_18 AND (NOT (fsm_output(4))) AND (fsm_output(1)) AND (NOT
      (fsm_output(2))) AND (NOT (fsm_output(6))) AND nor_697_cse;
  or_tmp_1845 <= and_418_cse OR (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(7))
      OR (fsm_output(5));
  and_tmp_12 <= (fsm_output(9)) AND ((fsm_output(6)) OR or_tmp_1845);
  mux_tmp_1610 <= MUX_s_1_2_2(or_2012_cse, or_1820_cse, fsm_output(7));
  or_1880_cse <= (fsm_output(2)) OR mux_tmp_1610;
  mux_tmp_1612 <= MUX_s_1_2_2(or_tmp_1794, mux_1583_cse, fsm_output(2));
  or_tmp_1854 <= (NOT (fsm_output(3))) OR (NOT (fsm_output(9))) OR (fsm_output(8));
  mux_tmp_1615 <= MUX_s_1_2_2(or_tmp_1854, or_2012_cse, fsm_output(7));
  or_tmp_1855 <= (fsm_output(2)) OR mux_tmp_1615;
  mux_tmp_1618 <= MUX_s_1_2_2(mux_tmp_1615, or_tmp_1793, fsm_output(2));
  nand_111_nl <= NOT((fsm_output(2)) AND (NOT mux_tmp_1610));
  mux_1671_nl <= MUX_s_1_2_2(nand_111_nl, mux_tmp_1612, fsm_output(1));
  nand_110_nl <= NOT((fsm_output(2)) AND (NOT mux_1583_cse));
  mux_1670_nl <= MUX_s_1_2_2(mux_tmp_1618, nand_110_nl, fsm_output(1));
  mux_tmp_1621 <= MUX_s_1_2_2(mux_1671_nl, mux_1670_nl, fsm_output(5));
  mux_tmp_1623 <= MUX_s_1_2_2(or_tmp_1788, mux_1583_cse, fsm_output(2));
  mux_tmp_1625 <= MUX_s_1_2_2(mux_tmp_1615, or_tmp_1796, fsm_output(2));
  mux_tmp_1626 <= MUX_s_1_2_2(mux_tmp_1625, or_1982_cse, fsm_output(1));
  mux_1679_nl <= MUX_s_1_2_2(or_tmp_1794, or_tmp_1796, fsm_output(2));
  mux_tmp_1629 <= MUX_s_1_2_2(mux_1679_nl, mux_tmp_1623, fsm_output(1));
  nand_151_nl <= NOT((fsm_output(1)) AND (fsm_output(0)) AND (fsm_output(4)));
  mux_tmp_1688 <= MUX_s_1_2_2(nand_151_nl, or_2348_cse, fsm_output(2));
  or_tmp_1899 <= and_375_cse OR (fsm_output(7)) OR (fsm_output(5));
  and_dcpl_183 <= and_dcpl_40 AND and_dcpl_28;
  nand_342_nl <= NOT((fsm_output(2)) AND (fsm_output(3)) AND (NOT (fsm_output(9)))
      AND (fsm_output(8)));
  or_2000_nl <= (NOT (fsm_output(2))) OR (fsm_output(3)) OR (NOT (fsm_output(9)))
      OR (fsm_output(8));
  mux_1768_cse <= MUX_s_1_2_2(nand_342_nl, or_2000_nl, fsm_output(7));
  or_1996_nl <= (fsm_output(2)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(3)))
      OR (NOT (fsm_output(9))) OR (fsm_output(8));
  mux_1803_nl <= MUX_s_1_2_2(or_1996_nl, nand_357_cse, fsm_output(6));
  mux_1804_nl <= MUX_s_1_2_2(mux_1803_nl, mux_1802_cse, fsm_output(4));
  and_261_nl <= (fsm_output(5)) AND (NOT mux_1804_nl);
  mux_1779_nl <= MUX_s_1_2_2(and_261_nl, nor_760_cse, fsm_output(1));
  mux_1769_nl <= MUX_s_1_2_2(or_279_cse, mux_1768_cse, fsm_output(6));
  and_263_nl <= (fsm_output(4)) AND (NOT mux_1769_nl);
  mux_1770_nl <= MUX_s_1_2_2(and_263_nl, nor_256_cse, fsm_output(5));
  mux_1774_nl <= MUX_s_1_2_2(mux_1909_cse, mux_1770_nl, fsm_output(1));
  not_tmp_402 <= MUX_s_1_2_2(mux_1779_nl, mux_1774_nl, fsm_output(0));
  nor_tmp_203 <= (fsm_output(6)) AND (fsm_output(7)) AND (fsm_output(9));
  not_tmp_418 <= NOT((fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(9)));
  nor_248_nl <= NOT((fsm_output(0)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(9)));
  mux_1827_nl <= MUX_s_1_2_2(nor_248_nl, nor_tmp_203, fsm_output(1));
  mux_1828_nl <= MUX_s_1_2_2(not_tmp_418, mux_1827_nl, fsm_output(2));
  mux_1829_nl <= MUX_s_1_2_2(mux_1828_nl, nor_tmp_203, fsm_output(3));
  mux_1830_nl <= MUX_s_1_2_2(not_tmp_418, mux_1829_nl, fsm_output(4));
  mux_1831_nl <= MUX_s_1_2_2(mux_1830_nl, nor_tmp_203, fsm_output(5));
  mux_1832_itm <= MUX_s_1_2_2(mux_1831_nl, (fsm_output(9)), fsm_output(8));
  or_tmp_1989 <= (fsm_output(5)) OR (NOT nor_tmp_203);
  or_tmp_1990 <= (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(9));
  mux_tmp_1782 <= MUX_s_1_2_2(or_tmp_1990, or_tmp_1989, fsm_output(4));
  mux_1834_itm <= MUX_s_1_2_2(not_tmp_418, nor_tmp_203, fsm_output(5));
  mux_tmp_1786 <= MUX_s_1_2_2((NOT mux_1834_itm), or_tmp_1990, fsm_output(4));
  mux_1843_nl <= MUX_s_1_2_2(or_tmp_1899, or_103_cse, or_2186_cse);
  mux_tmp_1793 <= MUX_s_1_2_2(or_tmp_1899, mux_1843_nl, fsm_output(2));
  mux_tmp_1799 <= MUX_s_1_2_2((NOT (fsm_output(5))), (fsm_output(5)), fsm_output(7));
  mux_tmp_1801 <= MUX_s_1_2_2(mux_tmp_1799, nor_tmp_40, fsm_output(4));
  mux_tmp_1803 <= MUX_s_1_2_2(mux_tmp_1799, nor_tmp_40, and_375_cse);
  mux_tmp_1808 <= MUX_s_1_2_2(nor_tmp_40, (fsm_output(7)), or_2040_cse);
  mux_tmp_1809 <= MUX_s_1_2_2(nor_tmp_40, (fsm_output(7)), fsm_output(4));
  not_tmp_431 <= NOT((fsm_output(6)) OR mux_tmp_1793);
  nor_tmp_215 <= (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(9));
  not_tmp_439 <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(9)));
  nor_244_nl <= NOT((fsm_output(7)) OR (fsm_output(9)));
  and_368_nl <= (fsm_output(9)) AND (fsm_output(7));
  mux_tmp_1839 <= MUX_s_1_2_2(nor_244_nl, and_368_nl, fsm_output(6));
  and_dcpl_199 <= and_dcpl_132 AND and_dcpl_28;
  and_dcpl_200 <= and_dcpl_19 AND and_dcpl_43;
  and_dcpl_201 <= and_dcpl_108 AND and_dcpl_39;
  and_dcpl_202 <= and_dcpl_112 AND and_dcpl_48;
  and_dcpl_203 <= and_dcpl_117 AND and_dcpl_60;
  and_dcpl_204 <= and_dcpl_19 AND and_dcpl_71;
  and_dcpl_206 <= and_dcpl_74 AND and_dcpl_32 AND and_dcpl_73;
  and_dcpl_207 <= and_dcpl_80 AND and_dcpl_29;
  and_dcpl_208 <= and_dcpl_207 AND and_dcpl_83;
  and_dcpl_210 <= and_dcpl_86 AND and_dcpl_32 AND and_dcpl_85;
  and_dcpl_212 <= and_dcpl_67 AND and_dcpl_29 AND and_dcpl_85;
  and_dcpl_214 <= and_dcpl_67 AND and_dcpl_32 AND and_dcpl_94;
  and_dcpl_215 <= and_dcpl_207 AND and_dcpl_101;
  and_dcpl_217 <= and_dcpl_80 AND and_dcpl_32 AND and_dcpl_103;
  and_dcpl_219 <= and_dcpl_74 AND and_dcpl_29 AND and_dcpl_103;
  and_dcpl_220 <= and_dcpl_55 AND and_dcpl_111;
  and_dcpl_221 <= and_dcpl_61 AND and_dcpl_107;
  or_tmp_2035 <= (NOT (fsm_output(2))) OR (fsm_output(9)) OR (fsm_output(8));
  mux_tmp_1861 <= MUX_s_1_2_2(or_tmp_2035, (fsm_output(8)), fsm_output(3));
  or_tmp_2037 <= and_376_cse OR CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"));
  mux_tmp_1863 <= MUX_s_1_2_2(mux_tmp_1861, or_tmp_2037, fsm_output(7));
  or_tmp_2040 <= (NOT((NOT (fsm_output(2))) OR (fsm_output(9)))) OR (fsm_output(8));
  or_tmp_2041 <= (fsm_output(3)) OR or_tmp_2040;
  mux_tmp_1866 <= MUX_s_1_2_2(or_tmp_2041, mux_tmp_1861, fsm_output(7));
  or_tmp_2043 <= (NOT (fsm_output(2))) OR (fsm_output(9)) OR (NOT (fsm_output(8)));
  or_tmp_2044 <= (fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(8));
  mux_1920_cse <= MUX_s_1_2_2(or_tmp_2044, or_tmp_2043, fsm_output(3));
  mux_tmp_1870 <= MUX_s_1_2_2(or_tmp_2037, mux_1920_cse, fsm_output(7));
  or_2086_cse <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"));
  mux_1922_cse <= MUX_s_1_2_2(or_2086_cse, or_tmp_2043, fsm_output(3));
  mux_tmp_1872 <= MUX_s_1_2_2(or_212_cse, mux_1922_cse, fsm_output(7));
  or_tmp_2047 <= (NOT((fsm_output(2)) OR (NOT (fsm_output(9))))) OR (fsm_output(8));
  mux_tmp_1874 <= MUX_s_1_2_2(or_tmp_2035, or_tmp_2047, fsm_output(3));
  mux_tmp_1875 <= MUX_s_1_2_2(mux_tmp_1874, or_tmp_2037, fsm_output(7));
  nand_tmp_134 <= NOT((fsm_output(3)) AND (NOT or_tmp_2047));
  mux_tmp_1876 <= MUX_s_1_2_2(nand_tmp_134, or_tmp_2037, fsm_output(7));
  mux_tmp_1877 <= MUX_s_1_2_2(mux_tmp_1876, mux_tmp_1875, fsm_output(0));
  mux_tmp_1882 <= MUX_s_1_2_2(or_212_cse, or_tmp_2041, fsm_output(7));
  mux_tmp_1883 <= MUX_s_1_2_2(mux_tmp_1882, mux_tmp_1872, fsm_output(0));
  mux_1938_cse <= MUX_s_1_2_2(or_tmp_2040, or_tmp_2044, fsm_output(3));
  mux_tmp_1888 <= MUX_s_1_2_2(mux_1938_cse, mux_tmp_1861, fsm_output(7));
  or_2091_nl <= (NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"));
  mux_tmp_1891 <= MUX_s_1_2_2(or_2091_nl, or_tmp_2041, fsm_output(7));
  STAGE_LOOP_i_3_0_sva_mx0c1 <= and_dcpl_19 AND and_dcpl_23 AND nor_tmp_14;
  VEC_LOOP_j_sva_9_0_mx0c1 <= and_dcpl_40 AND and_dcpl_27 AND nor_tmp_14;
  vec_rsc_0_0_i_d_d_pff <= modulo_dev_cmp_return_rsc_z;
  and_42_nl <= and_dcpl_30 AND and_dcpl_28;
  and_52_nl <= and_dcpl_40 AND and_dcpl_39;
  and_57_nl <= and_dcpl_45 AND and_dcpl_39;
  and_67_nl <= and_dcpl_55 AND and_dcpl_15;
  and_73_nl <= and_dcpl_61 AND and_dcpl_60;
  and_80_nl <= and_dcpl_68 AND and_dcpl_65;
  and_87_nl <= and_dcpl_75 AND and_dcpl_73;
  and_93_nl <= and_dcpl_81 AND and_dcpl_79;
  and_99_nl <= and_dcpl_87 AND and_dcpl_85;
  and_103_nl <= and_dcpl_68 AND and_dcpl_91;
  and_107_nl <= and_dcpl_95 AND and_dcpl_94;
  and_111_nl <= and_dcpl_81 AND and_dcpl_99;
  and_116_nl <= and_dcpl_80 AND and_dcpl_16 AND and_dcpl_103;
  and_120_nl <= and_dcpl_108 AND and_dcpl_107;
  and_124_nl <= and_dcpl_112 AND and_dcpl_111;
  and_129_nl <= and_dcpl_117 AND and_dcpl_116;
  vec_rsc_0_0_i_radr_d_pff <= MUX1HOT_v_6_17_2(z_out_4, (z_out_6_10_1(9 DOWNTO 4)),
      (COMP_LOOP_acc_1_cse_2_sva(9 DOWNTO 4)), (COMP_LOOP_acc_11_psp_sva(8 DOWNTO
      3)), (COMP_LOOP_acc_1_cse_4_sva(9 DOWNTO 4)), (COMP_LOOP_acc_13_psp_sva(7 DOWNTO
      2)), (COMP_LOOP_acc_1_cse_6_sva(9 DOWNTO 4)), (COMP_LOOP_acc_14_psp_sva(8 DOWNTO
      3)), (COMP_LOOP_acc_1_cse_8_sva(9 DOWNTO 4)), (COMP_LOOP_acc_16_psp_sva(6 DOWNTO
      1)), (COMP_LOOP_acc_1_cse_10_sva(9 DOWNTO 4)), (COMP_LOOP_acc_17_psp_sva(8
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_12_sva(9 DOWNTO 4)), (COMP_LOOP_acc_19_psp_sva(7
      DOWNTO 2)), (COMP_LOOP_acc_1_cse_14_sva(9 DOWNTO 4)), (COMP_LOOP_acc_20_psp_sva(8
      DOWNTO 3)), (COMP_LOOP_acc_1_cse_sva(9 DOWNTO 4)), STD_LOGIC_VECTOR'( and_42_nl
      & modExp_dev_while_or_2_cse & and_52_nl & and_57_nl & and_67_nl & and_73_nl
      & and_80_nl & and_87_nl & and_93_nl & and_99_nl & and_103_nl & and_107_nl &
      and_111_nl & and_116_nl & and_120_nl & and_124_nl & and_129_nl));
  and_131_nl <= and_dcpl_40 AND and_dcpl_60;
  mux_524_nl <= MUX_s_1_2_2(or_279_cse, nand_tmp_7, fsm_output(6));
  or_280_nl <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR mux_524_nl;
  mux_521_nl <= MUX_s_1_2_2(nand_tmp_7, or_tmp_239, fsm_output(6));
  mux_522_nl <= MUX_s_1_2_2(or_1973_cse, mux_521_nl, fsm_output(0));
  or_275_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(6))) OR (fsm_output(2))
      OR (fsm_output(7)) OR (fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(3));
  mux_523_nl <= MUX_s_1_2_2(mux_522_nl, or_275_nl, fsm_output(4));
  mux_525_nl <= MUX_s_1_2_2(or_280_nl, mux_523_nl, fsm_output(5));
  or_271_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(8))) OR (fsm_output(3));
  mux_516_nl <= MUX_s_1_2_2(or_271_nl, or_tmp_241, fsm_output(7));
  or_272_nl <= (fsm_output(2)) OR mux_516_nl;
  mux_517_nl <= MUX_s_1_2_2(or_272_nl, nand_tmp_6, fsm_output(6));
  mux_518_nl <= MUX_s_1_2_2(or_1967_cse, mux_517_nl, fsm_output(0));
  or_274_nl <= (fsm_output(4)) OR mux_518_nl;
  mux_515_nl <= MUX_s_1_2_2(or_tmp_239, nand_tmp_6, fsm_output(6));
  or_269_nl <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR mux_515_nl;
  mux_519_nl <= MUX_s_1_2_2(or_274_nl, or_269_nl, fsm_output(5));
  mux_526_nl <= MUX_s_1_2_2(mux_525_nl, mux_519_nl, fsm_output(1));
  and_132_nl <= and_dcpl_45 AND and_dcpl_60;
  and_134_nl <= and_dcpl_89 AND and_dcpl_122;
  and_135_nl <= and_dcpl_87 AND and_dcpl_65;
  and_136_nl <= and_dcpl_68 AND and_dcpl_43;
  and_137_nl <= and_dcpl_75 AND and_dcpl_85;
  and_138_nl <= and_dcpl_81 AND and_dcpl_94;
  and_139_nl <= and_dcpl_87 AND and_dcpl_91;
  and_140_nl <= and_dcpl_68 AND and_dcpl_71;
  and_142_nl <= and_dcpl_95 AND and_dcpl_130;
  and_144_nl <= and_dcpl_132 AND and_dcpl_111;
  and_145_nl <= and_dcpl_19 AND and_dcpl_107;
  and_146_nl <= and_dcpl_108 AND and_dcpl_116;
  and_148_nl <= and_dcpl_112 AND and_dcpl_136;
  and_150_nl <= and_dcpl_117 AND and_dcpl_138;
  and_152_nl <= and_dcpl_19 AND and_dcpl_47 AND nor_tmp_14;
  vec_rsc_0_0_i_wadr_d_pff <= MUX1HOT_v_6_17_2(COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_10_1_1_sva_9_5
      & (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(4))), (COMP_LOOP_acc_1_cse_2_sva(9 DOWNTO
      4)), (COMP_LOOP_acc_11_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_1_cse_4_sva(9 DOWNTO
      4)), (COMP_LOOP_acc_13_psp_sva(7 DOWNTO 2)), (COMP_LOOP_acc_1_cse_6_sva(9 DOWNTO
      4)), (COMP_LOOP_acc_14_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_1_cse_8_sva(9 DOWNTO
      4)), (COMP_LOOP_acc_16_psp_sva(6 DOWNTO 1)), (COMP_LOOP_acc_1_cse_10_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_17_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_1_cse_12_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_19_psp_sva(7 DOWNTO 2)), (COMP_LOOP_acc_1_cse_14_sva(9
      DOWNTO 4)), (COMP_LOOP_acc_20_psp_sva(8 DOWNTO 3)), (COMP_LOOP_acc_1_cse_sva(9
      DOWNTO 4)), STD_LOGIC_VECTOR'( and_131_nl & (NOT mux_526_nl) & and_132_nl &
      and_134_nl & and_135_nl & and_136_nl & and_137_nl & and_138_nl & and_139_nl
      & and_140_nl & and_142_nl & and_144_nl & and_145_nl & and_146_nl & and_148_nl
      & and_150_nl & and_152_nl));
  or_319_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_552_nl <= MUX_s_1_2_2(or_tmp_259, or_319_nl, fsm_output(0));
  or_318_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_551_nl <= MUX_s_1_2_2(or_318_nl, or_tmp_253, fsm_output(0));
  mux_553_nl <= MUX_s_1_2_2(mux_552_nl, mux_551_nl, fsm_output(4));
  nand_10_nl <= NOT((fsm_output(6)) AND (NOT mux_553_nl));
  or_317_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000"));
  mux_554_nl <= MUX_s_1_2_2(nand_10_nl, or_317_nl, fsm_output(7));
  nor_689_nl <= NOT((fsm_output(8)) OR mux_554_nl);
  nor_690_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT
      (fsm_output(1))));
  or_313_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_549_nl <= MUX_s_1_2_2(or_313_nl, or_tmp_259, fsm_output(0));
  nor_691_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_549_nl);
  mux_550_nl <= MUX_s_1_2_2(nor_690_nl, nor_691_nl, fsm_output(8));
  mux_555_nl <= MUX_s_1_2_2(nor_689_nl, mux_550_nl, fsm_output(9));
  or_310_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_308_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_544_nl <= MUX_s_1_2_2(or_308_nl, or_tmp_259, fsm_output(0));
  or_306_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_543_nl <= MUX_s_1_2_2(or_tmp_258, or_306_nl, fsm_output(0));
  mux_545_nl <= MUX_s_1_2_2(mux_544_nl, mux_543_nl, fsm_output(4));
  or_304_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_542_nl <= MUX_s_1_2_2(or_304_nl, or_tmp_253, fsm_output(0));
  or_305_nl <= (fsm_output(4)) OR mux_542_nl;
  mux_546_nl <= MUX_s_1_2_2(mux_545_nl, or_305_nl, fsm_output(6));
  mux_547_nl <= MUX_s_1_2_2(or_310_nl, mux_546_nl, fsm_output(7));
  and_344_nl <= (fsm_output(8)) AND (NOT mux_547_nl);
  nor_692_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
  mux_548_nl <= MUX_s_1_2_2(and_344_nl, nor_692_nl, fsm_output(9));
  mux_556_nl <= MUX_s_1_2_2(mux_555_nl, mux_548_nl, fsm_output(3));
  or_301_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_299_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_537_nl <= MUX_s_1_2_2(or_299_nl, or_tmp_259, fsm_output(0));
  or_297_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_536_nl <= MUX_s_1_2_2(or_tmp_258, or_297_nl, fsm_output(0));
  mux_538_nl <= MUX_s_1_2_2(mux_537_nl, mux_536_nl, fsm_output(4));
  mux_539_nl <= MUX_s_1_2_2(or_301_nl, mux_538_nl, fsm_output(6));
  or_295_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_534_nl <= MUX_s_1_2_2(or_295_nl, or_tmp_253, fsm_output(0));
  or_296_nl <= (fsm_output(4)) OR mux_534_nl;
  mux_535_nl <= MUX_s_1_2_2(or_296_nl, or_tmp_252, fsm_output(6));
  mux_540_nl <= MUX_s_1_2_2(mux_539_nl, mux_535_nl, fsm_output(7));
  nor_693_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_540_nl);
  or_292_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5))
      OR (NOT (fsm_output(1)));
  or_290_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_530_nl <= MUX_s_1_2_2(or_290_nl, or_tmp_259, fsm_output(0));
  or_286_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_529_nl <= MUX_s_1_2_2(or_tmp_258, or_286_nl, fsm_output(0));
  mux_531_nl <= MUX_s_1_2_2(mux_530_nl, mux_529_nl, fsm_output(4));
  mux_532_nl <= MUX_s_1_2_2(or_292_nl, mux_531_nl, fsm_output(6));
  nand_8_nl <= NOT((fsm_output(7)) AND (NOT mux_532_nl));
  or_283_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_527_nl <= MUX_s_1_2_2(or_283_nl, or_tmp_253, fsm_output(0));
  or_284_nl <= (fsm_output(4)) OR mux_527_nl;
  mux_528_nl <= MUX_s_1_2_2(or_284_nl, or_tmp_252, fsm_output(6));
  or_285_nl <= (fsm_output(7)) OR mux_528_nl;
  mux_533_nl <= MUX_s_1_2_2(nand_8_nl, or_285_nl, fsm_output(8));
  nor_694_nl <= NOT((fsm_output(9)) OR mux_533_nl);
  mux_541_nl <= MUX_s_1_2_2(nor_693_nl, nor_694_nl, fsm_output(3));
  vec_rsc_0_0_i_we_d_pff <= MUX_s_1_2_2(mux_556_nl, mux_541_nl, fsm_output(2));
  nor_678_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_368_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR not_tmp_133;
  or_369_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_372_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_371_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_583_nl <= MUX_s_1_2_2(or_371_nl, or_369_cse, fsm_output(0));
  mux_584_nl <= MUX_s_1_2_2(or_372_nl, mux_583_nl, fsm_output(6));
  or_366_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_581_nl <= MUX_s_1_2_2(or_368_cse, or_366_nl, fsm_output(0));
  or_365_nl <= (VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_363_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_580_nl <= MUX_s_1_2_2(or_365_nl, or_363_nl, fsm_output(0));
  mux_582_nl <= MUX_s_1_2_2(mux_581_nl, mux_580_nl, fsm_output(6));
  mux_585_nl <= MUX_s_1_2_2(mux_584_nl, mux_582_nl, fsm_output(1));
  nor_669_nl <= NOT((fsm_output(3)) OR mux_585_nl);
  or_361_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_359_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_577_nl <= MUX_s_1_2_2(or_361_nl, or_359_nl, fsm_output(0));
  or_358_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_578_nl <= MUX_s_1_2_2(mux_577_nl, or_358_nl, fsm_output(6));
  nor_670_nl <= NOT((fsm_output(1)) OR mux_578_nl);
  nor_671_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  mux_579_nl <= MUX_s_1_2_2(nor_670_nl, nor_671_nl, fsm_output(3));
  mux_586_nl <= MUX_s_1_2_2(nor_669_nl, mux_579_nl, fsm_output(2));
  nor_672_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_673_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_674_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_675_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR not_tmp_133);
  mux_573_nl <= MUX_s_1_2_2(nor_674_nl, nor_675_nl, fsm_output(0));
  mux_574_nl <= MUX_s_1_2_2(nor_673_nl, mux_573_nl, fsm_output(6));
  and_342_nl <= (fsm_output(1)) AND mux_574_nl;
  mux_575_nl <= MUX_s_1_2_2(nor_672_nl, and_342_nl, fsm_output(3));
  nor_676_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_677_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_570_nl <= MUX_s_1_2_2(nor_676_nl, nor_677_nl, fsm_output(0));
  nor_679_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_569_nl <= MUX_s_1_2_2(nor_678_cse, nor_679_nl, fsm_output(0));
  mux_571_nl <= MUX_s_1_2_2(mux_570_nl, mux_569_nl, fsm_output(6));
  nor_680_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_681_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_567_nl <= MUX_s_1_2_2(nor_680_nl, nor_681_nl, fsm_output(0));
  nor_682_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_568_nl <= MUX_s_1_2_2(mux_567_nl, nor_682_nl, fsm_output(6));
  mux_572_nl <= MUX_s_1_2_2(mux_571_nl, mux_568_nl, fsm_output(1));
  and_343_nl <= (fsm_output(3)) AND mux_572_nl;
  mux_576_nl <= MUX_s_1_2_2(mux_575_nl, and_343_nl, fsm_output(2));
  mux_587_nl <= MUX_s_1_2_2(mux_586_nl, mux_576_nl, fsm_output(8));
  nor_685_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_563_nl <= MUX_s_1_2_2(nor_678_cse, nor_685_nl, fsm_output(0));
  nor_686_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_687_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_562_nl <= MUX_s_1_2_2(nor_686_nl, nor_687_nl, fsm_output(0));
  mux_564_nl <= MUX_s_1_2_2(mux_563_nl, mux_562_nl, fsm_output(6));
  nor_688_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_565_nl <= MUX_s_1_2_2(mux_564_nl, nor_688_nl, fsm_output(1));
  nand_11_nl <= NOT((fsm_output(3)) AND mux_565_nl);
  or_328_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_326_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_559_nl <= MUX_s_1_2_2(or_326_nl, or_368_cse, fsm_output(0));
  or_322_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_558_nl <= MUX_s_1_2_2(or_369_cse, or_322_nl, fsm_output(0));
  mux_560_nl <= MUX_s_1_2_2(mux_559_nl, mux_558_nl, fsm_output(6));
  mux_561_nl <= MUX_s_1_2_2(or_328_nl, mux_560_nl, fsm_output(1));
  or_329_nl <= (fsm_output(3)) OR mux_561_nl;
  mux_566_nl <= MUX_s_1_2_2(nand_11_nl, or_329_nl, fsm_output(2));
  nor_683_nl <= NOT((fsm_output(8)) OR mux_566_nl);
  vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_587_nl, nor_683_nl,
      fsm_output(9));
  or_413_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(1)) OR (fsm_output(5));
  mux_614_nl <= MUX_s_1_2_2(or_tmp_353, or_413_nl, fsm_output(0));
  or_412_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_613_nl <= MUX_s_1_2_2(or_412_nl, or_tmp_346, fsm_output(0));
  mux_615_nl <= MUX_s_1_2_2(mux_614_nl, mux_613_nl, fsm_output(4));
  nor_661_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(6))) OR mux_615_nl);
  or_410_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_9_0(0)))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  or_409_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_610_nl <= MUX_s_1_2_2(or_409_nl, or_tmp_353, fsm_output(0));
  or_408_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_609_nl <= MUX_s_1_2_2(or_tmp_352, or_408_nl, fsm_output(0));
  mux_611_nl <= MUX_s_1_2_2(mux_610_nl, mux_609_nl, fsm_output(4));
  mux_612_nl <= MUX_s_1_2_2(or_410_nl, mux_611_nl, fsm_output(6));
  and_341_nl <= (fsm_output(9)) AND (NOT mux_612_nl);
  mux_616_nl <= MUX_s_1_2_2(nor_661_nl, and_341_nl, fsm_output(2));
  or_405_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_608_nl <= MUX_s_1_2_2(or_405_nl, or_tmp_353, fsm_output(0));
  nor_662_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR
      (fsm_output(4)) OR mux_608_nl);
  mux_617_nl <= MUX_s_1_2_2(mux_616_nl, nor_662_nl, fsm_output(8));
  or_402_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(1))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"));
  or_401_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_606_nl <= MUX_s_1_2_2(or_402_nl, or_401_nl, fsm_output(9));
  or_399_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_604_nl <= MUX_s_1_2_2(or_399_nl, or_tmp_346, fsm_output(0));
  or_400_nl <= (fsm_output(4)) OR mux_604_nl;
  mux_605_nl <= MUX_s_1_2_2(or_400_nl, or_tmp_362, fsm_output(6));
  nand_14_nl <= NOT((fsm_output(9)) AND (NOT mux_605_nl));
  mux_607_nl <= MUX_s_1_2_2(mux_606_nl, nand_14_nl, fsm_output(2));
  nor_663_nl <= NOT((fsm_output(8)) OR mux_607_nl);
  mux_618_nl <= MUX_s_1_2_2(mux_617_nl, nor_663_nl, fsm_output(7));
  nor_664_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR
      (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")));
  nor_665_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("000")) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(1)))
      OR (fsm_output(5)));
  or_393_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_599_nl <= MUX_s_1_2_2(or_393_nl, or_tmp_346, fsm_output(0));
  or_394_nl <= (fsm_output(4)) OR mux_599_nl;
  mux_600_nl <= MUX_s_1_2_2(or_394_nl, or_tmp_362, fsm_output(6));
  nor_666_nl <= NOT((fsm_output(9)) OR mux_600_nl);
  mux_601_nl <= MUX_s_1_2_2(nor_665_nl, nor_666_nl, fsm_output(2));
  mux_602_nl <= MUX_s_1_2_2(nor_664_nl, mux_601_nl, fsm_output(8));
  or_389_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT
      (fsm_output(1))) OR (fsm_output(5));
  or_388_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_595_nl <= MUX_s_1_2_2(or_388_nl, or_tmp_353, fsm_output(0));
  or_387_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_594_nl <= MUX_s_1_2_2(or_tmp_352, or_387_nl, fsm_output(0));
  mux_596_nl <= MUX_s_1_2_2(mux_595_nl, mux_594_nl, fsm_output(4));
  mux_597_nl <= MUX_s_1_2_2(or_389_nl, mux_596_nl, fsm_output(6));
  nor_667_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(9)) OR mux_597_nl);
  or_383_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_591_nl <= MUX_s_1_2_2(or_383_nl, or_tmp_353, fsm_output(0));
  or_380_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_590_nl <= MUX_s_1_2_2(or_tmp_352, or_380_nl, fsm_output(0));
  mux_592_nl <= MUX_s_1_2_2(mux_591_nl, mux_590_nl, fsm_output(4));
  or_377_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_589_nl <= MUX_s_1_2_2(or_377_nl, or_tmp_346, fsm_output(0));
  or_378_nl <= (fsm_output(4)) OR mux_589_nl;
  mux_593_nl <= MUX_s_1_2_2(mux_592_nl, or_378_nl, fsm_output(6));
  nor_668_nl <= NOT((fsm_output(2)) OR (fsm_output(9)) OR mux_593_nl);
  mux_598_nl <= MUX_s_1_2_2(nor_667_nl, nor_668_nl, fsm_output(8));
  mux_603_nl <= MUX_s_1_2_2(mux_602_nl, mux_598_nl, fsm_output(7));
  vec_rsc_0_1_i_we_d_pff <= MUX_s_1_2_2(mux_618_nl, mux_603_nl, fsm_output(3));
  nor_650_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_462_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_465_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_464_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_645_nl <= MUX_s_1_2_2(or_464_nl, or_462_cse, fsm_output(0));
  mux_646_nl <= MUX_s_1_2_2(or_465_nl, mux_645_nl, fsm_output(6));
  or_461_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")) OR
      nand_308_cse;
  or_459_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_643_nl <= MUX_s_1_2_2(or_461_nl, or_459_nl, fsm_output(0));
  or_458_nl <= (NOT (VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_456_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_642_nl <= MUX_s_1_2_2(or_458_nl, or_456_nl, fsm_output(0));
  mux_644_nl <= MUX_s_1_2_2(mux_643_nl, mux_642_nl, fsm_output(6));
  mux_647_nl <= MUX_s_1_2_2(mux_646_nl, mux_644_nl, fsm_output(1));
  nor_641_nl <= NOT((fsm_output(3)) OR mux_647_nl);
  or_454_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_452_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR
      (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_639_nl <= MUX_s_1_2_2(or_454_nl, or_452_nl, fsm_output(0));
  or_451_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_640_nl <= MUX_s_1_2_2(mux_639_nl, or_451_nl, fsm_output(6));
  nor_642_nl <= NOT((fsm_output(1)) OR mux_640_nl);
  nor_643_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  mux_641_nl <= MUX_s_1_2_2(nor_642_nl, nor_643_nl, fsm_output(3));
  mux_648_nl <= MUX_s_1_2_2(nor_641_nl, mux_641_nl, fsm_output(2));
  nor_644_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_645_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_646_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_647_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR not_tmp_133);
  mux_635_nl <= MUX_s_1_2_2(nor_646_nl, nor_647_nl, fsm_output(0));
  mux_636_nl <= MUX_s_1_2_2(nor_645_nl, mux_635_nl, fsm_output(6));
  and_339_nl <= (fsm_output(1)) AND mux_636_nl;
  mux_637_nl <= MUX_s_1_2_2(nor_644_nl, and_339_nl, fsm_output(3));
  nor_648_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_649_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_632_nl <= MUX_s_1_2_2(nor_648_nl, nor_649_nl, fsm_output(0));
  nor_651_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_631_nl <= MUX_s_1_2_2(nor_650_cse, nor_651_nl, fsm_output(0));
  mux_633_nl <= MUX_s_1_2_2(mux_632_nl, mux_631_nl, fsm_output(6));
  nor_652_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_653_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_629_nl <= MUX_s_1_2_2(nor_652_nl, nor_653_nl, fsm_output(0));
  nor_654_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_630_nl <= MUX_s_1_2_2(mux_629_nl, nor_654_nl, fsm_output(6));
  mux_634_nl <= MUX_s_1_2_2(mux_633_nl, mux_630_nl, fsm_output(1));
  and_340_nl <= (fsm_output(3)) AND mux_634_nl;
  mux_638_nl <= MUX_s_1_2_2(mux_637_nl, and_340_nl, fsm_output(2));
  mux_649_nl <= MUX_s_1_2_2(mux_648_nl, mux_638_nl, fsm_output(8));
  nor_657_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_625_nl <= MUX_s_1_2_2(nor_650_cse, nor_657_nl, fsm_output(0));
  nor_658_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_659_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_624_nl <= MUX_s_1_2_2(nor_658_nl, nor_659_nl, fsm_output(0));
  mux_626_nl <= MUX_s_1_2_2(mux_625_nl, mux_624_nl, fsm_output(6));
  nor_660_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_627_nl <= MUX_s_1_2_2(mux_626_nl, nor_660_nl, fsm_output(1));
  nand_17_nl <= NOT((fsm_output(3)) AND mux_627_nl);
  or_421_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_419_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_418_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001")) OR
      not_tmp_133;
  mux_621_nl <= MUX_s_1_2_2(or_419_nl, or_418_nl, fsm_output(0));
  or_415_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_620_nl <= MUX_s_1_2_2(or_462_cse, or_415_nl, fsm_output(0));
  mux_622_nl <= MUX_s_1_2_2(mux_621_nl, mux_620_nl, fsm_output(6));
  mux_623_nl <= MUX_s_1_2_2(or_421_nl, mux_622_nl, fsm_output(1));
  or_422_nl <= (fsm_output(3)) OR mux_623_nl;
  mux_628_nl <= MUX_s_1_2_2(nand_17_nl, or_422_nl, fsm_output(2));
  nor_655_nl <= NOT((fsm_output(8)) OR mux_628_nl);
  vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_649_nl, nor_655_nl,
      fsm_output(9));
  or_505_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_676_nl <= MUX_s_1_2_2(or_tmp_445, or_505_nl, fsm_output(0));
  or_504_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_675_nl <= MUX_s_1_2_2(or_504_nl, or_tmp_439, fsm_output(0));
  mux_677_nl <= MUX_s_1_2_2(mux_676_nl, mux_675_nl, fsm_output(4));
  nand_22_nl <= NOT((fsm_output(6)) AND (NOT mux_677_nl));
  or_503_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0010"));
  mux_678_nl <= MUX_s_1_2_2(nand_22_nl, or_503_nl, fsm_output(7));
  nor_635_nl <= NOT((fsm_output(8)) OR mux_678_nl);
  nor_636_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT
      (fsm_output(1))));
  or_499_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_673_nl <= MUX_s_1_2_2(or_499_nl, or_tmp_445, fsm_output(0));
  nor_637_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_673_nl);
  mux_674_nl <= MUX_s_1_2_2(nor_636_nl, nor_637_nl, fsm_output(8));
  mux_679_nl <= MUX_s_1_2_2(nor_635_nl, mux_674_nl, fsm_output(9));
  or_496_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_494_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_668_nl <= MUX_s_1_2_2(or_494_nl, or_tmp_445, fsm_output(0));
  or_492_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_667_nl <= MUX_s_1_2_2(or_tmp_444, or_492_nl, fsm_output(0));
  mux_669_nl <= MUX_s_1_2_2(mux_668_nl, mux_667_nl, fsm_output(4));
  or_490_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_666_nl <= MUX_s_1_2_2(or_490_nl, or_tmp_439, fsm_output(0));
  or_491_nl <= (fsm_output(4)) OR mux_666_nl;
  mux_670_nl <= MUX_s_1_2_2(mux_669_nl, or_491_nl, fsm_output(6));
  mux_671_nl <= MUX_s_1_2_2(or_496_nl, mux_670_nl, fsm_output(7));
  and_338_nl <= (fsm_output(8)) AND (NOT mux_671_nl);
  nor_638_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")));
  mux_672_nl <= MUX_s_1_2_2(and_338_nl, nor_638_nl, fsm_output(9));
  mux_680_nl <= MUX_s_1_2_2(mux_679_nl, mux_672_nl, fsm_output(3));
  or_487_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_485_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_661_nl <= MUX_s_1_2_2(or_485_nl, or_tmp_445, fsm_output(0));
  or_483_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_660_nl <= MUX_s_1_2_2(or_tmp_444, or_483_nl, fsm_output(0));
  mux_662_nl <= MUX_s_1_2_2(mux_661_nl, mux_660_nl, fsm_output(4));
  mux_663_nl <= MUX_s_1_2_2(or_487_nl, mux_662_nl, fsm_output(6));
  or_481_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_658_nl <= MUX_s_1_2_2(or_481_nl, or_tmp_439, fsm_output(0));
  or_482_nl <= (fsm_output(4)) OR mux_658_nl;
  mux_659_nl <= MUX_s_1_2_2(or_482_nl, or_tmp_438, fsm_output(6));
  mux_664_nl <= MUX_s_1_2_2(mux_663_nl, mux_659_nl, fsm_output(7));
  nor_639_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_664_nl);
  or_478_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5))
      OR (NOT (fsm_output(1)));
  or_476_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_654_nl <= MUX_s_1_2_2(or_476_nl, or_tmp_445, fsm_output(0));
  or_472_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_653_nl <= MUX_s_1_2_2(or_tmp_444, or_472_nl, fsm_output(0));
  mux_655_nl <= MUX_s_1_2_2(mux_654_nl, mux_653_nl, fsm_output(4));
  mux_656_nl <= MUX_s_1_2_2(or_478_nl, mux_655_nl, fsm_output(6));
  nand_20_nl <= NOT((fsm_output(7)) AND (NOT mux_656_nl));
  or_469_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_651_nl <= MUX_s_1_2_2(or_469_nl, or_tmp_439, fsm_output(0));
  or_470_nl <= (fsm_output(4)) OR mux_651_nl;
  mux_652_nl <= MUX_s_1_2_2(or_470_nl, or_tmp_438, fsm_output(6));
  or_471_nl <= (fsm_output(7)) OR mux_652_nl;
  mux_657_nl <= MUX_s_1_2_2(nand_20_nl, or_471_nl, fsm_output(8));
  nor_640_nl <= NOT((fsm_output(9)) OR mux_657_nl);
  mux_665_nl <= MUX_s_1_2_2(nor_639_nl, nor_640_nl, fsm_output(3));
  vec_rsc_0_2_i_we_d_pff <= MUX_s_1_2_2(mux_680_nl, mux_665_nl, fsm_output(2));
  nor_624_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_554_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR not_tmp_133;
  or_555_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_558_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_557_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_707_nl <= MUX_s_1_2_2(or_557_nl, or_555_cse, fsm_output(0));
  mux_708_nl <= MUX_s_1_2_2(or_558_nl, mux_707_nl, fsm_output(6));
  or_552_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_705_nl <= MUX_s_1_2_2(or_554_cse, or_552_nl, fsm_output(0));
  or_551_nl <= (VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_549_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_704_nl <= MUX_s_1_2_2(or_551_nl, or_549_nl, fsm_output(0));
  mux_706_nl <= MUX_s_1_2_2(mux_705_nl, mux_704_nl, fsm_output(6));
  mux_709_nl <= MUX_s_1_2_2(mux_708_nl, mux_706_nl, fsm_output(1));
  nor_615_nl <= NOT((fsm_output(3)) OR mux_709_nl);
  or_547_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_545_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR
      (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_701_nl <= MUX_s_1_2_2(or_547_nl, or_545_nl, fsm_output(0));
  or_544_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_702_nl <= MUX_s_1_2_2(mux_701_nl, or_544_nl, fsm_output(6));
  nor_616_nl <= NOT((fsm_output(1)) OR mux_702_nl);
  nor_617_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  mux_703_nl <= MUX_s_1_2_2(nor_616_nl, nor_617_nl, fsm_output(3));
  mux_710_nl <= MUX_s_1_2_2(nor_615_nl, mux_703_nl, fsm_output(2));
  nor_618_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0010")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_619_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_620_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_621_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR not_tmp_133);
  mux_697_nl <= MUX_s_1_2_2(nor_620_nl, nor_621_nl, fsm_output(0));
  mux_698_nl <= MUX_s_1_2_2(nor_619_nl, mux_697_nl, fsm_output(6));
  and_336_nl <= (fsm_output(1)) AND mux_698_nl;
  mux_699_nl <= MUX_s_1_2_2(nor_618_nl, and_336_nl, fsm_output(3));
  nor_622_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_623_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_694_nl <= MUX_s_1_2_2(nor_622_nl, nor_623_nl, fsm_output(0));
  nor_625_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_693_nl <= MUX_s_1_2_2(nor_624_cse, nor_625_nl, fsm_output(0));
  mux_695_nl <= MUX_s_1_2_2(mux_694_nl, mux_693_nl, fsm_output(6));
  nor_626_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_627_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_691_nl <= MUX_s_1_2_2(nor_626_nl, nor_627_nl, fsm_output(0));
  nor_628_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_692_nl <= MUX_s_1_2_2(mux_691_nl, nor_628_nl, fsm_output(6));
  mux_696_nl <= MUX_s_1_2_2(mux_695_nl, mux_692_nl, fsm_output(1));
  and_337_nl <= (fsm_output(3)) AND mux_696_nl;
  mux_700_nl <= MUX_s_1_2_2(mux_699_nl, and_337_nl, fsm_output(2));
  mux_711_nl <= MUX_s_1_2_2(mux_710_nl, mux_700_nl, fsm_output(8));
  nor_631_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_687_nl <= MUX_s_1_2_2(nor_624_cse, nor_631_nl, fsm_output(0));
  nor_632_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_633_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_686_nl <= MUX_s_1_2_2(nor_632_nl, nor_633_nl, fsm_output(0));
  mux_688_nl <= MUX_s_1_2_2(mux_687_nl, mux_686_nl, fsm_output(6));
  nor_634_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_689_nl <= MUX_s_1_2_2(mux_688_nl, nor_634_nl, fsm_output(1));
  nand_23_nl <= NOT((fsm_output(3)) AND mux_689_nl);
  or_514_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_512_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_683_nl <= MUX_s_1_2_2(or_512_nl, or_554_cse, fsm_output(0));
  or_508_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_682_nl <= MUX_s_1_2_2(or_555_cse, or_508_nl, fsm_output(0));
  mux_684_nl <= MUX_s_1_2_2(mux_683_nl, mux_682_nl, fsm_output(6));
  mux_685_nl <= MUX_s_1_2_2(or_514_nl, mux_684_nl, fsm_output(1));
  or_515_nl <= (fsm_output(3)) OR mux_685_nl;
  mux_690_nl <= MUX_s_1_2_2(nand_23_nl, or_515_nl, fsm_output(2));
  nor_629_nl <= NOT((fsm_output(8)) OR mux_690_nl);
  vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_711_nl, nor_629_nl,
      fsm_output(9));
  or_598_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_738_nl <= MUX_s_1_2_2(or_tmp_538, or_598_nl, fsm_output(0));
  or_597_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_737_nl <= MUX_s_1_2_2(or_597_nl, or_tmp_532, fsm_output(0));
  mux_739_nl <= MUX_s_1_2_2(mux_738_nl, mux_737_nl, fsm_output(4));
  nand_28_nl <= NOT((fsm_output(6)) AND (NOT mux_739_nl));
  or_596_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0011"));
  mux_740_nl <= MUX_s_1_2_2(nand_28_nl, or_596_nl, fsm_output(7));
  nor_609_nl <= NOT((fsm_output(8)) OR mux_740_nl);
  and_439_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("001"))
      AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT (fsm_output(5))) AND (fsm_output(1));
  or_592_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_735_nl <= MUX_s_1_2_2(or_592_nl, or_tmp_538, fsm_output(0));
  nor_611_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_735_nl);
  mux_736_nl <= MUX_s_1_2_2(and_439_nl, nor_611_nl, fsm_output(8));
  mux_741_nl <= MUX_s_1_2_2(nor_609_nl, mux_736_nl, fsm_output(9));
  or_589_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_587_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_730_nl <= MUX_s_1_2_2(or_587_nl, or_tmp_538, fsm_output(0));
  or_585_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_729_nl <= MUX_s_1_2_2(or_tmp_537, or_585_nl, fsm_output(0));
  mux_731_nl <= MUX_s_1_2_2(mux_730_nl, mux_729_nl, fsm_output(4));
  or_583_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_728_nl <= MUX_s_1_2_2(or_583_nl, or_tmp_532, fsm_output(0));
  or_584_nl <= (fsm_output(4)) OR mux_728_nl;
  mux_732_nl <= MUX_s_1_2_2(mux_731_nl, or_584_nl, fsm_output(6));
  mux_733_nl <= MUX_s_1_2_2(or_589_nl, mux_732_nl, fsm_output(7));
  and_335_nl <= (fsm_output(8)) AND (NOT mux_733_nl);
  nor_612_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")));
  mux_734_nl <= MUX_s_1_2_2(and_335_nl, nor_612_nl, fsm_output(9));
  mux_742_nl <= MUX_s_1_2_2(mux_741_nl, mux_734_nl, fsm_output(3));
  or_580_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_9_0(0)))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_578_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_723_nl <= MUX_s_1_2_2(or_578_nl, or_tmp_538, fsm_output(0));
  or_576_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_722_nl <= MUX_s_1_2_2(or_tmp_537, or_576_nl, fsm_output(0));
  mux_724_nl <= MUX_s_1_2_2(mux_723_nl, mux_722_nl, fsm_output(4));
  mux_725_nl <= MUX_s_1_2_2(or_580_nl, mux_724_nl, fsm_output(6));
  or_574_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_720_nl <= MUX_s_1_2_2(or_574_nl, or_tmp_532, fsm_output(0));
  or_575_nl <= (fsm_output(4)) OR mux_720_nl;
  mux_721_nl <= MUX_s_1_2_2(or_575_nl, or_tmp_531, fsm_output(6));
  mux_726_nl <= MUX_s_1_2_2(mux_725_nl, mux_721_nl, fsm_output(7));
  nor_613_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_726_nl);
  or_571_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (fsm_output(5))
      OR (NOT (fsm_output(1)));
  or_569_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_716_nl <= MUX_s_1_2_2(or_569_nl, or_tmp_538, fsm_output(0));
  or_565_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_715_nl <= MUX_s_1_2_2(or_tmp_537, or_565_nl, fsm_output(0));
  mux_717_nl <= MUX_s_1_2_2(mux_716_nl, mux_715_nl, fsm_output(4));
  mux_718_nl <= MUX_s_1_2_2(or_571_nl, mux_717_nl, fsm_output(6));
  nand_26_nl <= NOT((fsm_output(7)) AND (NOT mux_718_nl));
  or_562_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_713_nl <= MUX_s_1_2_2(or_562_nl, or_tmp_532, fsm_output(0));
  or_563_nl <= (fsm_output(4)) OR mux_713_nl;
  mux_714_nl <= MUX_s_1_2_2(or_563_nl, or_tmp_531, fsm_output(6));
  or_564_nl <= (fsm_output(7)) OR mux_714_nl;
  mux_719_nl <= MUX_s_1_2_2(nand_26_nl, or_564_nl, fsm_output(8));
  nor_614_nl <= NOT((fsm_output(9)) OR mux_719_nl);
  mux_727_nl <= MUX_s_1_2_2(nor_613_nl, nor_614_nl, fsm_output(3));
  vec_rsc_0_3_i_we_d_pff <= MUX_s_1_2_2(mux_742_nl, mux_727_nl, fsm_output(2));
  nor_598_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_648_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_651_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_650_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_769_nl <= MUX_s_1_2_2(or_650_nl, or_648_cse, fsm_output(0));
  mux_770_nl <= MUX_s_1_2_2(or_651_nl, mux_769_nl, fsm_output(6));
  or_647_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("001")) OR
      nand_308_cse;
  or_645_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_767_nl <= MUX_s_1_2_2(or_647_nl, or_645_nl, fsm_output(0));
  or_644_nl <= (NOT (VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_642_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_766_nl <= MUX_s_1_2_2(or_644_nl, or_642_nl, fsm_output(0));
  mux_768_nl <= MUX_s_1_2_2(mux_767_nl, mux_766_nl, fsm_output(6));
  mux_771_nl <= MUX_s_1_2_2(mux_770_nl, mux_768_nl, fsm_output(1));
  nor_589_nl <= NOT((fsm_output(3)) OR mux_771_nl);
  or_640_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_638_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR
      (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_763_nl <= MUX_s_1_2_2(or_640_nl, or_638_nl, fsm_output(0));
  or_637_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_764_nl <= MUX_s_1_2_2(mux_763_nl, or_637_nl, fsm_output(6));
  nor_590_nl <= NOT((fsm_output(1)) OR mux_764_nl);
  nor_591_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0011"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_765_nl <= MUX_s_1_2_2(nor_590_nl, nor_591_nl, fsm_output(3));
  mux_772_nl <= MUX_s_1_2_2(nor_589_nl, mux_765_nl, fsm_output(2));
  nor_592_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_593_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_594_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_595_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR not_tmp_133);
  mux_759_nl <= MUX_s_1_2_2(nor_594_nl, nor_595_nl, fsm_output(0));
  mux_760_nl <= MUX_s_1_2_2(nor_593_nl, mux_759_nl, fsm_output(6));
  and_333_nl <= (fsm_output(1)) AND mux_760_nl;
  mux_761_nl <= MUX_s_1_2_2(nor_592_nl, and_333_nl, fsm_output(3));
  nor_596_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_597_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_756_nl <= MUX_s_1_2_2(nor_596_nl, nor_597_nl, fsm_output(0));
  nor_599_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_755_nl <= MUX_s_1_2_2(nor_598_cse, nor_599_nl, fsm_output(0));
  mux_757_nl <= MUX_s_1_2_2(mux_756_nl, mux_755_nl, fsm_output(6));
  nor_600_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_601_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_753_nl <= MUX_s_1_2_2(nor_600_nl, nor_601_nl, fsm_output(0));
  nor_602_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_754_nl <= MUX_s_1_2_2(mux_753_nl, nor_602_nl, fsm_output(6));
  mux_758_nl <= MUX_s_1_2_2(mux_757_nl, mux_754_nl, fsm_output(1));
  and_334_nl <= (fsm_output(3)) AND mux_758_nl;
  mux_762_nl <= MUX_s_1_2_2(mux_761_nl, and_334_nl, fsm_output(2));
  mux_773_nl <= MUX_s_1_2_2(mux_772_nl, mux_762_nl, fsm_output(8));
  nor_605_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_749_nl <= MUX_s_1_2_2(nor_598_cse, nor_605_nl, fsm_output(0));
  nor_606_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_607_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_748_nl <= MUX_s_1_2_2(nor_606_nl, nor_607_nl, fsm_output(0));
  mux_750_nl <= MUX_s_1_2_2(mux_749_nl, mux_748_nl, fsm_output(6));
  nor_608_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_751_nl <= MUX_s_1_2_2(mux_750_nl, nor_608_nl, fsm_output(1));
  nand_29_nl <= NOT((fsm_output(3)) AND mux_751_nl);
  or_607_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_605_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_604_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011")) OR
      not_tmp_133;
  mux_745_nl <= MUX_s_1_2_2(or_605_nl, or_604_nl, fsm_output(0));
  or_601_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_744_nl <= MUX_s_1_2_2(or_648_cse, or_601_nl, fsm_output(0));
  mux_746_nl <= MUX_s_1_2_2(mux_745_nl, mux_744_nl, fsm_output(6));
  mux_747_nl <= MUX_s_1_2_2(or_607_nl, mux_746_nl, fsm_output(1));
  or_608_nl <= (fsm_output(3)) OR mux_747_nl;
  mux_752_nl <= MUX_s_1_2_2(nand_29_nl, or_608_nl, fsm_output(2));
  nor_603_nl <= NOT((fsm_output(8)) OR mux_752_nl);
  vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_773_nl, nor_603_nl,
      fsm_output(9));
  or_691_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_800_nl <= MUX_s_1_2_2(or_tmp_631, or_691_nl, fsm_output(0));
  or_690_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_799_nl <= MUX_s_1_2_2(or_690_nl, or_tmp_625, fsm_output(0));
  mux_801_nl <= MUX_s_1_2_2(mux_800_nl, mux_799_nl, fsm_output(4));
  nand_34_nl <= NOT((fsm_output(6)) AND (NOT mux_801_nl));
  or_689_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0100"));
  mux_802_nl <= MUX_s_1_2_2(nand_34_nl, or_689_nl, fsm_output(7));
  nor_583_nl <= NOT((fsm_output(8)) OR mux_802_nl);
  nor_584_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT
      (fsm_output(1))));
  or_685_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_797_nl <= MUX_s_1_2_2(or_685_nl, or_tmp_631, fsm_output(0));
  nor_585_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_797_nl);
  mux_798_nl <= MUX_s_1_2_2(nor_584_nl, nor_585_nl, fsm_output(8));
  mux_803_nl <= MUX_s_1_2_2(nor_583_nl, mux_798_nl, fsm_output(9));
  or_682_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_680_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_792_nl <= MUX_s_1_2_2(or_680_nl, or_tmp_631, fsm_output(0));
  or_678_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_791_nl <= MUX_s_1_2_2(or_tmp_630, or_678_nl, fsm_output(0));
  mux_793_nl <= MUX_s_1_2_2(mux_792_nl, mux_791_nl, fsm_output(4));
  or_676_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_790_nl <= MUX_s_1_2_2(or_676_nl, or_tmp_625, fsm_output(0));
  or_677_nl <= (fsm_output(4)) OR mux_790_nl;
  mux_794_nl <= MUX_s_1_2_2(mux_793_nl, or_677_nl, fsm_output(6));
  mux_795_nl <= MUX_s_1_2_2(or_682_nl, mux_794_nl, fsm_output(7));
  and_332_nl <= (fsm_output(8)) AND (NOT mux_795_nl);
  nor_586_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")));
  mux_796_nl <= MUX_s_1_2_2(and_332_nl, nor_586_nl, fsm_output(9));
  mux_804_nl <= MUX_s_1_2_2(mux_803_nl, mux_796_nl, fsm_output(3));
  or_673_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_671_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_785_nl <= MUX_s_1_2_2(or_671_nl, or_tmp_631, fsm_output(0));
  or_669_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_784_nl <= MUX_s_1_2_2(or_tmp_630, or_669_nl, fsm_output(0));
  mux_786_nl <= MUX_s_1_2_2(mux_785_nl, mux_784_nl, fsm_output(4));
  mux_787_nl <= MUX_s_1_2_2(or_673_nl, mux_786_nl, fsm_output(6));
  or_667_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_782_nl <= MUX_s_1_2_2(or_667_nl, or_tmp_625, fsm_output(0));
  or_668_nl <= (fsm_output(4)) OR mux_782_nl;
  mux_783_nl <= MUX_s_1_2_2(or_668_nl, or_tmp_624, fsm_output(6));
  mux_788_nl <= MUX_s_1_2_2(mux_787_nl, mux_783_nl, fsm_output(7));
  nor_587_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_788_nl);
  or_664_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5))
      OR (NOT (fsm_output(1)));
  or_662_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_778_nl <= MUX_s_1_2_2(or_662_nl, or_tmp_631, fsm_output(0));
  or_658_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_777_nl <= MUX_s_1_2_2(or_tmp_630, or_658_nl, fsm_output(0));
  mux_779_nl <= MUX_s_1_2_2(mux_778_nl, mux_777_nl, fsm_output(4));
  mux_780_nl <= MUX_s_1_2_2(or_664_nl, mux_779_nl, fsm_output(6));
  nand_32_nl <= NOT((fsm_output(7)) AND (NOT mux_780_nl));
  or_655_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_775_nl <= MUX_s_1_2_2(or_655_nl, or_tmp_625, fsm_output(0));
  or_656_nl <= (fsm_output(4)) OR mux_775_nl;
  mux_776_nl <= MUX_s_1_2_2(or_656_nl, or_tmp_624, fsm_output(6));
  or_657_nl <= (fsm_output(7)) OR mux_776_nl;
  mux_781_nl <= MUX_s_1_2_2(nand_32_nl, or_657_nl, fsm_output(8));
  nor_588_nl <= NOT((fsm_output(9)) OR mux_781_nl);
  mux_789_nl <= MUX_s_1_2_2(nor_587_nl, nor_588_nl, fsm_output(3));
  vec_rsc_0_4_i_we_d_pff <= MUX_s_1_2_2(mux_804_nl, mux_789_nl, fsm_output(2));
  nor_572_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_740_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR not_tmp_133;
  or_741_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_744_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_743_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_831_nl <= MUX_s_1_2_2(or_743_nl, or_741_cse, fsm_output(0));
  mux_832_nl <= MUX_s_1_2_2(or_744_nl, mux_831_nl, fsm_output(6));
  or_738_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_829_nl <= MUX_s_1_2_2(or_740_cse, or_738_nl, fsm_output(0));
  or_737_nl <= (VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_735_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_828_nl <= MUX_s_1_2_2(or_737_nl, or_735_nl, fsm_output(0));
  mux_830_nl <= MUX_s_1_2_2(mux_829_nl, mux_828_nl, fsm_output(6));
  mux_833_nl <= MUX_s_1_2_2(mux_832_nl, mux_830_nl, fsm_output(1));
  nor_563_nl <= NOT((fsm_output(3)) OR mux_833_nl);
  or_733_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_731_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR
      (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_825_nl <= MUX_s_1_2_2(or_733_nl, or_731_nl, fsm_output(0));
  or_730_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_826_nl <= MUX_s_1_2_2(mux_825_nl, or_730_nl, fsm_output(6));
  nor_564_nl <= NOT((fsm_output(1)) OR mux_826_nl);
  nor_565_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  mux_827_nl <= MUX_s_1_2_2(nor_564_nl, nor_565_nl, fsm_output(3));
  mux_834_nl <= MUX_s_1_2_2(nor_563_nl, mux_827_nl, fsm_output(2));
  nor_566_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0100")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_567_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_568_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_569_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR not_tmp_133);
  mux_821_nl <= MUX_s_1_2_2(nor_568_nl, nor_569_nl, fsm_output(0));
  mux_822_nl <= MUX_s_1_2_2(nor_567_nl, mux_821_nl, fsm_output(6));
  and_330_nl <= (fsm_output(1)) AND mux_822_nl;
  mux_823_nl <= MUX_s_1_2_2(nor_566_nl, and_330_nl, fsm_output(3));
  nor_570_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_571_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_818_nl <= MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output(0));
  nor_573_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_817_nl <= MUX_s_1_2_2(nor_572_cse, nor_573_nl, fsm_output(0));
  mux_819_nl <= MUX_s_1_2_2(mux_818_nl, mux_817_nl, fsm_output(6));
  nor_574_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_575_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_815_nl <= MUX_s_1_2_2(nor_574_nl, nor_575_nl, fsm_output(0));
  nor_576_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_816_nl <= MUX_s_1_2_2(mux_815_nl, nor_576_nl, fsm_output(6));
  mux_820_nl <= MUX_s_1_2_2(mux_819_nl, mux_816_nl, fsm_output(1));
  and_331_nl <= (fsm_output(3)) AND mux_820_nl;
  mux_824_nl <= MUX_s_1_2_2(mux_823_nl, and_331_nl, fsm_output(2));
  mux_835_nl <= MUX_s_1_2_2(mux_834_nl, mux_824_nl, fsm_output(8));
  nor_579_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_811_nl <= MUX_s_1_2_2(nor_572_cse, nor_579_nl, fsm_output(0));
  nor_580_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_581_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_810_nl <= MUX_s_1_2_2(nor_580_nl, nor_581_nl, fsm_output(0));
  mux_812_nl <= MUX_s_1_2_2(mux_811_nl, mux_810_nl, fsm_output(6));
  nor_582_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_813_nl <= MUX_s_1_2_2(mux_812_nl, nor_582_nl, fsm_output(1));
  nand_35_nl <= NOT((fsm_output(3)) AND mux_813_nl);
  or_700_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_698_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_807_nl <= MUX_s_1_2_2(or_698_nl, or_740_cse, fsm_output(0));
  or_694_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_806_nl <= MUX_s_1_2_2(or_741_cse, or_694_nl, fsm_output(0));
  mux_808_nl <= MUX_s_1_2_2(mux_807_nl, mux_806_nl, fsm_output(6));
  mux_809_nl <= MUX_s_1_2_2(or_700_nl, mux_808_nl, fsm_output(1));
  or_701_nl <= (fsm_output(3)) OR mux_809_nl;
  mux_814_nl <= MUX_s_1_2_2(nand_35_nl, or_701_nl, fsm_output(2));
  nor_577_nl <= NOT((fsm_output(8)) OR mux_814_nl);
  vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_835_nl, nor_577_nl,
      fsm_output(9));
  or_785_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(1)) OR (fsm_output(5));
  mux_862_nl <= MUX_s_1_2_2(or_tmp_725, or_785_nl, fsm_output(0));
  or_784_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_861_nl <= MUX_s_1_2_2(or_784_nl, or_tmp_718, fsm_output(0));
  mux_863_nl <= MUX_s_1_2_2(mux_862_nl, mux_861_nl, fsm_output(4));
  nor_555_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(6))) OR mux_863_nl);
  or_782_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_9_0(0)))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  or_781_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_858_nl <= MUX_s_1_2_2(or_781_nl, or_tmp_725, fsm_output(0));
  or_780_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_857_nl <= MUX_s_1_2_2(or_tmp_724, or_780_nl, fsm_output(0));
  mux_859_nl <= MUX_s_1_2_2(mux_858_nl, mux_857_nl, fsm_output(4));
  mux_860_nl <= MUX_s_1_2_2(or_782_nl, mux_859_nl, fsm_output(6));
  and_329_nl <= (fsm_output(9)) AND (NOT mux_860_nl);
  mux_864_nl <= MUX_s_1_2_2(nor_555_nl, and_329_nl, fsm_output(2));
  or_777_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_856_nl <= MUX_s_1_2_2(or_777_nl, or_tmp_725, fsm_output(0));
  nor_556_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR
      (fsm_output(4)) OR mux_856_nl);
  mux_865_nl <= MUX_s_1_2_2(mux_864_nl, nor_556_nl, fsm_output(8));
  or_774_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(1))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"));
  or_773_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_854_nl <= MUX_s_1_2_2(or_774_nl, or_773_nl, fsm_output(9));
  or_771_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_852_nl <= MUX_s_1_2_2(or_771_nl, or_tmp_718, fsm_output(0));
  or_772_nl <= (fsm_output(4)) OR mux_852_nl;
  mux_853_nl <= MUX_s_1_2_2(or_772_nl, or_tmp_734, fsm_output(6));
  nand_38_nl <= NOT((fsm_output(9)) AND (NOT mux_853_nl));
  mux_855_nl <= MUX_s_1_2_2(mux_854_nl, nand_38_nl, fsm_output(2));
  nor_557_nl <= NOT((fsm_output(8)) OR mux_855_nl);
  mux_866_nl <= MUX_s_1_2_2(mux_865_nl, nor_557_nl, fsm_output(7));
  nor_558_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR
      (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")));
  nor_559_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("010")) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(1)))
      OR (fsm_output(5)));
  or_765_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_847_nl <= MUX_s_1_2_2(or_765_nl, or_tmp_718, fsm_output(0));
  or_766_nl <= (fsm_output(4)) OR mux_847_nl;
  mux_848_nl <= MUX_s_1_2_2(or_766_nl, or_tmp_734, fsm_output(6));
  nor_560_nl <= NOT((fsm_output(9)) OR mux_848_nl);
  mux_849_nl <= MUX_s_1_2_2(nor_559_nl, nor_560_nl, fsm_output(2));
  mux_850_nl <= MUX_s_1_2_2(nor_558_nl, mux_849_nl, fsm_output(8));
  or_761_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT
      (fsm_output(1))) OR (fsm_output(5));
  or_760_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_843_nl <= MUX_s_1_2_2(or_760_nl, or_tmp_725, fsm_output(0));
  or_759_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_842_nl <= MUX_s_1_2_2(or_tmp_724, or_759_nl, fsm_output(0));
  mux_844_nl <= MUX_s_1_2_2(mux_843_nl, mux_842_nl, fsm_output(4));
  mux_845_nl <= MUX_s_1_2_2(or_761_nl, mux_844_nl, fsm_output(6));
  nor_561_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(9)) OR mux_845_nl);
  or_755_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_839_nl <= MUX_s_1_2_2(or_755_nl, or_tmp_725, fsm_output(0));
  or_752_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_838_nl <= MUX_s_1_2_2(or_tmp_724, or_752_nl, fsm_output(0));
  mux_840_nl <= MUX_s_1_2_2(mux_839_nl, mux_838_nl, fsm_output(4));
  or_749_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_837_nl <= MUX_s_1_2_2(or_749_nl, or_tmp_718, fsm_output(0));
  or_750_nl <= (fsm_output(4)) OR mux_837_nl;
  mux_841_nl <= MUX_s_1_2_2(mux_840_nl, or_750_nl, fsm_output(6));
  nor_562_nl <= NOT((fsm_output(2)) OR (fsm_output(9)) OR mux_841_nl);
  mux_846_nl <= MUX_s_1_2_2(nor_561_nl, nor_562_nl, fsm_output(8));
  mux_851_nl <= MUX_s_1_2_2(mux_850_nl, mux_846_nl, fsm_output(7));
  vec_rsc_0_5_i_we_d_pff <= MUX_s_1_2_2(mux_866_nl, mux_851_nl, fsm_output(3));
  nor_544_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_834_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_837_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_836_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_893_nl <= MUX_s_1_2_2(or_836_nl, or_834_cse, fsm_output(0));
  mux_894_nl <= MUX_s_1_2_2(or_837_nl, mux_893_nl, fsm_output(6));
  or_833_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("010")) OR
      nand_308_cse;
  or_831_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_891_nl <= MUX_s_1_2_2(or_833_nl, or_831_nl, fsm_output(0));
  or_830_nl <= (NOT (VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_828_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_890_nl <= MUX_s_1_2_2(or_830_nl, or_828_nl, fsm_output(0));
  mux_892_nl <= MUX_s_1_2_2(mux_891_nl, mux_890_nl, fsm_output(6));
  mux_895_nl <= MUX_s_1_2_2(mux_894_nl, mux_892_nl, fsm_output(1));
  nor_535_nl <= NOT((fsm_output(3)) OR mux_895_nl);
  or_826_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_824_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR
      (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_887_nl <= MUX_s_1_2_2(or_826_nl, or_824_nl, fsm_output(0));
  or_823_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_888_nl <= MUX_s_1_2_2(mux_887_nl, or_823_nl, fsm_output(6));
  nor_536_nl <= NOT((fsm_output(1)) OR mux_888_nl);
  nor_537_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0101"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_889_nl <= MUX_s_1_2_2(nor_536_nl, nor_537_nl, fsm_output(3));
  mux_896_nl <= MUX_s_1_2_2(nor_535_nl, mux_889_nl, fsm_output(2));
  nor_538_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_539_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_540_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_541_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR not_tmp_133);
  mux_883_nl <= MUX_s_1_2_2(nor_540_nl, nor_541_nl, fsm_output(0));
  mux_884_nl <= MUX_s_1_2_2(nor_539_nl, mux_883_nl, fsm_output(6));
  and_327_nl <= (fsm_output(1)) AND mux_884_nl;
  mux_885_nl <= MUX_s_1_2_2(nor_538_nl, and_327_nl, fsm_output(3));
  nor_542_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_543_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_880_nl <= MUX_s_1_2_2(nor_542_nl, nor_543_nl, fsm_output(0));
  nor_545_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_879_nl <= MUX_s_1_2_2(nor_544_cse, nor_545_nl, fsm_output(0));
  mux_881_nl <= MUX_s_1_2_2(mux_880_nl, mux_879_nl, fsm_output(6));
  nor_546_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_547_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_877_nl <= MUX_s_1_2_2(nor_546_nl, nor_547_nl, fsm_output(0));
  nor_548_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_878_nl <= MUX_s_1_2_2(mux_877_nl, nor_548_nl, fsm_output(6));
  mux_882_nl <= MUX_s_1_2_2(mux_881_nl, mux_878_nl, fsm_output(1));
  and_328_nl <= (fsm_output(3)) AND mux_882_nl;
  mux_886_nl <= MUX_s_1_2_2(mux_885_nl, and_328_nl, fsm_output(2));
  mux_897_nl <= MUX_s_1_2_2(mux_896_nl, mux_886_nl, fsm_output(8));
  nor_551_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_873_nl <= MUX_s_1_2_2(nor_544_cse, nor_551_nl, fsm_output(0));
  nor_552_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_553_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_872_nl <= MUX_s_1_2_2(nor_552_nl, nor_553_nl, fsm_output(0));
  mux_874_nl <= MUX_s_1_2_2(mux_873_nl, mux_872_nl, fsm_output(6));
  nor_554_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_875_nl <= MUX_s_1_2_2(mux_874_nl, nor_554_nl, fsm_output(1));
  nand_41_nl <= NOT((fsm_output(3)) AND mux_875_nl);
  or_793_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_791_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_790_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101")) OR
      not_tmp_133;
  mux_869_nl <= MUX_s_1_2_2(or_791_nl, or_790_nl, fsm_output(0));
  or_787_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_868_nl <= MUX_s_1_2_2(or_834_cse, or_787_nl, fsm_output(0));
  mux_870_nl <= MUX_s_1_2_2(mux_869_nl, mux_868_nl, fsm_output(6));
  mux_871_nl <= MUX_s_1_2_2(or_793_nl, mux_870_nl, fsm_output(1));
  or_794_nl <= (fsm_output(3)) OR mux_871_nl;
  mux_876_nl <= MUX_s_1_2_2(nand_41_nl, or_794_nl, fsm_output(2));
  nor_549_nl <= NOT((fsm_output(8)) OR mux_876_nl);
  vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_897_nl, nor_549_nl,
      fsm_output(9));
  or_877_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_924_nl <= MUX_s_1_2_2(or_tmp_817, or_877_nl, fsm_output(0));
  or_876_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_923_nl <= MUX_s_1_2_2(or_876_nl, or_tmp_811, fsm_output(0));
  mux_925_nl <= MUX_s_1_2_2(mux_924_nl, mux_923_nl, fsm_output(4));
  nand_46_nl <= NOT((fsm_output(6)) AND (NOT mux_925_nl));
  or_875_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0110"));
  mux_926_nl <= MUX_s_1_2_2(nand_46_nl, or_875_nl, fsm_output(7));
  nor_529_nl <= NOT((fsm_output(8)) OR mux_926_nl);
  and_438_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (NOT (VEC_LOOP_j_sva_9_0(0))) AND (NOT (fsm_output(5))) AND (fsm_output(1));
  or_871_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_921_nl <= MUX_s_1_2_2(or_871_nl, or_tmp_817, fsm_output(0));
  nor_531_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_921_nl);
  mux_922_nl <= MUX_s_1_2_2(and_438_nl, nor_531_nl, fsm_output(8));
  mux_927_nl <= MUX_s_1_2_2(nor_529_nl, mux_922_nl, fsm_output(9));
  or_868_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_866_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_916_nl <= MUX_s_1_2_2(or_866_nl, or_tmp_817, fsm_output(0));
  or_864_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_915_nl <= MUX_s_1_2_2(or_tmp_816, or_864_nl, fsm_output(0));
  mux_917_nl <= MUX_s_1_2_2(mux_916_nl, mux_915_nl, fsm_output(4));
  or_862_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_914_nl <= MUX_s_1_2_2(or_862_nl, or_tmp_811, fsm_output(0));
  or_863_nl <= (fsm_output(4)) OR mux_914_nl;
  mux_918_nl <= MUX_s_1_2_2(mux_917_nl, or_863_nl, fsm_output(6));
  mux_919_nl <= MUX_s_1_2_2(or_868_nl, mux_918_nl, fsm_output(7));
  and_326_nl <= (fsm_output(8)) AND (NOT mux_919_nl);
  nor_532_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")));
  mux_920_nl <= MUX_s_1_2_2(and_326_nl, nor_532_nl, fsm_output(9));
  mux_928_nl <= MUX_s_1_2_2(mux_927_nl, mux_920_nl, fsm_output(3));
  or_859_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_857_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_909_nl <= MUX_s_1_2_2(or_857_nl, or_tmp_817, fsm_output(0));
  or_855_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_908_nl <= MUX_s_1_2_2(or_tmp_816, or_855_nl, fsm_output(0));
  mux_910_nl <= MUX_s_1_2_2(mux_909_nl, mux_908_nl, fsm_output(4));
  mux_911_nl <= MUX_s_1_2_2(or_859_nl, mux_910_nl, fsm_output(6));
  or_853_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_906_nl <= MUX_s_1_2_2(or_853_nl, or_tmp_811, fsm_output(0));
  or_854_nl <= (fsm_output(4)) OR mux_906_nl;
  mux_907_nl <= MUX_s_1_2_2(or_854_nl, or_tmp_810, fsm_output(6));
  mux_912_nl <= MUX_s_1_2_2(mux_911_nl, mux_907_nl, fsm_output(7));
  nor_533_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_912_nl);
  or_850_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5))
      OR (NOT (fsm_output(1)));
  or_848_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_902_nl <= MUX_s_1_2_2(or_848_nl, or_tmp_817, fsm_output(0));
  or_844_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_901_nl <= MUX_s_1_2_2(or_tmp_816, or_844_nl, fsm_output(0));
  mux_903_nl <= MUX_s_1_2_2(mux_902_nl, mux_901_nl, fsm_output(4));
  mux_904_nl <= MUX_s_1_2_2(or_850_nl, mux_903_nl, fsm_output(6));
  nand_44_nl <= NOT((fsm_output(7)) AND (NOT mux_904_nl));
  or_841_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_899_nl <= MUX_s_1_2_2(or_841_nl, or_tmp_811, fsm_output(0));
  or_842_nl <= (fsm_output(4)) OR mux_899_nl;
  mux_900_nl <= MUX_s_1_2_2(or_842_nl, or_tmp_810, fsm_output(6));
  or_843_nl <= (fsm_output(7)) OR mux_900_nl;
  mux_905_nl <= MUX_s_1_2_2(nand_44_nl, or_843_nl, fsm_output(8));
  nor_534_nl <= NOT((fsm_output(9)) OR mux_905_nl);
  mux_913_nl <= MUX_s_1_2_2(nor_533_nl, nor_534_nl, fsm_output(3));
  vec_rsc_0_6_i_we_d_pff <= MUX_s_1_2_2(mux_928_nl, mux_913_nl, fsm_output(2));
  nor_518_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_926_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR not_tmp_133;
  or_927_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_930_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_929_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_955_nl <= MUX_s_1_2_2(or_929_nl, or_927_cse, fsm_output(0));
  mux_956_nl <= MUX_s_1_2_2(or_930_nl, mux_955_nl, fsm_output(6));
  or_924_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR
      (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_953_nl <= MUX_s_1_2_2(or_926_cse, or_924_nl, fsm_output(0));
  or_923_nl <= (VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_921_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_952_nl <= MUX_s_1_2_2(or_923_nl, or_921_nl, fsm_output(0));
  mux_954_nl <= MUX_s_1_2_2(mux_953_nl, mux_952_nl, fsm_output(6));
  mux_957_nl <= MUX_s_1_2_2(mux_956_nl, mux_954_nl, fsm_output(1));
  nor_509_nl <= NOT((fsm_output(3)) OR mux_957_nl);
  or_919_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_917_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR
      (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_949_nl <= MUX_s_1_2_2(or_919_nl, or_917_nl, fsm_output(0));
  or_916_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_950_nl <= MUX_s_1_2_2(mux_949_nl, or_916_nl, fsm_output(6));
  nor_510_nl <= NOT((fsm_output(1)) OR mux_950_nl);
  nor_511_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0110"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_951_nl <= MUX_s_1_2_2(nor_510_nl, nor_511_nl, fsm_output(3));
  mux_958_nl <= MUX_s_1_2_2(nor_509_nl, mux_951_nl, fsm_output(2));
  nor_512_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0110")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_513_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_514_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_515_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR not_tmp_133);
  mux_945_nl <= MUX_s_1_2_2(nor_514_nl, nor_515_nl, fsm_output(0));
  mux_946_nl <= MUX_s_1_2_2(nor_513_nl, mux_945_nl, fsm_output(6));
  and_324_nl <= (fsm_output(1)) AND mux_946_nl;
  mux_947_nl <= MUX_s_1_2_2(nor_512_nl, and_324_nl, fsm_output(3));
  nor_516_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_517_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_942_nl <= MUX_s_1_2_2(nor_516_nl, nor_517_nl, fsm_output(0));
  nor_519_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_941_nl <= MUX_s_1_2_2(nor_518_cse, nor_519_nl, fsm_output(0));
  mux_943_nl <= MUX_s_1_2_2(mux_942_nl, mux_941_nl, fsm_output(6));
  nor_520_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_521_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_939_nl <= MUX_s_1_2_2(nor_520_nl, nor_521_nl, fsm_output(0));
  nor_522_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_940_nl <= MUX_s_1_2_2(mux_939_nl, nor_522_nl, fsm_output(6));
  mux_944_nl <= MUX_s_1_2_2(mux_943_nl, mux_940_nl, fsm_output(1));
  and_325_nl <= (fsm_output(3)) AND mux_944_nl;
  mux_948_nl <= MUX_s_1_2_2(mux_947_nl, and_325_nl, fsm_output(2));
  mux_959_nl <= MUX_s_1_2_2(mux_958_nl, mux_948_nl, fsm_output(8));
  nor_525_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_935_nl <= MUX_s_1_2_2(nor_518_cse, nor_525_nl, fsm_output(0));
  nor_526_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_527_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_934_nl <= MUX_s_1_2_2(nor_526_nl, nor_527_nl, fsm_output(0));
  mux_936_nl <= MUX_s_1_2_2(mux_935_nl, mux_934_nl, fsm_output(6));
  nor_528_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_937_nl <= MUX_s_1_2_2(mux_936_nl, nor_528_nl, fsm_output(1));
  nand_47_nl <= NOT((fsm_output(3)) AND mux_937_nl);
  or_886_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_884_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_931_nl <= MUX_s_1_2_2(or_884_nl, or_926_cse, fsm_output(0));
  or_880_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_930_nl <= MUX_s_1_2_2(or_927_cse, or_880_nl, fsm_output(0));
  mux_932_nl <= MUX_s_1_2_2(mux_931_nl, mux_930_nl, fsm_output(6));
  mux_933_nl <= MUX_s_1_2_2(or_886_nl, mux_932_nl, fsm_output(1));
  or_887_nl <= (fsm_output(3)) OR mux_933_nl;
  mux_938_nl <= MUX_s_1_2_2(nand_47_nl, or_887_nl, fsm_output(2));
  nor_523_nl <= NOT((fsm_output(8)) OR mux_938_nl);
  vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_959_nl, nor_523_nl,
      fsm_output(9));
  or_970_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_986_nl <= MUX_s_1_2_2(or_tmp_910, or_970_nl, fsm_output(0));
  or_969_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_985_nl <= MUX_s_1_2_2(or_969_nl, or_tmp_904, fsm_output(0));
  mux_987_nl <= MUX_s_1_2_2(mux_986_nl, mux_985_nl, fsm_output(4));
  nand_52_nl <= NOT((fsm_output(6)) AND (NOT mux_987_nl));
  or_968_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0111"));
  mux_988_nl <= MUX_s_1_2_2(nand_52_nl, or_968_nl, fsm_output(7));
  nor_503_nl <= NOT((fsm_output(8)) OR mux_988_nl);
  and_437_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT (fsm_output(5))) AND (fsm_output(1));
  or_964_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_983_nl <= MUX_s_1_2_2(or_964_nl, or_tmp_910, fsm_output(0));
  nor_505_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_983_nl);
  mux_984_nl <= MUX_s_1_2_2(and_437_nl, nor_505_nl, fsm_output(8));
  mux_989_nl <= MUX_s_1_2_2(nor_503_nl, mux_984_nl, fsm_output(9));
  nand_376_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0))
      AND (NOT (fsm_output(5))) AND (fsm_output(1)));
  or_959_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_978_nl <= MUX_s_1_2_2(or_959_nl, or_tmp_910, fsm_output(0));
  or_957_nl <= (COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_977_nl <= MUX_s_1_2_2(or_tmp_909, or_957_nl, fsm_output(0));
  mux_979_nl <= MUX_s_1_2_2(mux_978_nl, mux_977_nl, fsm_output(4));
  or_955_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_976_nl <= MUX_s_1_2_2(or_955_nl, or_tmp_904, fsm_output(0));
  or_956_nl <= (fsm_output(4)) OR mux_976_nl;
  mux_980_nl <= MUX_s_1_2_2(mux_979_nl, or_956_nl, fsm_output(6));
  mux_981_nl <= MUX_s_1_2_2(nand_376_nl, mux_980_nl, fsm_output(7));
  and_323_nl <= (fsm_output(8)) AND (NOT mux_981_nl);
  nor_506_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")));
  mux_982_nl <= MUX_s_1_2_2(and_323_nl, nor_506_nl, fsm_output(9));
  mux_990_nl <= MUX_s_1_2_2(mux_989_nl, mux_982_nl, fsm_output(3));
  nand_371_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (fsm_output(4)) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT
      (fsm_output(5))) AND (fsm_output(1)));
  or_950_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_971_nl <= MUX_s_1_2_2(or_950_nl, or_tmp_910, fsm_output(0));
  or_948_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_970_nl <= MUX_s_1_2_2(or_tmp_909, or_948_nl, fsm_output(0));
  mux_972_nl <= MUX_s_1_2_2(mux_971_nl, mux_970_nl, fsm_output(4));
  mux_973_nl <= MUX_s_1_2_2(nand_371_nl, mux_972_nl, fsm_output(6));
  or_946_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_968_nl <= MUX_s_1_2_2(or_946_nl, or_tmp_904, fsm_output(0));
  or_947_nl <= (fsm_output(4)) OR mux_968_nl;
  mux_969_nl <= MUX_s_1_2_2(or_947_nl, or_tmp_903, fsm_output(6));
  mux_974_nl <= MUX_s_1_2_2(mux_973_nl, mux_969_nl, fsm_output(7));
  nor_507_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_974_nl);
  nand_360_nl <= NOT((fsm_output(4)) AND (fsm_output(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("011")) AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT (fsm_output(5)))
      AND (fsm_output(1)));
  or_941_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_964_nl <= MUX_s_1_2_2(or_941_nl, or_tmp_910, fsm_output(0));
  or_937_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_963_nl <= MUX_s_1_2_2(or_tmp_909, or_937_nl, fsm_output(0));
  mux_965_nl <= MUX_s_1_2_2(mux_964_nl, mux_963_nl, fsm_output(4));
  mux_966_nl <= MUX_s_1_2_2(nand_360_nl, mux_965_nl, fsm_output(6));
  nand_50_nl <= NOT((fsm_output(7)) AND (NOT mux_966_nl));
  or_934_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_961_nl <= MUX_s_1_2_2(or_934_nl, or_tmp_904, fsm_output(0));
  or_935_nl <= (fsm_output(4)) OR mux_961_nl;
  mux_962_nl <= MUX_s_1_2_2(or_935_nl, or_tmp_903, fsm_output(6));
  or_936_nl <= (fsm_output(7)) OR mux_962_nl;
  mux_967_nl <= MUX_s_1_2_2(nand_50_nl, or_936_nl, fsm_output(8));
  nor_508_nl <= NOT((fsm_output(9)) OR mux_967_nl);
  mux_975_nl <= MUX_s_1_2_2(nor_507_nl, nor_508_nl, fsm_output(3));
  vec_rsc_0_7_i_we_d_pff <= MUX_s_1_2_2(mux_990_nl, mux_975_nl, fsm_output(2));
  nor_492_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nand_280_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111")));
  nand_275_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  nand_274_nl <= NOT((fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND
      CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_1022_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_1017_nl <= MUX_s_1_2_2(or_1022_nl, nand_275_cse, fsm_output(0));
  mux_1018_nl <= MUX_s_1_2_2(nand_274_nl, mux_1017_nl, fsm_output(6));
  or_1019_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("011")) OR
      nand_308_cse;
  or_1017_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_1015_nl <= MUX_s_1_2_2(or_1019_nl, or_1017_nl, fsm_output(0));
  nand_370_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("011")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4)));
  or_1014_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1014_nl <= MUX_s_1_2_2(nand_370_nl, or_1014_nl, fsm_output(0));
  mux_1016_nl <= MUX_s_1_2_2(mux_1015_nl, mux_1014_nl, fsm_output(6));
  mux_1019_nl <= MUX_s_1_2_2(mux_1018_nl, mux_1016_nl, fsm_output(1));
  nor_484_nl <= NOT((fsm_output(3)) OR mux_1019_nl);
  or_1012_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1010_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_1011_nl <= MUX_s_1_2_2(or_1012_nl, or_1010_nl, fsm_output(0));
  or_1009_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1012_nl <= MUX_s_1_2_2(mux_1011_nl, or_1009_nl, fsm_output(6));
  nor_485_nl <= NOT((fsm_output(1)) OR mux_1012_nl);
  nor_486_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_1013_nl <= MUX_s_1_2_2(nor_485_nl, nor_486_nl, fsm_output(3));
  mux_1020_nl <= MUX_s_1_2_2(nor_484_nl, mux_1013_nl, fsm_output(2));
  nor_487_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0111")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_488_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) OR not_tmp_133);
  and_321_nl <= (VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("011")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4)));
  nor_489_nl <= NOT(nand_280_cse OR not_tmp_133);
  mux_1007_nl <= MUX_s_1_2_2(and_321_nl, nor_489_nl, fsm_output(0));
  mux_1008_nl <= MUX_s_1_2_2(nor_488_nl, mux_1007_nl, fsm_output(6));
  and_320_nl <= (fsm_output(1)) AND mux_1008_nl;
  mux_1009_nl <= MUX_s_1_2_2(nor_487_nl, and_320_nl, fsm_output(3));
  nor_490_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("111")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_491_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_1004_nl <= MUX_s_1_2_2(nor_490_nl, nor_491_nl, fsm_output(0));
  nor_493_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1003_nl <= MUX_s_1_2_2(nor_492_cse, nor_493_nl, fsm_output(0));
  mux_1005_nl <= MUX_s_1_2_2(mux_1004_nl, mux_1003_nl, fsm_output(6));
  nor_494_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  and_432_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111")) AND
      (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4));
  mux_1001_nl <= MUX_s_1_2_2(nor_494_nl, and_432_nl, fsm_output(0));
  nor_496_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1002_nl <= MUX_s_1_2_2(mux_1001_nl, nor_496_nl, fsm_output(6));
  mux_1006_nl <= MUX_s_1_2_2(mux_1005_nl, mux_1002_nl, fsm_output(1));
  and_322_nl <= (fsm_output(3)) AND mux_1006_nl;
  mux_1010_nl <= MUX_s_1_2_2(mux_1009_nl, and_322_nl, fsm_output(2));
  mux_1021_nl <= MUX_s_1_2_2(mux_1020_nl, mux_1010_nl, fsm_output(8));
  nor_499_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_997_nl <= MUX_s_1_2_2(nor_492_cse, nor_499_nl, fsm_output(0));
  nor_500_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_501_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_996_nl <= MUX_s_1_2_2(nor_500_nl, nor_501_nl, fsm_output(0));
  mux_998_nl <= MUX_s_1_2_2(mux_997_nl, mux_996_nl, fsm_output(6));
  nor_502_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0111"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_999_nl <= MUX_s_1_2_2(mux_998_nl, nor_502_nl, fsm_output(1));
  nand_53_nl <= NOT((fsm_output(3)) AND mux_999_nl);
  or_979_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      AND (NOT (fsm_output(5))))) OR not_tmp_134;
  nand_282_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))
      AND (VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5))
      AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_976_nl <= nand_280_cse OR not_tmp_133;
  mux_993_nl <= MUX_s_1_2_2(nand_282_nl, or_976_nl, fsm_output(0));
  nand_354_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5)) AND (NOT (fsm_output(7)))
      AND (fsm_output(4)));
  mux_992_nl <= MUX_s_1_2_2(nand_275_cse, nand_354_nl, fsm_output(0));
  mux_994_nl <= MUX_s_1_2_2(mux_993_nl, mux_992_nl, fsm_output(6));
  mux_995_nl <= MUX_s_1_2_2(or_979_nl, mux_994_nl, fsm_output(1));
  or_980_nl <= (fsm_output(3)) OR mux_995_nl;
  mux_1000_nl <= MUX_s_1_2_2(nand_53_nl, or_980_nl, fsm_output(2));
  nor_497_nl <= NOT((fsm_output(8)) OR mux_1000_nl);
  vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1021_nl, nor_497_nl,
      fsm_output(9));
  or_1069_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_1048_nl <= MUX_s_1_2_2(or_tmp_1007, or_1069_nl, fsm_output(0));
  or_1068_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1047_nl <= MUX_s_1_2_2(or_1068_nl, or_tmp_999, fsm_output(0));
  mux_1049_nl <= MUX_s_1_2_2(mux_1048_nl, mux_1047_nl, fsm_output(4));
  nand_58_nl <= NOT((fsm_output(6)) AND (NOT mux_1049_nl));
  or_1067_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1000"));
  mux_1050_nl <= MUX_s_1_2_2(nand_58_nl, or_1067_nl, fsm_output(7));
  nor_478_nl <= NOT((fsm_output(8)) OR mux_1050_nl);
  nor_479_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(7))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT
      (fsm_output(1))));
  or_1062_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1045_nl <= MUX_s_1_2_2(or_1062_nl, or_tmp_1007, fsm_output(0));
  nor_480_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_1045_nl);
  mux_1046_nl <= MUX_s_1_2_2(nor_479_nl, nor_480_nl, fsm_output(8));
  mux_1051_nl <= MUX_s_1_2_2(nor_478_nl, mux_1046_nl, fsm_output(9));
  or_1059_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_1057_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1040_nl <= MUX_s_1_2_2(or_1057_nl, or_tmp_1007, fsm_output(0));
  or_1055_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1039_nl <= MUX_s_1_2_2(or_tmp_1005, or_1055_nl, fsm_output(0));
  mux_1041_nl <= MUX_s_1_2_2(mux_1040_nl, mux_1039_nl, fsm_output(4));
  or_1053_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1038_nl <= MUX_s_1_2_2(or_1053_nl, or_tmp_999, fsm_output(0));
  or_1054_nl <= (fsm_output(4)) OR mux_1038_nl;
  mux_1042_nl <= MUX_s_1_2_2(mux_1041_nl, or_1054_nl, fsm_output(6));
  mux_1043_nl <= MUX_s_1_2_2(or_1059_nl, mux_1042_nl, fsm_output(7));
  and_319_nl <= (fsm_output(8)) AND (NOT mux_1043_nl);
  nor_481_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")));
  mux_1044_nl <= MUX_s_1_2_2(and_319_nl, nor_481_nl, fsm_output(9));
  mux_1052_nl <= MUX_s_1_2_2(mux_1051_nl, mux_1044_nl, fsm_output(3));
  or_1049_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_1047_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1033_nl <= MUX_s_1_2_2(or_1047_nl, or_tmp_1007, fsm_output(0));
  or_1045_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1032_nl <= MUX_s_1_2_2(or_tmp_1005, or_1045_nl, fsm_output(0));
  mux_1034_nl <= MUX_s_1_2_2(mux_1033_nl, mux_1032_nl, fsm_output(4));
  mux_1035_nl <= MUX_s_1_2_2(or_1049_nl, mux_1034_nl, fsm_output(6));
  or_1043_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1030_nl <= MUX_s_1_2_2(or_1043_nl, or_tmp_999, fsm_output(0));
  or_1044_nl <= (fsm_output(4)) OR mux_1030_nl;
  mux_1031_nl <= MUX_s_1_2_2(or_1044_nl, or_tmp_997, fsm_output(6));
  mux_1036_nl <= MUX_s_1_2_2(mux_1035_nl, mux_1031_nl, fsm_output(7));
  nor_482_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1036_nl);
  or_1040_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5))
      OR (NOT (fsm_output(1)));
  or_1038_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1026_nl <= MUX_s_1_2_2(or_1038_nl, or_tmp_1007, fsm_output(0));
  or_1032_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1025_nl <= MUX_s_1_2_2(or_tmp_1005, or_1032_nl, fsm_output(0));
  mux_1027_nl <= MUX_s_1_2_2(mux_1026_nl, mux_1025_nl, fsm_output(4));
  mux_1028_nl <= MUX_s_1_2_2(or_1040_nl, mux_1027_nl, fsm_output(6));
  nand_56_nl <= NOT((fsm_output(7)) AND (NOT mux_1028_nl));
  or_1029_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1023_nl <= MUX_s_1_2_2(or_1029_nl, or_tmp_999, fsm_output(0));
  or_1030_nl <= (fsm_output(4)) OR mux_1023_nl;
  mux_1024_nl <= MUX_s_1_2_2(or_1030_nl, or_tmp_997, fsm_output(6));
  or_1031_nl <= (fsm_output(7)) OR mux_1024_nl;
  mux_1029_nl <= MUX_s_1_2_2(nand_56_nl, or_1031_nl, fsm_output(8));
  nor_483_nl <= NOT((fsm_output(9)) OR mux_1029_nl);
  mux_1037_nl <= MUX_s_1_2_2(nor_482_nl, nor_483_nl, fsm_output(3));
  vec_rsc_0_8_i_we_d_pff <= MUX_s_1_2_2(mux_1052_nl, mux_1037_nl, fsm_output(2));
  nor_467_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_1119_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1122_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1121_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_1079_nl <= MUX_s_1_2_2(or_1121_nl, or_1119_cse, fsm_output(0));
  mux_1080_nl <= MUX_s_1_2_2(or_1122_nl, mux_1079_nl, fsm_output(6));
  or_1118_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR not_tmp_133;
  or_1116_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_1077_nl <= MUX_s_1_2_2(or_1118_nl, or_1116_nl, fsm_output(0));
  or_1115_nl <= (VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1113_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1076_nl <= MUX_s_1_2_2(or_1115_nl, or_1113_nl, fsm_output(0));
  mux_1078_nl <= MUX_s_1_2_2(mux_1077_nl, mux_1076_nl, fsm_output(6));
  mux_1081_nl <= MUX_s_1_2_2(mux_1080_nl, mux_1078_nl, fsm_output(1));
  nor_458_nl <= NOT((fsm_output(3)) OR mux_1081_nl);
  or_1111_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1109_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_1073_nl <= MUX_s_1_2_2(or_1111_nl, or_1109_nl, fsm_output(0));
  or_1108_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1074_nl <= MUX_s_1_2_2(mux_1073_nl, or_1108_nl, fsm_output(6));
  nor_459_nl <= NOT((fsm_output(1)) OR mux_1074_nl);
  nor_460_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0)))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  mux_1075_nl <= MUX_s_1_2_2(nor_459_nl, nor_460_nl, fsm_output(3));
  mux_1082_nl <= MUX_s_1_2_2(nor_458_nl, mux_1075_nl, fsm_output(2));
  nor_461_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1000")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_462_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_463_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_464_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_270_cse_1);
  mux_1069_nl <= MUX_s_1_2_2(nor_463_nl, nor_464_nl, fsm_output(0));
  mux_1070_nl <= MUX_s_1_2_2(nor_462_nl, mux_1069_nl, fsm_output(6));
  and_317_nl <= (fsm_output(1)) AND mux_1070_nl;
  mux_1071_nl <= MUX_s_1_2_2(nor_461_nl, and_317_nl, fsm_output(3));
  nor_465_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_466_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_1066_nl <= MUX_s_1_2_2(nor_465_nl, nor_466_nl, fsm_output(0));
  nor_468_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1065_nl <= MUX_s_1_2_2(nor_467_cse, nor_468_nl, fsm_output(0));
  mux_1067_nl <= MUX_s_1_2_2(mux_1066_nl, mux_1065_nl, fsm_output(6));
  nor_469_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_470_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1063_nl <= MUX_s_1_2_2(nor_469_nl, nor_470_nl, fsm_output(0));
  nor_471_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1064_nl <= MUX_s_1_2_2(mux_1063_nl, nor_471_nl, fsm_output(6));
  mux_1068_nl <= MUX_s_1_2_2(mux_1067_nl, mux_1064_nl, fsm_output(1));
  and_318_nl <= (fsm_output(3)) AND mux_1068_nl;
  mux_1072_nl <= MUX_s_1_2_2(mux_1071_nl, and_318_nl, fsm_output(2));
  mux_1083_nl <= MUX_s_1_2_2(mux_1082_nl, mux_1072_nl, fsm_output(8));
  nor_474_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1059_nl <= MUX_s_1_2_2(nor_467_cse, nor_474_nl, fsm_output(0));
  nor_475_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_476_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1058_nl <= MUX_s_1_2_2(nor_475_nl, nor_476_nl, fsm_output(0));
  mux_1060_nl <= MUX_s_1_2_2(mux_1059_nl, mux_1058_nl, fsm_output(6));
  nor_477_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_1061_nl <= MUX_s_1_2_2(mux_1060_nl, nor_477_nl, fsm_output(1));
  nand_59_nl <= NOT((fsm_output(3)) AND mux_1061_nl);
  or_1078_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_1076_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1075_nl <= CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR
      nand_270_cse_1;
  mux_1055_nl <= MUX_s_1_2_2(or_1076_nl, or_1075_nl, fsm_output(0));
  or_1072_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_1054_nl <= MUX_s_1_2_2(or_1119_cse, or_1072_nl, fsm_output(0));
  mux_1056_nl <= MUX_s_1_2_2(mux_1055_nl, mux_1054_nl, fsm_output(6));
  mux_1057_nl <= MUX_s_1_2_2(or_1078_nl, mux_1056_nl, fsm_output(1));
  or_1079_nl <= (fsm_output(3)) OR mux_1057_nl;
  mux_1062_nl <= MUX_s_1_2_2(nand_59_nl, or_1079_nl, fsm_output(2));
  nor_472_nl <= NOT((fsm_output(8)) OR mux_1062_nl);
  vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1083_nl, nor_472_nl,
      fsm_output(9));
  or_1169_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(1)) OR (fsm_output(5));
  mux_1110_nl <= MUX_s_1_2_2(or_tmp_1106, or_1169_nl, fsm_output(0));
  or_1168_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1109_nl <= MUX_s_1_2_2(or_1168_nl, or_tmp_1097, fsm_output(0));
  mux_1111_nl <= MUX_s_1_2_2(mux_1110_nl, mux_1109_nl, fsm_output(4));
  nor_450_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(6))) OR mux_1111_nl);
  or_1166_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_9_0(0)))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  or_1165_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1106_nl <= MUX_s_1_2_2(or_1165_nl, or_tmp_1106, fsm_output(0));
  or_1164_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1105_nl <= MUX_s_1_2_2(or_tmp_1104, or_1164_nl, fsm_output(0));
  mux_1107_nl <= MUX_s_1_2_2(mux_1106_nl, mux_1105_nl, fsm_output(4));
  mux_1108_nl <= MUX_s_1_2_2(or_1166_nl, mux_1107_nl, fsm_output(6));
  and_316_nl <= (fsm_output(9)) AND (NOT mux_1108_nl);
  mux_1112_nl <= MUX_s_1_2_2(nor_450_nl, and_316_nl, fsm_output(2));
  or_1161_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1104_nl <= MUX_s_1_2_2(or_1161_nl, or_tmp_1106, fsm_output(0));
  nor_451_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR
      (fsm_output(4)) OR mux_1104_nl);
  mux_1113_nl <= MUX_s_1_2_2(mux_1112_nl, nor_451_nl, fsm_output(8));
  or_1158_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(1))
      OR (NOT (fsm_output(5))) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"));
  or_1156_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1102_nl <= MUX_s_1_2_2(or_1158_nl, or_1156_nl, fsm_output(9));
  or_1154_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1100_nl <= MUX_s_1_2_2(or_1154_nl, or_tmp_1097, fsm_output(0));
  or_1155_nl <= (fsm_output(4)) OR mux_1100_nl;
  mux_1101_nl <= MUX_s_1_2_2(or_1155_nl, or_tmp_1116, fsm_output(6));
  nand_62_nl <= NOT((fsm_output(9)) AND (NOT mux_1101_nl));
  mux_1103_nl <= MUX_s_1_2_2(mux_1102_nl, nand_62_nl, fsm_output(2));
  nor_452_nl <= NOT((fsm_output(8)) OR mux_1103_nl);
  mux_1114_nl <= MUX_s_1_2_2(mux_1113_nl, nor_452_nl, fsm_output(7));
  nor_453_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR
      (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))
      OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")));
  nor_454_nl <= NOT((fsm_output(9)) OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("100")) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(0))) OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT (fsm_output(1)))
      OR (fsm_output(5)));
  or_1147_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1095_nl <= MUX_s_1_2_2(or_1147_nl, or_tmp_1097, fsm_output(0));
  or_1148_nl <= (fsm_output(4)) OR mux_1095_nl;
  mux_1096_nl <= MUX_s_1_2_2(or_1148_nl, or_tmp_1116, fsm_output(6));
  nor_455_nl <= NOT((fsm_output(9)) OR mux_1096_nl);
  mux_1097_nl <= MUX_s_1_2_2(nor_454_nl, nor_455_nl, fsm_output(2));
  mux_1098_nl <= MUX_s_1_2_2(nor_453_nl, mux_1097_nl, fsm_output(8));
  or_1142_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT
      (fsm_output(1))) OR (fsm_output(5));
  or_1141_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1091_nl <= MUX_s_1_2_2(or_1141_nl, or_tmp_1106, fsm_output(0));
  or_1140_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1090_nl <= MUX_s_1_2_2(or_tmp_1104, or_1140_nl, fsm_output(0));
  mux_1092_nl <= MUX_s_1_2_2(mux_1091_nl, mux_1090_nl, fsm_output(4));
  mux_1093_nl <= MUX_s_1_2_2(or_1142_nl, mux_1092_nl, fsm_output(6));
  nor_456_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(9)) OR mux_1093_nl);
  or_1136_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1087_nl <= MUX_s_1_2_2(or_1136_nl, or_tmp_1106, fsm_output(0));
  or_1131_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1086_nl <= MUX_s_1_2_2(or_tmp_1104, or_1131_nl, fsm_output(0));
  mux_1088_nl <= MUX_s_1_2_2(mux_1087_nl, mux_1086_nl, fsm_output(4));
  or_1128_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1085_nl <= MUX_s_1_2_2(or_1128_nl, or_tmp_1097, fsm_output(0));
  or_1129_nl <= (fsm_output(4)) OR mux_1085_nl;
  mux_1089_nl <= MUX_s_1_2_2(mux_1088_nl, or_1129_nl, fsm_output(6));
  nor_457_nl <= NOT((fsm_output(2)) OR (fsm_output(9)) OR mux_1089_nl);
  mux_1094_nl <= MUX_s_1_2_2(nor_456_nl, nor_457_nl, fsm_output(8));
  mux_1099_nl <= MUX_s_1_2_2(mux_1098_nl, mux_1094_nl, fsm_output(7));
  vec_rsc_0_9_i_we_d_pff <= MUX_s_1_2_2(mux_1114_nl, mux_1099_nl, fsm_output(3));
  nor_439_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_1218_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1221_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1220_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_1141_nl <= MUX_s_1_2_2(or_1220_nl, or_1218_cse, fsm_output(0));
  mux_1142_nl <= MUX_s_1_2_2(or_1221_nl, mux_1141_nl, fsm_output(6));
  or_1217_nl <= CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR
      nand_264_cse;
  or_1215_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_1139_nl <= MUX_s_1_2_2(or_1217_nl, or_1215_nl, fsm_output(0));
  or_1214_nl <= (NOT (VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1212_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1138_nl <= MUX_s_1_2_2(or_1214_nl, or_1212_nl, fsm_output(0));
  mux_1140_nl <= MUX_s_1_2_2(mux_1139_nl, mux_1138_nl, fsm_output(6));
  mux_1143_nl <= MUX_s_1_2_2(mux_1142_nl, mux_1140_nl, fsm_output(1));
  nor_430_nl <= NOT((fsm_output(3)) OR mux_1143_nl);
  or_1210_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1208_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_1135_nl <= MUX_s_1_2_2(or_1210_nl, or_1208_nl, fsm_output(0));
  or_1207_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1136_nl <= MUX_s_1_2_2(mux_1135_nl, or_1207_nl, fsm_output(6));
  nor_431_nl <= NOT((fsm_output(1)) OR mux_1136_nl);
  nor_432_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1001"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_1137_nl <= MUX_s_1_2_2(nor_431_nl, nor_432_nl, fsm_output(3));
  mux_1144_nl <= MUX_s_1_2_2(nor_430_nl, mux_1137_nl, fsm_output(2));
  nor_433_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1001")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_434_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_435_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_436_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_270_cse_1);
  mux_1131_nl <= MUX_s_1_2_2(nor_435_nl, nor_436_nl, fsm_output(0));
  mux_1132_nl <= MUX_s_1_2_2(nor_434_nl, mux_1131_nl, fsm_output(6));
  and_314_nl <= (fsm_output(1)) AND mux_1132_nl;
  mux_1133_nl <= MUX_s_1_2_2(nor_433_nl, and_314_nl, fsm_output(3));
  nor_437_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_438_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_1128_nl <= MUX_s_1_2_2(nor_437_nl, nor_438_nl, fsm_output(0));
  nor_440_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1127_nl <= MUX_s_1_2_2(nor_439_cse, nor_440_nl, fsm_output(0));
  mux_1129_nl <= MUX_s_1_2_2(mux_1128_nl, mux_1127_nl, fsm_output(6));
  nor_441_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_442_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1125_nl <= MUX_s_1_2_2(nor_441_nl, nor_442_nl, fsm_output(0));
  nor_443_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1126_nl <= MUX_s_1_2_2(mux_1125_nl, nor_443_nl, fsm_output(6));
  mux_1130_nl <= MUX_s_1_2_2(mux_1129_nl, mux_1126_nl, fsm_output(1));
  and_315_nl <= (fsm_output(3)) AND mux_1130_nl;
  mux_1134_nl <= MUX_s_1_2_2(mux_1133_nl, and_315_nl, fsm_output(2));
  mux_1145_nl <= MUX_s_1_2_2(mux_1144_nl, mux_1134_nl, fsm_output(8));
  nor_446_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1121_nl <= MUX_s_1_2_2(nor_439_cse, nor_446_nl, fsm_output(0));
  nor_447_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_448_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1120_nl <= MUX_s_1_2_2(nor_447_nl, nor_448_nl, fsm_output(0));
  mux_1122_nl <= MUX_s_1_2_2(mux_1121_nl, mux_1120_nl, fsm_output(6));
  nor_449_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_1123_nl <= MUX_s_1_2_2(mux_1122_nl, nor_449_nl, fsm_output(1));
  nand_65_nl <= NOT((fsm_output(3)) AND mux_1123_nl);
  or_1177_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_1175_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1174_nl <= CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR
      nand_270_cse_1;
  mux_1117_nl <= MUX_s_1_2_2(or_1175_nl, or_1174_nl, fsm_output(0));
  or_1171_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_1116_nl <= MUX_s_1_2_2(or_1218_cse, or_1171_nl, fsm_output(0));
  mux_1118_nl <= MUX_s_1_2_2(mux_1117_nl, mux_1116_nl, fsm_output(6));
  mux_1119_nl <= MUX_s_1_2_2(or_1177_nl, mux_1118_nl, fsm_output(1));
  or_1178_nl <= (fsm_output(3)) OR mux_1119_nl;
  mux_1124_nl <= MUX_s_1_2_2(nand_65_nl, or_1178_nl, fsm_output(2));
  nor_444_nl <= NOT((fsm_output(8)) OR mux_1124_nl);
  vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1145_nl, nor_444_nl,
      fsm_output(9));
  or_1267_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_1172_nl <= MUX_s_1_2_2(or_tmp_1205, or_1267_nl, fsm_output(0));
  or_1266_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1171_nl <= MUX_s_1_2_2(or_1266_nl, or_tmp_1197, fsm_output(0));
  mux_1173_nl <= MUX_s_1_2_2(mux_1172_nl, mux_1171_nl, fsm_output(4));
  nand_70_nl <= NOT((fsm_output(6)) AND (NOT mux_1173_nl));
  or_1265_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1010"));
  mux_1174_nl <= MUX_s_1_2_2(nand_70_nl, or_1265_nl, fsm_output(7));
  nor_424_nl <= NOT((fsm_output(8)) OR mux_1174_nl);
  and_442_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (NOT (VEC_LOOP_j_sva_9_0(0))) AND (NOT (fsm_output(5))) AND (fsm_output(1));
  or_1260_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1169_nl <= MUX_s_1_2_2(or_1260_nl, or_tmp_1205, fsm_output(0));
  nor_426_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_1169_nl);
  mux_1170_nl <= MUX_s_1_2_2(and_442_nl, nor_426_nl, fsm_output(8));
  mux_1175_nl <= MUX_s_1_2_2(nor_424_nl, mux_1170_nl, fsm_output(9));
  or_1257_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_1255_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1164_nl <= MUX_s_1_2_2(or_1255_nl, or_tmp_1205, fsm_output(0));
  or_1253_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1163_nl <= MUX_s_1_2_2(or_tmp_1203, or_1253_nl, fsm_output(0));
  mux_1165_nl <= MUX_s_1_2_2(mux_1164_nl, mux_1163_nl, fsm_output(4));
  or_1251_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1162_nl <= MUX_s_1_2_2(or_1251_nl, or_tmp_1197, fsm_output(0));
  or_1252_nl <= (fsm_output(4)) OR mux_1162_nl;
  mux_1166_nl <= MUX_s_1_2_2(mux_1165_nl, or_1252_nl, fsm_output(6));
  mux_1167_nl <= MUX_s_1_2_2(or_1257_nl, mux_1166_nl, fsm_output(7));
  and_313_nl <= (fsm_output(8)) AND (NOT mux_1167_nl);
  nor_427_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")));
  mux_1168_nl <= MUX_s_1_2_2(and_313_nl, nor_427_nl, fsm_output(9));
  mux_1176_nl <= MUX_s_1_2_2(mux_1175_nl, mux_1168_nl, fsm_output(3));
  or_1247_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_1245_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1157_nl <= MUX_s_1_2_2(or_1245_nl, or_tmp_1205, fsm_output(0));
  or_1243_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1156_nl <= MUX_s_1_2_2(or_tmp_1203, or_1243_nl, fsm_output(0));
  mux_1158_nl <= MUX_s_1_2_2(mux_1157_nl, mux_1156_nl, fsm_output(4));
  mux_1159_nl <= MUX_s_1_2_2(or_1247_nl, mux_1158_nl, fsm_output(6));
  or_1241_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1154_nl <= MUX_s_1_2_2(or_1241_nl, or_tmp_1197, fsm_output(0));
  or_1242_nl <= (fsm_output(4)) OR mux_1154_nl;
  mux_1155_nl <= MUX_s_1_2_2(or_1242_nl, or_tmp_1195, fsm_output(6));
  mux_1160_nl <= MUX_s_1_2_2(mux_1159_nl, mux_1155_nl, fsm_output(7));
  nor_428_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1160_nl);
  or_1238_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5))
      OR (NOT (fsm_output(1)));
  or_1236_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1150_nl <= MUX_s_1_2_2(or_1236_nl, or_tmp_1205, fsm_output(0));
  or_1230_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1149_nl <= MUX_s_1_2_2(or_tmp_1203, or_1230_nl, fsm_output(0));
  mux_1151_nl <= MUX_s_1_2_2(mux_1150_nl, mux_1149_nl, fsm_output(4));
  mux_1152_nl <= MUX_s_1_2_2(or_1238_nl, mux_1151_nl, fsm_output(6));
  nand_68_nl <= NOT((fsm_output(7)) AND (NOT mux_1152_nl));
  or_1227_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1147_nl <= MUX_s_1_2_2(or_1227_nl, or_tmp_1197, fsm_output(0));
  or_1228_nl <= (fsm_output(4)) OR mux_1147_nl;
  mux_1148_nl <= MUX_s_1_2_2(or_1228_nl, or_tmp_1195, fsm_output(6));
  or_1229_nl <= (fsm_output(7)) OR mux_1148_nl;
  mux_1153_nl <= MUX_s_1_2_2(nand_68_nl, or_1229_nl, fsm_output(8));
  nor_429_nl <= NOT((fsm_output(9)) OR mux_1153_nl);
  mux_1161_nl <= MUX_s_1_2_2(nor_428_nl, nor_429_nl, fsm_output(3));
  vec_rsc_0_10_i_we_d_pff <= MUX_s_1_2_2(mux_1176_nl, mux_1161_nl, fsm_output(2));
  nor_413_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_1317_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1320_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1319_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_1203_nl <= MUX_s_1_2_2(or_1319_nl, or_1317_cse, fsm_output(0));
  mux_1204_nl <= MUX_s_1_2_2(or_1320_nl, mux_1203_nl, fsm_output(6));
  or_1316_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR not_tmp_133;
  or_1314_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_1201_nl <= MUX_s_1_2_2(or_1316_nl, or_1314_nl, fsm_output(0));
  or_1313_nl <= (VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1311_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1200_nl <= MUX_s_1_2_2(or_1313_nl, or_1311_nl, fsm_output(0));
  mux_1202_nl <= MUX_s_1_2_2(mux_1201_nl, mux_1200_nl, fsm_output(6));
  mux_1205_nl <= MUX_s_1_2_2(mux_1204_nl, mux_1202_nl, fsm_output(1));
  nor_404_nl <= NOT((fsm_output(3)) OR mux_1205_nl);
  or_1309_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1307_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_1197_nl <= MUX_s_1_2_2(or_1309_nl, or_1307_nl, fsm_output(0));
  or_1306_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1198_nl <= MUX_s_1_2_2(mux_1197_nl, or_1306_nl, fsm_output(6));
  nor_405_nl <= NOT((fsm_output(1)) OR mux_1198_nl);
  nor_406_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1010"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_1199_nl <= MUX_s_1_2_2(nor_405_nl, nor_406_nl, fsm_output(3));
  mux_1206_nl <= MUX_s_1_2_2(nor_404_nl, mux_1199_nl, fsm_output(2));
  nor_407_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1010")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_408_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_409_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_410_nl <= NOT((z_out_6_10_1(0)) OR (z_out_6_10_1(2)) OR nand_260_cse_1);
  mux_1193_nl <= MUX_s_1_2_2(nor_409_nl, nor_410_nl, fsm_output(0));
  mux_1194_nl <= MUX_s_1_2_2(nor_408_nl, mux_1193_nl, fsm_output(6));
  and_311_nl <= (fsm_output(1)) AND mux_1194_nl;
  mux_1195_nl <= MUX_s_1_2_2(nor_407_nl, and_311_nl, fsm_output(3));
  nor_411_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_412_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_1190_nl <= MUX_s_1_2_2(nor_411_nl, nor_412_nl, fsm_output(0));
  nor_414_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1189_nl <= MUX_s_1_2_2(nor_413_cse, nor_414_nl, fsm_output(0));
  mux_1191_nl <= MUX_s_1_2_2(mux_1190_nl, mux_1189_nl, fsm_output(6));
  nor_415_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_416_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1187_nl <= MUX_s_1_2_2(nor_415_nl, nor_416_nl, fsm_output(0));
  nor_417_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1188_nl <= MUX_s_1_2_2(mux_1187_nl, nor_417_nl, fsm_output(6));
  mux_1192_nl <= MUX_s_1_2_2(mux_1191_nl, mux_1188_nl, fsm_output(1));
  and_312_nl <= (fsm_output(3)) AND mux_1192_nl;
  mux_1196_nl <= MUX_s_1_2_2(mux_1195_nl, and_312_nl, fsm_output(2));
  mux_1207_nl <= MUX_s_1_2_2(mux_1206_nl, mux_1196_nl, fsm_output(8));
  nor_420_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1183_nl <= MUX_s_1_2_2(nor_413_cse, nor_420_nl, fsm_output(0));
  nor_421_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_422_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1182_nl <= MUX_s_1_2_2(nor_421_nl, nor_422_nl, fsm_output(0));
  mux_1184_nl <= MUX_s_1_2_2(mux_1183_nl, mux_1182_nl, fsm_output(6));
  nor_423_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_1185_nl <= MUX_s_1_2_2(mux_1184_nl, nor_423_nl, fsm_output(1));
  nand_71_nl <= NOT((fsm_output(3)) AND mux_1185_nl);
  or_1276_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_1274_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1273_nl <= (z_out_6_10_1(0)) OR (z_out_6_10_1(2)) OR nand_260_cse_1;
  mux_1179_nl <= MUX_s_1_2_2(or_1274_nl, or_1273_nl, fsm_output(0));
  or_1270_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_1178_nl <= MUX_s_1_2_2(or_1317_cse, or_1270_nl, fsm_output(0));
  mux_1180_nl <= MUX_s_1_2_2(mux_1179_nl, mux_1178_nl, fsm_output(6));
  mux_1181_nl <= MUX_s_1_2_2(or_1276_nl, mux_1180_nl, fsm_output(1));
  or_1277_nl <= (fsm_output(3)) OR mux_1181_nl;
  mux_1186_nl <= MUX_s_1_2_2(nand_71_nl, or_1277_nl, fsm_output(2));
  nor_418_nl <= NOT((fsm_output(8)) OR mux_1186_nl);
  vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1207_nl, nor_418_nl,
      fsm_output(9));
  or_1366_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_1234_nl <= MUX_s_1_2_2(or_tmp_1304, or_1366_nl, fsm_output(0));
  or_1365_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1233_nl <= MUX_s_1_2_2(or_1365_nl, or_tmp_1296, fsm_output(0));
  mux_1235_nl <= MUX_s_1_2_2(mux_1234_nl, mux_1233_nl, fsm_output(4));
  nand_76_nl <= NOT((fsm_output(6)) AND (NOT mux_1235_nl));
  or_1364_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("1011"));
  mux_1236_nl <= MUX_s_1_2_2(nand_76_nl, or_1364_nl, fsm_output(7));
  nor_398_nl <= NOT((fsm_output(8)) OR mux_1236_nl);
  and_441_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT (fsm_output(5))) AND (fsm_output(1));
  or_1359_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1231_nl <= MUX_s_1_2_2(or_1359_nl, or_tmp_1304, fsm_output(0));
  nor_400_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_1231_nl);
  mux_1232_nl <= MUX_s_1_2_2(and_441_nl, nor_400_nl, fsm_output(8));
  mux_1237_nl <= MUX_s_1_2_2(nor_398_nl, mux_1232_nl, fsm_output(9));
  nand_378_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0))
      AND (NOT (fsm_output(5))) AND (fsm_output(1)));
  or_1354_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1226_nl <= MUX_s_1_2_2(or_1354_nl, or_tmp_1304, fsm_output(0));
  or_1352_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1225_nl <= MUX_s_1_2_2(or_tmp_1302, or_1352_nl, fsm_output(0));
  mux_1227_nl <= MUX_s_1_2_2(mux_1226_nl, mux_1225_nl, fsm_output(4));
  or_1350_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1224_nl <= MUX_s_1_2_2(or_1350_nl, or_tmp_1296, fsm_output(0));
  or_1351_nl <= (fsm_output(4)) OR mux_1224_nl;
  mux_1228_nl <= MUX_s_1_2_2(mux_1227_nl, or_1351_nl, fsm_output(6));
  mux_1229_nl <= MUX_s_1_2_2(nand_378_nl, mux_1228_nl, fsm_output(7));
  and_310_nl <= (fsm_output(8)) AND (NOT mux_1229_nl);
  nor_401_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")));
  mux_1230_nl <= MUX_s_1_2_2(and_310_nl, nor_401_nl, fsm_output(9));
  mux_1238_nl <= MUX_s_1_2_2(mux_1237_nl, mux_1230_nl, fsm_output(3));
  nand_373_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (fsm_output(4)) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT
      (fsm_output(5))) AND (fsm_output(1)));
  or_1344_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1219_nl <= MUX_s_1_2_2(or_1344_nl, or_tmp_1304, fsm_output(0));
  or_1342_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1218_nl <= MUX_s_1_2_2(or_tmp_1302, or_1342_nl, fsm_output(0));
  mux_1220_nl <= MUX_s_1_2_2(mux_1219_nl, mux_1218_nl, fsm_output(4));
  mux_1221_nl <= MUX_s_1_2_2(nand_373_nl, mux_1220_nl, fsm_output(6));
  or_1340_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1216_nl <= MUX_s_1_2_2(or_1340_nl, or_tmp_1296, fsm_output(0));
  or_1341_nl <= (fsm_output(4)) OR mux_1216_nl;
  mux_1217_nl <= MUX_s_1_2_2(or_1341_nl, or_tmp_1294, fsm_output(6));
  mux_1222_nl <= MUX_s_1_2_2(mux_1221_nl, mux_1217_nl, fsm_output(7));
  nor_402_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1222_nl);
  nand_363_nl <= NOT((fsm_output(4)) AND (fsm_output(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("101")) AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT (fsm_output(5)))
      AND (fsm_output(1)));
  or_1335_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1212_nl <= MUX_s_1_2_2(or_1335_nl, or_tmp_1304, fsm_output(0));
  or_1329_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1211_nl <= MUX_s_1_2_2(or_tmp_1302, or_1329_nl, fsm_output(0));
  mux_1213_nl <= MUX_s_1_2_2(mux_1212_nl, mux_1211_nl, fsm_output(4));
  mux_1214_nl <= MUX_s_1_2_2(nand_363_nl, mux_1213_nl, fsm_output(6));
  nand_74_nl <= NOT((fsm_output(7)) AND (NOT mux_1214_nl));
  or_1326_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1209_nl <= MUX_s_1_2_2(or_1326_nl, or_tmp_1296, fsm_output(0));
  or_1327_nl <= (fsm_output(4)) OR mux_1209_nl;
  mux_1210_nl <= MUX_s_1_2_2(or_1327_nl, or_tmp_1294, fsm_output(6));
  or_1328_nl <= (fsm_output(7)) OR mux_1210_nl;
  mux_1215_nl <= MUX_s_1_2_2(nand_74_nl, or_1328_nl, fsm_output(8));
  nor_403_nl <= NOT((fsm_output(9)) OR mux_1215_nl);
  mux_1223_nl <= MUX_s_1_2_2(nor_402_nl, nor_403_nl, fsm_output(3));
  vec_rsc_0_11_i_we_d_pff <= MUX_s_1_2_2(mux_1238_nl, mux_1223_nl, fsm_output(2));
  nor_387_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nand_241_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  nand_240_nl <= NOT((fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND
      CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_1418_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_1265_nl <= MUX_s_1_2_2(or_1418_nl, nand_241_cse, fsm_output(0));
  mux_1266_nl <= MUX_s_1_2_2(nand_240_nl, mux_1265_nl, fsm_output(6));
  or_1415_nl <= CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      nand_264_cse;
  or_1413_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_1263_nl <= MUX_s_1_2_2(or_1415_nl, or_1413_nl, fsm_output(0));
  nand_369_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("101")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4)));
  or_1410_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1262_nl <= MUX_s_1_2_2(nand_369_nl, or_1410_nl, fsm_output(0));
  mux_1264_nl <= MUX_s_1_2_2(mux_1263_nl, mux_1262_nl, fsm_output(6));
  mux_1267_nl <= MUX_s_1_2_2(mux_1266_nl, mux_1264_nl, fsm_output(1));
  nor_379_nl <= NOT((fsm_output(3)) OR mux_1267_nl);
  or_1408_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1406_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_1259_nl <= MUX_s_1_2_2(or_1408_nl, or_1406_nl, fsm_output(0));
  or_1405_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1260_nl <= MUX_s_1_2_2(mux_1259_nl, or_1405_nl, fsm_output(6));
  nor_380_nl <= NOT((fsm_output(1)) OR mux_1260_nl);
  nor_381_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_1261_nl <= MUX_s_1_2_2(nor_380_nl, nor_381_nl, fsm_output(3));
  mux_1268_nl <= MUX_s_1_2_2(nor_379_nl, mux_1261_nl, fsm_output(2));
  nor_382_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1011")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_383_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) OR not_tmp_133);
  and_308_nl <= (VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("101")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4)));
  nor_384_nl <= NOT((NOT (z_out_6_10_1(0))) OR (z_out_6_10_1(2)) OR nand_260_cse_1);
  mux_1255_nl <= MUX_s_1_2_2(and_308_nl, nor_384_nl, fsm_output(0));
  mux_1256_nl <= MUX_s_1_2_2(nor_383_nl, mux_1255_nl, fsm_output(6));
  and_307_nl <= (fsm_output(1)) AND mux_1256_nl;
  mux_1257_nl <= MUX_s_1_2_2(nor_382_nl, and_307_nl, fsm_output(3));
  nor_385_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_386_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_1252_nl <= MUX_s_1_2_2(nor_385_nl, nor_386_nl, fsm_output(0));
  nor_388_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1251_nl <= MUX_s_1_2_2(nor_387_cse, nor_388_nl, fsm_output(0));
  mux_1253_nl <= MUX_s_1_2_2(mux_1252_nl, mux_1251_nl, fsm_output(6));
  nor_389_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  and_431_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011")) AND
      (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4));
  mux_1249_nl <= MUX_s_1_2_2(nor_389_nl, and_431_nl, fsm_output(0));
  nor_391_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1250_nl <= MUX_s_1_2_2(mux_1249_nl, nor_391_nl, fsm_output(6));
  mux_1254_nl <= MUX_s_1_2_2(mux_1253_nl, mux_1250_nl, fsm_output(1));
  and_309_nl <= (fsm_output(3)) AND mux_1254_nl;
  mux_1258_nl <= MUX_s_1_2_2(mux_1257_nl, and_309_nl, fsm_output(2));
  mux_1269_nl <= MUX_s_1_2_2(mux_1268_nl, mux_1258_nl, fsm_output(8));
  nor_394_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1245_nl <= MUX_s_1_2_2(nor_387_cse, nor_394_nl, fsm_output(0));
  nor_395_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_396_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1244_nl <= MUX_s_1_2_2(nor_395_nl, nor_396_nl, fsm_output(0));
  mux_1246_nl <= MUX_s_1_2_2(mux_1245_nl, mux_1244_nl, fsm_output(6));
  nor_397_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1011"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_1247_nl <= MUX_s_1_2_2(mux_1246_nl, nor_397_nl, fsm_output(1));
  nand_77_nl <= NOT((fsm_output(3)) AND mux_1247_nl);
  or_1375_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      AND (NOT (fsm_output(5))))) OR not_tmp_134;
  nand_248_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("101"))
      AND (VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5))
      AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_1372_nl <= (NOT (z_out_6_10_1(0))) OR (z_out_6_10_1(2)) OR nand_260_cse_1;
  mux_1241_nl <= MUX_s_1_2_2(nand_248_nl, or_1372_nl, fsm_output(0));
  nand_352_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5)) AND (NOT (fsm_output(7)))
      AND (fsm_output(4)));
  mux_1240_nl <= MUX_s_1_2_2(nand_241_cse, nand_352_nl, fsm_output(0));
  mux_1242_nl <= MUX_s_1_2_2(mux_1241_nl, mux_1240_nl, fsm_output(6));
  mux_1243_nl <= MUX_s_1_2_2(or_1375_nl, mux_1242_nl, fsm_output(1));
  or_1376_nl <= (fsm_output(3)) OR mux_1243_nl;
  mux_1248_nl <= MUX_s_1_2_2(nand_77_nl, or_1376_nl, fsm_output(2));
  nor_392_nl <= NOT((fsm_output(8)) OR mux_1248_nl);
  vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1269_nl, nor_392_nl,
      fsm_output(9));
  or_1465_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_1296_nl <= MUX_s_1_2_2(or_tmp_1403, or_1465_nl, fsm_output(0));
  or_1464_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1295_nl <= MUX_s_1_2_2(or_1464_nl, or_tmp_1395, fsm_output(0));
  mux_1297_nl <= MUX_s_1_2_2(mux_1296_nl, mux_1295_nl, fsm_output(4));
  nand_82_nl <= NOT((fsm_output(6)) AND (NOT mux_1297_nl));
  or_1463_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("00")) OR not_tmp_289;
  mux_1298_nl <= MUX_s_1_2_2(nand_82_nl, or_1463_nl, fsm_output(7));
  nor_373_nl <= NOT((fsm_output(8)) OR mux_1298_nl);
  and_436_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (NOT (VEC_LOOP_j_sva_9_0(0))) AND (NOT (fsm_output(5))) AND (fsm_output(1));
  or_1458_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1293_nl <= MUX_s_1_2_2(or_1458_nl, or_tmp_1403, fsm_output(0));
  nor_375_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_1293_nl);
  mux_1294_nl <= MUX_s_1_2_2(and_436_nl, nor_375_nl, fsm_output(8));
  mux_1299_nl <= MUX_s_1_2_2(nor_373_nl, mux_1294_nl, fsm_output(9));
  or_1455_nl <= CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0)))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_1453_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1288_nl <= MUX_s_1_2_2(or_1453_nl, or_tmp_1403, fsm_output(0));
  or_1451_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1287_nl <= MUX_s_1_2_2(or_tmp_1401, or_1451_nl, fsm_output(0));
  mux_1289_nl <= MUX_s_1_2_2(mux_1288_nl, mux_1287_nl, fsm_output(4));
  or_1449_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1286_nl <= MUX_s_1_2_2(or_1449_nl, or_tmp_1395, fsm_output(0));
  or_1450_nl <= (fsm_output(4)) OR mux_1286_nl;
  mux_1290_nl <= MUX_s_1_2_2(mux_1289_nl, or_1450_nl, fsm_output(6));
  mux_1291_nl <= MUX_s_1_2_2(or_1455_nl, mux_1290_nl, fsm_output(7));
  and_306_nl <= (fsm_output(8)) AND (NOT mux_1291_nl);
  nor_376_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_289);
  mux_1292_nl <= MUX_s_1_2_2(and_306_nl, nor_376_nl, fsm_output(9));
  mux_1300_nl <= MUX_s_1_2_2(mux_1299_nl, mux_1292_nl, fsm_output(3));
  or_1445_nl <= CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (VEC_LOOP_j_sva_9_0(0))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  or_1443_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1281_nl <= MUX_s_1_2_2(or_1443_nl, or_tmp_1403, fsm_output(0));
  or_1441_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1280_nl <= MUX_s_1_2_2(or_tmp_1401, or_1441_nl, fsm_output(0));
  mux_1282_nl <= MUX_s_1_2_2(mux_1281_nl, mux_1280_nl, fsm_output(4));
  mux_1283_nl <= MUX_s_1_2_2(or_1445_nl, mux_1282_nl, fsm_output(6));
  or_1439_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1278_nl <= MUX_s_1_2_2(or_1439_nl, or_tmp_1395, fsm_output(0));
  or_1440_nl <= (fsm_output(4)) OR mux_1278_nl;
  mux_1279_nl <= MUX_s_1_2_2(or_1440_nl, or_tmp_1393, fsm_output(6));
  mux_1284_nl <= MUX_s_1_2_2(mux_1283_nl, mux_1279_nl, fsm_output(7));
  nor_377_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1284_nl);
  or_1436_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (VEC_LOOP_j_sva_9_0(0)) OR (fsm_output(5))
      OR (NOT (fsm_output(1)));
  or_1434_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1274_nl <= MUX_s_1_2_2(or_1434_nl, or_tmp_1403, fsm_output(0));
  or_1428_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1273_nl <= MUX_s_1_2_2(or_tmp_1401, or_1428_nl, fsm_output(0));
  mux_1275_nl <= MUX_s_1_2_2(mux_1274_nl, mux_1273_nl, fsm_output(4));
  mux_1276_nl <= MUX_s_1_2_2(or_1436_nl, mux_1275_nl, fsm_output(6));
  nand_80_nl <= NOT((fsm_output(7)) AND (NOT mux_1276_nl));
  or_1425_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1271_nl <= MUX_s_1_2_2(or_1425_nl, or_tmp_1395, fsm_output(0));
  or_1426_nl <= (fsm_output(4)) OR mux_1271_nl;
  mux_1272_nl <= MUX_s_1_2_2(or_1426_nl, or_tmp_1393, fsm_output(6));
  or_1427_nl <= (fsm_output(7)) OR mux_1272_nl;
  mux_1277_nl <= MUX_s_1_2_2(nand_80_nl, or_1427_nl, fsm_output(8));
  nor_378_nl <= NOT((fsm_output(9)) OR mux_1277_nl);
  mux_1285_nl <= MUX_s_1_2_2(nor_377_nl, nor_378_nl, fsm_output(3));
  vec_rsc_0_12_i_we_d_pff <= MUX_s_1_2_2(mux_1300_nl, mux_1285_nl, fsm_output(2));
  nor_362_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  or_1515_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1518_nl <= (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1517_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_1327_nl <= MUX_s_1_2_2(or_1517_nl, or_1515_cse, fsm_output(0));
  mux_1328_nl <= MUX_s_1_2_2(or_1518_nl, mux_1327_nl, fsm_output(6));
  or_1514_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR not_tmp_133;
  or_1512_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_1325_nl <= MUX_s_1_2_2(or_1514_nl, or_1512_nl, fsm_output(0));
  or_1511_nl <= (VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1509_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1324_nl <= MUX_s_1_2_2(or_1511_nl, or_1509_nl, fsm_output(0));
  mux_1326_nl <= MUX_s_1_2_2(mux_1325_nl, mux_1324_nl, fsm_output(6));
  mux_1329_nl <= MUX_s_1_2_2(mux_1328_nl, mux_1326_nl, fsm_output(1));
  nor_353_nl <= NOT((fsm_output(3)) OR mux_1329_nl);
  or_1507_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1505_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_1321_nl <= MUX_s_1_2_2(or_1507_nl, or_1505_nl, fsm_output(0));
  or_1504_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1322_nl <= MUX_s_1_2_2(mux_1321_nl, or_1504_nl, fsm_output(6));
  nor_354_nl <= NOT((fsm_output(1)) OR mux_1322_nl);
  nor_355_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1100"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_1323_nl <= MUX_s_1_2_2(nor_354_nl, nor_355_nl, fsm_output(3));
  mux_1330_nl <= MUX_s_1_2_2(nor_353_nl, mux_1323_nl, fsm_output(2));
  nor_356_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1100")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_357_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR not_tmp_133);
  nor_358_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_359_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100"))
      OR nand_270_cse_1);
  mux_1317_nl <= MUX_s_1_2_2(nor_358_nl, nor_359_nl, fsm_output(0));
  mux_1318_nl <= MUX_s_1_2_2(nor_357_nl, mux_1317_nl, fsm_output(6));
  and_304_nl <= (fsm_output(1)) AND mux_1318_nl;
  mux_1319_nl <= MUX_s_1_2_2(nor_356_nl, and_304_nl, fsm_output(3));
  nor_360_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_361_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_1314_nl <= MUX_s_1_2_2(nor_360_nl, nor_361_nl, fsm_output(0));
  nor_363_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1313_nl <= MUX_s_1_2_2(nor_362_cse, nor_363_nl, fsm_output(0));
  mux_1315_nl <= MUX_s_1_2_2(mux_1314_nl, mux_1313_nl, fsm_output(6));
  nor_364_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  nor_365_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1311_nl <= MUX_s_1_2_2(nor_364_nl, nor_365_nl, fsm_output(0));
  nor_366_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1312_nl <= MUX_s_1_2_2(mux_1311_nl, nor_366_nl, fsm_output(6));
  mux_1316_nl <= MUX_s_1_2_2(mux_1315_nl, mux_1312_nl, fsm_output(1));
  and_305_nl <= (fsm_output(3)) AND mux_1316_nl;
  mux_1320_nl <= MUX_s_1_2_2(mux_1319_nl, and_305_nl, fsm_output(2));
  mux_1331_nl <= MUX_s_1_2_2(mux_1330_nl, mux_1320_nl, fsm_output(8));
  nor_369_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1307_nl <= MUX_s_1_2_2(nor_362_cse, nor_369_nl, fsm_output(0));
  nor_370_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_371_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1306_nl <= MUX_s_1_2_2(nor_370_nl, nor_371_nl, fsm_output(0));
  mux_1308_nl <= MUX_s_1_2_2(mux_1307_nl, mux_1306_nl, fsm_output(6));
  nor_372_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_1309_nl <= MUX_s_1_2_2(mux_1308_nl, nor_372_nl, fsm_output(1));
  nand_83_nl <= NOT((fsm_output(3)) AND mux_1309_nl);
  or_1474_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      OR (fsm_output(5)) OR not_tmp_134;
  or_1472_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR
      (NOT (fsm_output(5))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_1471_nl <= CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("100")) OR
      nand_270_cse_1;
  mux_1303_nl <= MUX_s_1_2_2(or_1472_nl, or_1471_nl, fsm_output(0));
  or_1468_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (NOT (fsm_output(4)));
  mux_1302_nl <= MUX_s_1_2_2(or_1515_cse, or_1468_nl, fsm_output(0));
  mux_1304_nl <= MUX_s_1_2_2(mux_1303_nl, mux_1302_nl, fsm_output(6));
  mux_1305_nl <= MUX_s_1_2_2(or_1474_nl, mux_1304_nl, fsm_output(1));
  or_1475_nl <= (fsm_output(3)) OR mux_1305_nl;
  mux_1310_nl <= MUX_s_1_2_2(nand_83_nl, or_1475_nl, fsm_output(2));
  nor_367_nl <= NOT((fsm_output(8)) OR mux_1310_nl);
  vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1331_nl, nor_367_nl,
      fsm_output(9));
  or_1565_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(1)) OR (fsm_output(5));
  mux_1358_nl <= MUX_s_1_2_2(or_tmp_1502, or_1565_nl, fsm_output(0));
  or_1564_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1357_nl <= MUX_s_1_2_2(or_1564_nl, or_tmp_1493, fsm_output(0));
  mux_1359_nl <= MUX_s_1_2_2(mux_1358_nl, mux_1357_nl, fsm_output(4));
  nor_346_nl <= NOT((fsm_output(9)) OR (NOT (fsm_output(6))) OR mux_1359_nl);
  nand_230_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (fsm_output(4)) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0)) AND (fsm_output(1))
      AND (NOT (fsm_output(5))));
  or_1561_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1354_nl <= MUX_s_1_2_2(or_1561_nl, or_tmp_1502, fsm_output(0));
  or_1560_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1353_nl <= MUX_s_1_2_2(or_tmp_1500, or_1560_nl, fsm_output(0));
  mux_1355_nl <= MUX_s_1_2_2(mux_1354_nl, mux_1353_nl, fsm_output(4));
  mux_1356_nl <= MUX_s_1_2_2(nand_230_nl, mux_1355_nl, fsm_output(6));
  and_302_nl <= (fsm_output(9)) AND (NOT mux_1356_nl);
  mux_1360_nl <= MUX_s_1_2_2(nor_346_nl, and_302_nl, fsm_output(2));
  or_1557_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1352_nl <= MUX_s_1_2_2(or_1557_nl, or_tmp_1502, fsm_output(0));
  nor_347_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR
      (fsm_output(4)) OR mux_1352_nl);
  mux_1361_nl <= MUX_s_1_2_2(mux_1360_nl, nor_347_nl, fsm_output(8));
  or_1554_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(1))
      OR (NOT (fsm_output(5))) OR (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1)) OR not_tmp_304;
  nand_231_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0))
      AND (fsm_output(1)) AND (NOT (fsm_output(5))));
  mux_1350_nl <= MUX_s_1_2_2(or_1554_nl, nand_231_nl, fsm_output(9));
  or_1550_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1348_nl <= MUX_s_1_2_2(or_1550_nl, or_tmp_1493, fsm_output(0));
  or_1551_nl <= (fsm_output(4)) OR mux_1348_nl;
  mux_1349_nl <= MUX_s_1_2_2(or_1551_nl, or_tmp_1512, fsm_output(6));
  nand_86_nl <= NOT((fsm_output(9)) AND (NOT mux_1349_nl));
  mux_1351_nl <= MUX_s_1_2_2(mux_1350_nl, nand_86_nl, fsm_output(2));
  nor_348_nl <= NOT((fsm_output(8)) OR mux_1351_nl);
  mux_1362_nl <= MUX_s_1_2_2(mux_1361_nl, nor_348_nl, fsm_output(7));
  nor_349_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(9))) OR (fsm_output(6)) OR
      (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(5))
      OR (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1)) OR not_tmp_304);
  and_303_nl <= (NOT (fsm_output(9))) AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("110")) AND (fsm_output(6)) AND (fsm_output(4))
      AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0)) AND (fsm_output(1)) AND (NOT
      (fsm_output(5)));
  or_1543_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1343_nl <= MUX_s_1_2_2(or_1543_nl, or_tmp_1493, fsm_output(0));
  or_1544_nl <= (fsm_output(4)) OR mux_1343_nl;
  mux_1344_nl <= MUX_s_1_2_2(or_1544_nl, or_tmp_1512, fsm_output(6));
  nor_350_nl <= NOT((fsm_output(9)) OR mux_1344_nl);
  mux_1345_nl <= MUX_s_1_2_2(and_303_nl, nor_350_nl, fsm_output(2));
  mux_1346_nl <= MUX_s_1_2_2(nor_349_nl, mux_1345_nl, fsm_output(8));
  nand_232_nl <= NOT((fsm_output(4)) AND (fsm_output(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("110")) AND (VEC_LOOP_j_sva_9_0(0)) AND (fsm_output(1))
      AND (NOT (fsm_output(5))));
  or_1537_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1339_nl <= MUX_s_1_2_2(or_1537_nl, or_tmp_1502, fsm_output(0));
  or_1536_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1338_nl <= MUX_s_1_2_2(or_tmp_1500, or_1536_nl, fsm_output(0));
  mux_1340_nl <= MUX_s_1_2_2(mux_1339_nl, mux_1338_nl, fsm_output(4));
  mux_1341_nl <= MUX_s_1_2_2(nand_232_nl, mux_1340_nl, fsm_output(6));
  nor_351_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(9)) OR mux_1341_nl);
  or_1532_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(1))) OR (fsm_output(5));
  mux_1335_nl <= MUX_s_1_2_2(or_1532_nl, or_tmp_1502, fsm_output(0));
  or_1527_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1334_nl <= MUX_s_1_2_2(or_tmp_1500, or_1527_nl, fsm_output(0));
  mux_1336_nl <= MUX_s_1_2_2(mux_1335_nl, mux_1334_nl, fsm_output(4));
  or_1524_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_1333_nl <= MUX_s_1_2_2(or_1524_nl, or_tmp_1493, fsm_output(0));
  or_1525_nl <= (fsm_output(4)) OR mux_1333_nl;
  mux_1337_nl <= MUX_s_1_2_2(mux_1336_nl, or_1525_nl, fsm_output(6));
  nor_352_nl <= NOT((fsm_output(2)) OR (fsm_output(9)) OR mux_1337_nl);
  mux_1342_nl <= MUX_s_1_2_2(nor_351_nl, nor_352_nl, fsm_output(8));
  mux_1347_nl <= MUX_s_1_2_2(mux_1346_nl, mux_1342_nl, fsm_output(7));
  vec_rsc_0_13_i_we_d_pff <= MUX_s_1_2_2(mux_1362_nl, mux_1347_nl, fsm_output(3));
  nor_335_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nand_217_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  nand_216_nl <= NOT((fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND
      CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_1615_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_1389_nl <= MUX_s_1_2_2(or_1615_nl, nand_217_cse, fsm_output(0));
  mux_1390_nl <= MUX_s_1_2_2(nand_216_nl, mux_1389_nl, fsm_output(6));
  or_1612_nl <= (z_out_6_10_1(1)) OR (NOT((z_out_6_10_1(2)) AND (z_out_6_10_1(3))
      AND (z_out_6_10_1(0)) AND (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(4))));
  or_1611_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_1387_nl <= MUX_s_1_2_2(or_1612_nl, or_1611_nl, fsm_output(0));
  nand_368_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("110")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4)));
  or_1608_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1386_nl <= MUX_s_1_2_2(nand_368_nl, or_1608_nl, fsm_output(0));
  mux_1388_nl <= MUX_s_1_2_2(mux_1387_nl, mux_1386_nl, fsm_output(6));
  mux_1391_nl <= MUX_s_1_2_2(mux_1390_nl, mux_1388_nl, fsm_output(1));
  nor_327_nl <= NOT((fsm_output(3)) OR mux_1391_nl);
  or_1606_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1604_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_1383_nl <= MUX_s_1_2_2(or_1606_nl, or_1604_nl, fsm_output(0));
  or_1603_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1384_nl <= MUX_s_1_2_2(mux_1383_nl, or_1603_nl, fsm_output(6));
  nor_328_nl <= NOT((fsm_output(1)) OR mux_1384_nl);
  nor_329_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_1385_nl <= MUX_s_1_2_2(nor_328_nl, nor_329_nl, fsm_output(3));
  mux_1392_nl <= MUX_s_1_2_2(nor_327_nl, mux_1385_nl, fsm_output(2));
  nor_330_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1101")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_331_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) OR not_tmp_133);
  and_300_nl <= (VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("110")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4)));
  nor_332_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101"))
      OR nand_270_cse_1);
  mux_1379_nl <= MUX_s_1_2_2(and_300_nl, nor_332_nl, fsm_output(0));
  mux_1380_nl <= MUX_s_1_2_2(nor_331_nl, mux_1379_nl, fsm_output(6));
  and_299_nl <= (fsm_output(1)) AND mux_1380_nl;
  mux_1381_nl <= MUX_s_1_2_2(nor_330_nl, and_299_nl, fsm_output(3));
  nor_333_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_334_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_1376_nl <= MUX_s_1_2_2(nor_333_nl, nor_334_nl, fsm_output(0));
  nor_336_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1375_nl <= MUX_s_1_2_2(nor_335_cse, nor_336_nl, fsm_output(0));
  mux_1377_nl <= MUX_s_1_2_2(mux_1376_nl, mux_1375_nl, fsm_output(6));
  nor_337_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  and_430_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101")) AND
      (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4));
  mux_1373_nl <= MUX_s_1_2_2(nor_337_nl, and_430_nl, fsm_output(0));
  nor_339_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1374_nl <= MUX_s_1_2_2(mux_1373_nl, nor_339_nl, fsm_output(6));
  mux_1378_nl <= MUX_s_1_2_2(mux_1377_nl, mux_1374_nl, fsm_output(1));
  and_301_nl <= (fsm_output(3)) AND mux_1378_nl;
  mux_1382_nl <= MUX_s_1_2_2(mux_1381_nl, and_301_nl, fsm_output(2));
  mux_1393_nl <= MUX_s_1_2_2(mux_1392_nl, mux_1382_nl, fsm_output(8));
  nor_342_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1369_nl <= MUX_s_1_2_2(nor_335_cse, nor_342_nl, fsm_output(0));
  nor_343_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_344_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1368_nl <= MUX_s_1_2_2(nor_343_nl, nor_344_nl, fsm_output(0));
  mux_1370_nl <= MUX_s_1_2_2(mux_1369_nl, mux_1368_nl, fsm_output(6));
  nor_345_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1101"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_1371_nl <= MUX_s_1_2_2(mux_1370_nl, nor_345_nl, fsm_output(1));
  nand_89_nl <= NOT((fsm_output(3)) AND mux_1371_nl);
  or_1573_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      AND (NOT (fsm_output(5))))) OR not_tmp_134;
  nand_224_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("110"))
      AND (VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5))
      AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_1570_nl <= CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101")) OR
      nand_270_cse_1;
  mux_1365_nl <= MUX_s_1_2_2(nand_224_nl, or_1570_nl, fsm_output(0));
  nand_351_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5)) AND (NOT (fsm_output(7)))
      AND (fsm_output(4)));
  mux_1364_nl <= MUX_s_1_2_2(nand_217_cse, nand_351_nl, fsm_output(0));
  mux_1366_nl <= MUX_s_1_2_2(mux_1365_nl, mux_1364_nl, fsm_output(6));
  mux_1367_nl <= MUX_s_1_2_2(or_1573_nl, mux_1366_nl, fsm_output(1));
  or_1574_nl <= (fsm_output(3)) OR mux_1367_nl;
  mux_1372_nl <= MUX_s_1_2_2(nand_89_nl, or_1574_nl, fsm_output(2));
  nor_340_nl <= NOT((fsm_output(8)) OR mux_1372_nl);
  vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1393_nl, nor_340_nl,
      fsm_output(9));
  or_1662_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_1420_nl <= MUX_s_1_2_2(or_tmp_1600, or_1662_nl, fsm_output(0));
  or_1661_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1419_nl <= MUX_s_1_2_2(or_1661_nl, or_tmp_1592, fsm_output(0));
  mux_1421_nl <= MUX_s_1_2_2(mux_1420_nl, mux_1419_nl, fsm_output(4));
  nand_94_nl <= NOT((fsm_output(6)) AND (NOT mux_1421_nl));
  or_1660_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("10")) OR not_tmp_289;
  mux_1422_nl <= MUX_s_1_2_2(nand_94_nl, or_1660_nl, fsm_output(7));
  nor_321_nl <= NOT((fsm_output(8)) OR mux_1422_nl);
  and_435_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (NOT (VEC_LOOP_j_sva_9_0(0))) AND (NOT (fsm_output(5))) AND (fsm_output(1));
  or_1655_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1417_nl <= MUX_s_1_2_2(or_1655_nl, or_tmp_1600, fsm_output(0));
  nor_323_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_1417_nl);
  mux_1418_nl <= MUX_s_1_2_2(and_435_nl, nor_323_nl, fsm_output(8));
  mux_1423_nl <= MUX_s_1_2_2(nor_321_nl, mux_1418_nl, fsm_output(9));
  nand_375_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0)) AND (NOT (VEC_LOOP_j_sva_9_0(0)))
      AND (NOT (fsm_output(5))) AND (fsm_output(1)));
  or_1650_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1412_nl <= MUX_s_1_2_2(or_1650_nl, or_tmp_1600, fsm_output(0));
  or_1648_nl <= (NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1411_nl <= MUX_s_1_2_2(or_tmp_1598, or_1648_nl, fsm_output(0));
  mux_1413_nl <= MUX_s_1_2_2(mux_1412_nl, mux_1411_nl, fsm_output(4));
  or_1646_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1410_nl <= MUX_s_1_2_2(or_1646_nl, or_tmp_1592, fsm_output(0));
  or_1647_nl <= (fsm_output(4)) OR mux_1410_nl;
  mux_1414_nl <= MUX_s_1_2_2(mux_1413_nl, or_1647_nl, fsm_output(6));
  mux_1415_nl <= MUX_s_1_2_2(nand_375_nl, mux_1414_nl, fsm_output(7));
  and_298_nl <= (fsm_output(8)) AND (NOT mux_1415_nl);
  nor_324_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      CONV_SL_1_1(COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"))
      OR not_tmp_289);
  mux_1416_nl <= MUX_s_1_2_2(and_298_nl, nor_324_nl, fsm_output(9));
  mux_1424_nl <= MUX_s_1_2_2(mux_1423_nl, mux_1416_nl, fsm_output(3));
  nand_367_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(4)) AND (fsm_output(0)) AND (NOT (VEC_LOOP_j_sva_9_0(0))) AND
      (NOT (fsm_output(5))) AND (fsm_output(1)));
  or_1640_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1405_nl <= MUX_s_1_2_2(or_1640_nl, or_tmp_1600, fsm_output(0));
  or_1638_nl <= CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1404_nl <= MUX_s_1_2_2(or_tmp_1598, or_1638_nl, fsm_output(0));
  mux_1406_nl <= MUX_s_1_2_2(mux_1405_nl, mux_1404_nl, fsm_output(4));
  mux_1407_nl <= MUX_s_1_2_2(nand_367_nl, mux_1406_nl, fsm_output(6));
  or_1636_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1402_nl <= MUX_s_1_2_2(or_1636_nl, or_tmp_1592, fsm_output(0));
  or_1637_nl <= (fsm_output(4)) OR mux_1402_nl;
  mux_1403_nl <= MUX_s_1_2_2(or_1637_nl, or_tmp_1590, fsm_output(6));
  mux_1408_nl <= MUX_s_1_2_2(mux_1407_nl, mux_1403_nl, fsm_output(7));
  nor_325_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1408_nl);
  nand_359_nl <= NOT((fsm_output(4)) AND (fsm_output(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (NOT (VEC_LOOP_j_sva_9_0(0))) AND (NOT
      (fsm_output(5))) AND (fsm_output(1)));
  or_1631_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_1398_nl <= MUX_s_1_2_2(or_1631_nl, or_tmp_1600, fsm_output(0));
  or_1625_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1397_nl <= MUX_s_1_2_2(or_tmp_1598, or_1625_nl, fsm_output(0));
  mux_1399_nl <= MUX_s_1_2_2(mux_1398_nl, mux_1397_nl, fsm_output(4));
  mux_1400_nl <= MUX_s_1_2_2(nand_359_nl, mux_1399_nl, fsm_output(6));
  nand_92_nl <= NOT((fsm_output(7)) AND (NOT mux_1400_nl));
  or_1622_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_1395_nl <= MUX_s_1_2_2(or_1622_nl, or_tmp_1592, fsm_output(0));
  or_1623_nl <= (fsm_output(4)) OR mux_1395_nl;
  mux_1396_nl <= MUX_s_1_2_2(or_1623_nl, or_tmp_1590, fsm_output(6));
  or_1624_nl <= (fsm_output(7)) OR mux_1396_nl;
  mux_1401_nl <= MUX_s_1_2_2(nand_92_nl, or_1624_nl, fsm_output(8));
  nor_326_nl <= NOT((fsm_output(9)) OR mux_1401_nl);
  mux_1409_nl <= MUX_s_1_2_2(nor_325_nl, nor_326_nl, fsm_output(3));
  vec_rsc_0_14_i_we_d_pff <= MUX_s_1_2_2(mux_1424_nl, mux_1409_nl, fsm_output(2));
  nor_310_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nand_202_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(4)));
  nand_197_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  nand_196_nl <= NOT((fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND
      CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_1712_nl <= CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR not_tmp_134;
  mux_1451_nl <= MUX_s_1_2_2(or_1712_nl, nand_197_cse, fsm_output(0));
  mux_1452_nl <= MUX_s_1_2_2(nand_196_nl, mux_1451_nl, fsm_output(6));
  or_1709_nl <= (NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))))
      OR not_tmp_133;
  or_1707_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  mux_1449_nl <= MUX_s_1_2_2(or_1709_nl, or_1707_nl, fsm_output(0));
  nand_366_nl <= NOT((NOT (VEC_LOOP_j_sva_9_0(0))) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4)));
  or_1704_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1448_nl <= MUX_s_1_2_2(nand_366_nl, or_1704_nl, fsm_output(0));
  mux_1450_nl <= MUX_s_1_2_2(mux_1449_nl, mux_1448_nl, fsm_output(6));
  mux_1453_nl <= MUX_s_1_2_2(mux_1452_nl, mux_1450_nl, fsm_output(1));
  nor_302_nl <= NOT((fsm_output(3)) OR mux_1453_nl);
  or_1702_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  or_1700_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4));
  mux_1445_nl <= MUX_s_1_2_2(or_1702_nl, or_1700_nl, fsm_output(0));
  or_1699_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1446_nl <= MUX_s_1_2_2(mux_1445_nl, or_1699_nl, fsm_output(6));
  nor_303_nl <= NOT((fsm_output(1)) OR mux_1446_nl);
  nor_304_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_1447_nl <= MUX_s_1_2_2(nor_303_nl, nor_304_nl, fsm_output(3));
  mux_1454_nl <= MUX_s_1_2_2(nor_302_nl, mux_1447_nl, fsm_output(2));
  nor_305_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1110")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_306_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) OR not_tmp_133);
  and_296_nl <= (NOT (VEC_LOOP_j_sva_9_0(0))) AND CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4)));
  nor_307_nl <= NOT((z_out_6_10_1(0)) OR nand_202_cse);
  mux_1441_nl <= MUX_s_1_2_2(and_296_nl, nor_307_nl, fsm_output(0));
  mux_1442_nl <= MUX_s_1_2_2(nor_306_nl, mux_1441_nl, fsm_output(6));
  and_295_nl <= (fsm_output(1)) AND mux_1442_nl;
  mux_1443_nl <= MUX_s_1_2_2(nor_305_nl, and_295_nl, fsm_output(3));
  nor_308_nl <= NOT((NOT (COMP_LOOP_acc_16_psp_sva(0))) OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("110")) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR (fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(4)));
  nor_309_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR not_tmp_134);
  mux_1438_nl <= MUX_s_1_2_2(nor_308_nl, nor_309_nl, fsm_output(0));
  nor_311_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1437_nl <= MUX_s_1_2_2(nor_310_cse, nor_311_nl, fsm_output(0));
  mux_1439_nl <= MUX_s_1_2_2(mux_1438_nl, mux_1437_nl, fsm_output(6));
  nor_312_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      OR CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("111"))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  and_429_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110")) AND
      (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4));
  mux_1435_nl <= MUX_s_1_2_2(nor_312_nl, and_429_nl, fsm_output(0));
  nor_314_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1436_nl <= MUX_s_1_2_2(mux_1435_nl, nor_314_nl, fsm_output(6));
  mux_1440_nl <= MUX_s_1_2_2(mux_1439_nl, mux_1436_nl, fsm_output(1));
  and_297_nl <= (fsm_output(3)) AND mux_1440_nl;
  mux_1444_nl <= MUX_s_1_2_2(mux_1443_nl, and_297_nl, fsm_output(2));
  mux_1455_nl <= MUX_s_1_2_2(mux_1454_nl, mux_1444_nl, fsm_output(8));
  nor_317_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  mux_1431_nl <= MUX_s_1_2_2(nor_310_cse, nor_317_nl, fsm_output(0));
  nor_318_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  nor_319_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4))));
  mux_1430_nl <= MUX_s_1_2_2(nor_318_nl, nor_319_nl, fsm_output(0));
  mux_1432_nl <= MUX_s_1_2_2(mux_1431_nl, mux_1430_nl, fsm_output(6));
  nor_320_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1110"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_1433_nl <= MUX_s_1_2_2(mux_1432_nl, nor_320_nl, fsm_output(1));
  nand_95_nl <= NOT((fsm_output(3)) AND mux_1433_nl);
  or_1670_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      AND (NOT (fsm_output(5))))) OR not_tmp_134;
  nand_204_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (NOT (VEC_LOOP_j_sva_9_0(0))) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_1667_nl <= (z_out_6_10_1(0)) OR nand_202_cse;
  mux_1427_nl <= MUX_s_1_2_2(nand_204_nl, or_1667_nl, fsm_output(0));
  nand_350_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5)) AND (NOT (fsm_output(7)))
      AND (fsm_output(4)));
  mux_1426_nl <= MUX_s_1_2_2(nand_197_cse, nand_350_nl, fsm_output(0));
  mux_1428_nl <= MUX_s_1_2_2(mux_1427_nl, mux_1426_nl, fsm_output(6));
  mux_1429_nl <= MUX_s_1_2_2(or_1670_nl, mux_1428_nl, fsm_output(1));
  or_1671_nl <= (fsm_output(3)) OR mux_1429_nl;
  mux_1434_nl <= MUX_s_1_2_2(nand_95_nl, or_1671_nl, fsm_output(2));
  nor_315_nl <= NOT((fsm_output(8)) OR mux_1434_nl);
  vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1455_nl, nor_315_nl,
      fsm_output(9));
  or_1756_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(5)) OR (fsm_output(1));
  mux_1482_nl <= MUX_s_1_2_2(or_tmp_1694, or_1756_nl, fsm_output(0));
  nand_178_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(5)) AND (NOT (fsm_output(1))));
  mux_1481_nl <= MUX_s_1_2_2(nand_178_nl, or_tmp_1689, fsm_output(0));
  mux_1483_nl <= MUX_s_1_2_2(mux_1482_nl, mux_1481_nl, fsm_output(4));
  nand_100_nl <= NOT((fsm_output(6)) AND (NOT mux_1483_nl));
  or_1754_nl <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(5)))
      OR (fsm_output(1)) OR not_tmp_335;
  mux_1484_nl <= MUX_s_1_2_2(nand_100_nl, or_1754_nl, fsm_output(7));
  nor_296_nl <= NOT((fsm_output(8)) OR mux_1484_nl);
  and_434_nl <= CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(7)) AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT (fsm_output(5))) AND (fsm_output(1));
  nand_377_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(5))) AND (fsm_output(1)));
  mux_1479_nl <= MUX_s_1_2_2(nand_377_nl, or_tmp_1694, fsm_output(0));
  nor_298_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(4)) OR mux_1479_nl);
  mux_1480_nl <= MUX_s_1_2_2(and_434_nl, nor_298_nl, fsm_output(8));
  mux_1485_nl <= MUX_s_1_2_2(nor_296_nl, mux_1480_nl, fsm_output(9));
  nand_374_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0))
      AND (NOT (fsm_output(5))) AND (fsm_output(1)));
  nand_372_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(5))) AND (fsm_output(1)));
  mux_1474_nl <= MUX_s_1_2_2(nand_372_nl, or_tmp_1694, fsm_output(0));
  nand_183_nl <= NOT((COMP_LOOP_acc_16_psp_sva(0)) AND CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (fsm_output(5)) AND (NOT (fsm_output(1))));
  mux_1473_nl <= MUX_s_1_2_2(not_tmp_336, nand_183_nl, fsm_output(0));
  mux_1475_nl <= MUX_s_1_2_2(mux_1474_nl, mux_1473_nl, fsm_output(4));
  nand_184_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(5)) AND (NOT (fsm_output(1))));
  mux_1472_nl <= MUX_s_1_2_2(nand_184_nl, or_tmp_1689, fsm_output(0));
  or_1741_nl <= (fsm_output(4)) OR mux_1472_nl;
  mux_1476_nl <= MUX_s_1_2_2(mux_1475_nl, or_1741_nl, fsm_output(6));
  mux_1477_nl <= MUX_s_1_2_2(nand_374_nl, mux_1476_nl, fsm_output(7));
  and_294_nl <= (fsm_output(8)) AND (NOT mux_1477_nl);
  nor_299_nl <= NOT((fsm_output(8)) OR (fsm_output(7)) OR (fsm_output(6)) OR (NOT
      (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(5)) OR (fsm_output(1)) OR
      not_tmp_335);
  mux_1478_nl <= MUX_s_1_2_2(and_294_nl, nor_299_nl, fsm_output(9));
  mux_1486_nl <= MUX_s_1_2_2(mux_1485_nl, mux_1478_nl, fsm_output(3));
  nand_365_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(4)) AND (fsm_output(0)) AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT
      (fsm_output(5))) AND (fsm_output(1)));
  nand_362_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(5))) AND (fsm_output(1)));
  mux_1467_nl <= MUX_s_1_2_2(nand_362_nl, or_tmp_1694, fsm_output(0));
  nand_187_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      (fsm_output(5)) AND (NOT (fsm_output(1))));
  mux_1466_nl <= MUX_s_1_2_2(not_tmp_336, nand_187_nl, fsm_output(0));
  mux_1468_nl <= MUX_s_1_2_2(mux_1467_nl, mux_1466_nl, fsm_output(4));
  mux_1469_nl <= MUX_s_1_2_2(nand_365_nl, mux_1468_nl, fsm_output(6));
  nand_188_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(5)) AND (NOT (fsm_output(1))));
  mux_1464_nl <= MUX_s_1_2_2(nand_188_nl, or_tmp_1689, fsm_output(0));
  or_1731_nl <= (fsm_output(4)) OR mux_1464_nl;
  mux_1465_nl <= MUX_s_1_2_2(or_1731_nl, or_tmp_1687, fsm_output(6));
  mux_1470_nl <= MUX_s_1_2_2(mux_1469_nl, mux_1465_nl, fsm_output(7));
  nor_300_nl <= NOT(CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"))
      OR mux_1470_nl);
  nand_358_nl <= NOT((fsm_output(4)) AND (fsm_output(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND (VEC_LOOP_j_sva_9_0(0)) AND (NOT (fsm_output(5)))
      AND (fsm_output(1)));
  nand_349_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(5))) AND (fsm_output(1)));
  mux_1460_nl <= MUX_s_1_2_2(nand_349_nl, or_tmp_1694, fsm_output(0));
  nand_191_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      (fsm_output(5)) AND (NOT (fsm_output(1))));
  mux_1459_nl <= MUX_s_1_2_2(not_tmp_336, nand_191_nl, fsm_output(0));
  mux_1461_nl <= MUX_s_1_2_2(mux_1460_nl, mux_1459_nl, fsm_output(4));
  mux_1462_nl <= MUX_s_1_2_2(nand_358_nl, mux_1461_nl, fsm_output(6));
  nand_98_nl <= NOT((fsm_output(7)) AND (NOT mux_1462_nl));
  nand_192_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(5)) AND (NOT (fsm_output(1))));
  mux_1457_nl <= MUX_s_1_2_2(nand_192_nl, or_tmp_1689, fsm_output(0));
  or_1720_nl <= (fsm_output(4)) OR mux_1457_nl;
  mux_1458_nl <= MUX_s_1_2_2(or_1720_nl, or_tmp_1687, fsm_output(6));
  or_1721_nl <= (fsm_output(7)) OR mux_1458_nl;
  mux_1463_nl <= MUX_s_1_2_2(nand_98_nl, or_1721_nl, fsm_output(8));
  nor_301_nl <= NOT((fsm_output(9)) OR mux_1463_nl);
  mux_1471_nl <= MUX_s_1_2_2(nor_300_nl, nor_301_nl, fsm_output(3));
  vec_rsc_0_15_i_we_d_pff <= MUX_s_1_2_2(mux_1486_nl, mux_1471_nl, fsm_output(2));
  and_291_cse <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(5))) AND (fsm_output(7)) AND (NOT (fsm_output(4)));
  nand_161_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(4)));
  nand_160_cse <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  nand_158_nl <= NOT((fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND
      CONV_SL_1_1(COMP_LOOP_acc_1_cse_4_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  or_1802_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_13_psp_sva(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (NOT (fsm_output(5))))) OR not_tmp_134;
  mux_1513_nl <= MUX_s_1_2_2(or_1802_nl, nand_160_cse, fsm_output(0));
  mux_1514_nl <= MUX_s_1_2_2(nand_158_nl, mux_1513_nl, fsm_output(6));
  nand_162_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(5))) AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  mux_1511_nl <= MUX_s_1_2_2(nand_161_cse, nand_162_nl, fsm_output(0));
  nand_364_nl <= NOT((VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_11_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4)));
  or_1796_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4));
  mux_1510_nl <= MUX_s_1_2_2(nand_364_nl, or_1796_nl, fsm_output(0));
  mux_1512_nl <= MUX_s_1_2_2(mux_1511_nl, mux_1510_nl, fsm_output(6));
  mux_1515_nl <= MUX_s_1_2_2(mux_1514_nl, mux_1512_nl, fsm_output(1));
  nor_282_nl <= NOT((fsm_output(3)) OR mux_1515_nl);
  nand_361_nl <= NOT(CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(5))) AND (NOT (fsm_output(7))) AND (fsm_output(4)));
  nand_164_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(5)) AND (NOT (fsm_output(7))) AND (NOT (fsm_output(4))));
  mux_1507_nl <= MUX_s_1_2_2(nand_361_nl, nand_164_nl, fsm_output(0));
  or_1791_nl <= (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(5)) OR (fsm_output(7)) OR (NOT (fsm_output(4)));
  mux_1508_nl <= MUX_s_1_2_2(mux_1507_nl, or_1791_nl, fsm_output(6));
  nor_283_nl <= NOT((fsm_output(1)) OR mux_1508_nl);
  nor_284_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_6_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm))
      OR not_tmp_133);
  mux_1509_nl <= MUX_s_1_2_2(nor_283_nl, nor_284_nl, fsm_output(3));
  mux_1516_nl <= MUX_s_1_2_2(nor_282_nl, mux_1509_nl, fsm_output(2));
  nor_285_nl <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(0)) OR CONV_SL_1_1(z_out_6_10_1(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("1111")) OR (fsm_output(5)) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_286_nl <= NOT((NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_10_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)) OR not_tmp_133);
  and_287_nl <= (VEC_LOOP_j_sva_9_0(0)) AND CONV_SL_1_1(COMP_LOOP_acc_17_psp_sva(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (fsm_output(5)) AND (fsm_output(7)) AND (NOT (fsm_output(4)));
  and_288_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND
      (fsm_output(5)) AND (fsm_output(7)) AND (fsm_output(4));
  mux_1503_nl <= MUX_s_1_2_2(and_287_nl, and_288_nl, fsm_output(0));
  mux_1504_nl <= MUX_s_1_2_2(nor_286_nl, mux_1503_nl, fsm_output(6));
  and_286_nl <= (fsm_output(1)) AND mux_1504_nl;
  mux_1505_nl <= MUX_s_1_2_2(nor_285_nl, and_286_nl, fsm_output(3));
  and_290_nl <= (COMP_LOOP_acc_16_psp_sva(0)) AND CONV_SL_1_1(VEC_LOOP_j_sva_9_0(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND (NOT (fsm_output(5))) AND (fsm_output(7)) AND (NOT (fsm_output(4)));
  nor_287_nl <= NOT((NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (NOT (fsm_output(5))))) OR not_tmp_134);
  mux_1500_nl <= MUX_s_1_2_2(and_290_nl, nor_287_nl, fsm_output(0));
  and_427_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_8_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(5))) AND (NOT
      (fsm_output(7))) AND (fsm_output(4));
  mux_1499_nl <= MUX_s_1_2_2(and_291_cse, and_427_nl, fsm_output(0));
  mux_1501_nl <= MUX_s_1_2_2(mux_1500_nl, mux_1499_nl, fsm_output(6));
  and_292_nl <= (VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      AND CONV_SL_1_1(COMP_LOOP_acc_14_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(5)) AND (NOT (fsm_output(7))) AND (NOT (fsm_output(4)));
  and_428_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND
      (fsm_output(5)) AND (NOT (fsm_output(7))) AND (fsm_output(4));
  mux_1497_nl <= MUX_s_1_2_2(and_292_nl, and_428_nl, fsm_output(0));
  nor_290_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(4)));
  mux_1498_nl <= MUX_s_1_2_2(mux_1497_nl, nor_290_nl, fsm_output(6));
  mux_1502_nl <= MUX_s_1_2_2(mux_1501_nl, mux_1498_nl, fsm_output(1));
  and_289_nl <= (fsm_output(3)) AND mux_1502_nl;
  mux_1506_nl <= MUX_s_1_2_2(mux_1505_nl, and_289_nl, fsm_output(2));
  mux_1517_nl <= MUX_s_1_2_2(mux_1516_nl, mux_1506_nl, fsm_output(8));
  and_433_nl <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_12_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm AND (NOT (fsm_output(5))) AND (NOT
      (fsm_output(7))) AND (fsm_output(4));
  mux_1493_nl <= MUX_s_1_2_2(and_291_cse, and_433_nl, fsm_output(0));
  nor_293_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_19_psp_sva(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(VEC_LOOP_j_sva_9_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR
      (NOT COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) OR (fsm_output(5)) OR (fsm_output(7))
      OR (fsm_output(4)));
  and_440_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111")) AND
      (NOT (fsm_output(5))) AND (NOT (fsm_output(7))) AND (fsm_output(4));
  mux_1492_nl <= MUX_s_1_2_2(nor_293_nl, and_440_nl, fsm_output(0));
  mux_1494_nl <= MUX_s_1_2_2(mux_1493_nl, mux_1492_nl, fsm_output(6));
  nor_295_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1111"))
      OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR (fsm_output(4)));
  mux_1495_nl <= MUX_s_1_2_2(mux_1494_nl, nor_295_nl, fsm_output(1));
  nand_101_nl <= NOT((fsm_output(3)) AND mux_1495_nl);
  or_1763_nl <= (NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND (fsm_output(6)) AND (fsm_output(0)) AND COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      AND (NOT (fsm_output(5))))) OR not_tmp_134;
  nand_172_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_20_psp_sva(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"))
      AND (VEC_LOOP_j_sva_9_0(0)) AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5))
      AND (fsm_output(7)) AND (NOT (fsm_output(4))));
  mux_1489_nl <= MUX_s_1_2_2(nand_172_nl, nand_161_cse, fsm_output(0));
  nand_348_nl <= NOT(CONV_SL_1_1(COMP_LOOP_acc_1_cse_14_sva(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))
      AND COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm AND (fsm_output(5)) AND (NOT (fsm_output(7)))
      AND (fsm_output(4)));
  mux_1488_nl <= MUX_s_1_2_2(nand_160_cse, nand_348_nl, fsm_output(0));
  mux_1490_nl <= MUX_s_1_2_2(mux_1489_nl, mux_1488_nl, fsm_output(6));
  mux_1491_nl <= MUX_s_1_2_2(or_1763_nl, mux_1490_nl, fsm_output(1));
  or_1764_nl <= (fsm_output(3)) OR mux_1491_nl;
  mux_1496_nl <= MUX_s_1_2_2(nand_101_nl, or_1764_nl, fsm_output(2));
  nor_291_nl <= NOT((fsm_output(8)) OR mux_1496_nl);
  vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d <= MUX_s_1_2_2(mux_1517_nl, nor_291_nl,
      fsm_output(9));
  or_2213_nl <= (fsm_output(0)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(3))) OR (NOT (fsm_output(8))) OR (fsm_output(9));
  mux_2057_nl <= MUX_s_1_2_2(or_1977_cse, or_279_cse, fsm_output(0));
  mux_tmp_2006 <= MUX_s_1_2_2(or_2213_nl, mux_2057_nl, fsm_output(4));
  or_2219_nl <= (fsm_output(4)) OR (NOT (fsm_output(0))) OR (fsm_output(7)) OR (fsm_output(2))
      OR (fsm_output(3)) OR (NOT (fsm_output(8))) OR (fsm_output(9));
  or_2218_nl <= (fsm_output(0)) OR (NOT (fsm_output(7))) OR (fsm_output(2)) OR (NOT
      (fsm_output(3))) OR (fsm_output(8)) OR (NOT (fsm_output(9)));
  mux_2062_nl <= MUX_s_1_2_2(or_1995_cse, nand_357_cse, fsm_output(0));
  mux_2063_nl <= MUX_s_1_2_2(or_2218_nl, mux_2062_nl, fsm_output(4));
  mux_2064_nl <= MUX_s_1_2_2(or_2219_nl, mux_2063_nl, fsm_output(5));
  or_2214_nl <= (fsm_output(4)) OR (NOT (fsm_output(0))) OR (fsm_output(7)) OR (NOT
      (fsm_output(2))) OR (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(9));
  mux_2061_nl <= MUX_s_1_2_2(or_2214_nl, mux_tmp_2006, fsm_output(5));
  mux_2065_nl <= MUX_s_1_2_2(mux_2064_nl, mux_2061_nl, fsm_output(6));
  or_2209_nl <= (fsm_output(4)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(7)))
      OR (fsm_output(2)) OR (fsm_output(3)) OR (fsm_output(8)) OR (fsm_output(9));
  mux_2059_nl <= MUX_s_1_2_2(mux_tmp_2006, or_2209_nl, fsm_output(5));
  or_2207_nl <= (fsm_output(0)) OR (fsm_output(7)) OR (fsm_output(2)) OR (NOT (fsm_output(3)))
      OR (fsm_output(8)) OR (NOT (fsm_output(9)));
  mux_2055_nl <= MUX_s_1_2_2(or_1976_cse, mux_1768_cse, fsm_output(0));
  mux_2056_nl <= MUX_s_1_2_2(or_2207_nl, mux_2055_nl, fsm_output(4));
  or_2208_nl <= (fsm_output(5)) OR mux_2056_nl;
  mux_2060_nl <= MUX_s_1_2_2(mux_2059_nl, or_2208_nl, fsm_output(6));
  mux_2066_cse <= MUX_s_1_2_2(mux_2065_nl, mux_2060_nl, fsm_output(1));
  and_dcpl_231 <= NOT((fsm_output(1)) OR (fsm_output(6)));
  and_dcpl_232 <= and_dcpl_231 AND (NOT (fsm_output(5)));
  and_dcpl_233 <= and_dcpl_232 AND and_dcpl_29;
  and_dcpl_234 <= (NOT (fsm_output(7))) AND (fsm_output(2));
  and_dcpl_236 <= NOT((fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(3)));
  and_dcpl_237 <= and_dcpl_236 AND and_dcpl_234;
  and_dcpl_238 <= and_dcpl_237 AND and_dcpl_233;
  and_dcpl_242 <= and_dcpl_237 AND and_dcpl_231 AND (fsm_output(5)) AND and_dcpl_32;
  and_dcpl_243 <= (NOT (fsm_output(1))) AND (fsm_output(6));
  and_dcpl_244 <= and_dcpl_243 AND (NOT (fsm_output(5)));
  and_dcpl_246 <= and_dcpl_237 AND and_dcpl_244 AND and_dcpl_29;
  and_dcpl_248 <= (fsm_output(1)) AND (NOT (fsm_output(6))) AND (fsm_output(5));
  and_dcpl_250 <= (fsm_output(7)) AND (NOT (fsm_output(2)));
  and_dcpl_251 <= and_dcpl_236 AND and_dcpl_250;
  and_dcpl_252 <= and_dcpl_251 AND and_dcpl_248 AND and_dcpl_29;
  and_dcpl_255 <= and_dcpl_251 AND and_dcpl_243 AND (fsm_output(5)) AND and_dcpl_32;
  and_dcpl_256 <= NOT((fsm_output(7)) OR (fsm_output(2)));
  and_dcpl_260 <= and_dcpl_70 AND (NOT (fsm_output(3))) AND and_dcpl_256 AND and_dcpl_233;
  and_dcpl_265 <= and_dcpl_70 AND (fsm_output(3));
  and_dcpl_267 <= and_dcpl_265 AND and_dcpl_234 AND (fsm_output(1)) AND (fsm_output(6))
      AND (fsm_output(5)) AND and_dcpl_16;
  and_dcpl_271 <= and_dcpl_265 AND (fsm_output(7)) AND (fsm_output(2));
  and_dcpl_272 <= and_dcpl_271 AND and_dcpl_232 AND and_dcpl_66;
  and_dcpl_274 <= and_dcpl_271 AND and_dcpl_244 AND and_dcpl_16;
  and_dcpl_277 <= (fsm_output(9)) AND (NOT (fsm_output(8))) AND (fsm_output(3));
  and_dcpl_278 <= and_dcpl_277 AND and_dcpl_256;
  and_dcpl_279 <= and_dcpl_278 AND and_dcpl_248 AND and_dcpl_16;
  and_dcpl_281 <= and_dcpl_278 AND and_dcpl_244 AND and_dcpl_66;
  and_dcpl_284 <= and_dcpl_277 AND and_dcpl_250 AND and_dcpl_232 AND and_dcpl_16;
  and_dcpl_293 <= and_dcpl_236 AND (NOT (fsm_output(7))) AND (fsm_output(2)) AND
      (NOT (fsm_output(1))) AND (NOT (fsm_output(6))) AND (NOT (fsm_output(5))) AND
      (NOT (fsm_output(0))) AND (fsm_output(4));
  and_dcpl_300 <= and_dcpl_236 AND and_dcpl_250 AND (fsm_output(1)) AND (NOT (fsm_output(6)))
      AND (NOT (fsm_output(5))) AND (fsm_output(0)) AND (NOT (fsm_output(4)));
  and_dcpl_308 <= (fsm_output(8)) AND (NOT (fsm_output(9))) AND (fsm_output(3)) AND
      and_dcpl_250 AND (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(5)) AND
      (fsm_output(0)) AND (fsm_output(4));
  and_dcpl_344 <= NOT(CONV_SL_1_1(fsm_output/=STD_LOGIC_VECTOR'("0000010100")));
  and_dcpl_361 <= (NOT (fsm_output(9))) AND (fsm_output(8)) AND (fsm_output(3)) AND
      and_dcpl_234 AND (fsm_output(1)) AND (NOT (fsm_output(6))) AND (fsm_output(5))
      AND (fsm_output(0)) AND (fsm_output(4));
  and_dcpl_376 <= (fsm_output(1)) AND (NOT (fsm_output(6)));
  and_dcpl_382 <= and_dcpl_376 AND (fsm_output(5));
  and_dcpl_396 <= and_dcpl_382 AND and_dcpl_66;
  and_dcpl_398 <= and_dcpl_265 AND and_dcpl_234;
  and_dcpl_402 <= (fsm_output(1)) AND (fsm_output(6)) AND (fsm_output(5));
  and_dcpl_403 <= and_dcpl_402 AND and_dcpl_16;
  and_dcpl_406 <= (fsm_output(7)) AND (fsm_output(2));
  and_dcpl_407 <= and_dcpl_265 AND and_dcpl_406;
  and_dcpl_416 <= and_dcpl_98 AND (fsm_output(3));
  and_dcpl_417 <= and_dcpl_416 AND and_dcpl_256;
  and_dcpl_425 <= and_dcpl_98 AND (NOT (fsm_output(3))) AND and_dcpl_406;
  and_dcpl_444 <= NOT((fsm_output(9)) OR (fsm_output(8)) OR (fsm_output(3)) OR (NOT
      and_dcpl_234) OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(5)) OR (NOT
      (fsm_output(0))) OR (fsm_output(4)));
  and_dcpl_460 <= (fsm_output(8)) AND (fsm_output(9)) AND (NOT (fsm_output(3))) AND
      (NOT (fsm_output(7))) AND (fsm_output(2)) AND (fsm_output(1)) AND (NOT (fsm_output(6)))
      AND (NOT (fsm_output(5))) AND and_dcpl_16;
  nor_761_cse <= NOT((fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(5)));
  and_dcpl_464 <= nor_761_cse AND (fsm_output(0)) AND (NOT (fsm_output(4)));
  and_551_ssc <= (fsm_output(9)) AND (NOT (fsm_output(8))) AND (NOT (fsm_output(3)))
      AND (fsm_output(7)) AND (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(6))
      AND (fsm_output(5)) AND and_dcpl_16;
  nand_tmp_139 <= NOT((fsm_output(3)) AND (NOT(and_dcpl_16 OR CONV_SL_1_1(fsm_output(9
      DOWNTO 8)/=STD_LOGIC_VECTOR'("01")))));
  or_tmp_2154 <= (fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(8)) OR (fsm_output(9));
  or_2261_nl <= (NOT (fsm_output(3))) OR (fsm_output(4)) OR (fsm_output(0)) OR (NOT
      (fsm_output(8))) OR (fsm_output(9));
  mux_tmp_2041 <= MUX_s_1_2_2(or_tmp_2154, or_2261_nl, fsm_output(2));
  or_tmp_2156 <= nor_810_cse OR CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"));
  or_2267_nl <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(8)) OR (fsm_output(9));
  or_2266_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(8))) OR (fsm_output(9));
  mux_tmp_2043 <= MUX_s_1_2_2(or_2267_nl, or_2266_nl, fsm_output(3));
  or_2271_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(0))) OR (fsm_output(8))
      OR (fsm_output(9));
  or_2270_nl <= (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(8)) OR (NOT (fsm_output(9)));
  mux_2097_nl <= MUX_s_1_2_2(or_2271_nl, or_2270_nl, fsm_output(3));
  nand_388_nl <= NOT((fsm_output(3)) AND (NOT(nor_810_cse OR CONV_SL_1_1(fsm_output(9
      DOWNTO 8)/=STD_LOGIC_VECTOR'("01")))));
  mux_tmp_2046 <= MUX_s_1_2_2(mux_2097_nl, nand_388_nl, fsm_output(2));
  or_tmp_2166 <= (NOT (fsm_output(0))) OR (fsm_output(8)) OR (NOT (fsm_output(9)));
  or_tmp_2168 <= (fsm_output(3)) OR and_dcpl_66 OR CONV_SL_1_1(fsm_output(9 DOWNTO
      8)/=STD_LOGIC_VECTOR'("00"));
  nand_389_nl <= NOT((fsm_output(3)) AND (NOT or_tmp_2156));
  mux_2103_nl <= MUX_s_1_2_2(nand_389_nl, mux_tmp_2043, fsm_output(2));
  or_2272_nl <= (fsm_output(4)) OR (fsm_output(0)) OR (NOT (fsm_output(8))) OR (fsm_output(9));
  mux_2101_nl <= MUX_s_1_2_2(or_tmp_2166, or_2272_nl, fsm_output(3));
  mux_2102_nl <= MUX_s_1_2_2(or_tmp_2168, mux_2101_nl, fsm_output(2));
  mux_tmp_2052 <= MUX_s_1_2_2(mux_2103_nl, mux_2102_nl, fsm_output(7));
  or_tmp_2171 <= and_dcpl_16 OR CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("10"));
  or_2282_nl <= (NOT (fsm_output(3))) OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(8))
      OR (NOT (fsm_output(9)));
  mux_tmp_2058 <= MUX_s_1_2_2(or_2282_nl, nand_tmp_139, fsm_output(2));
  or_tmp_2183 <= NOT((fsm_output(4)) AND (fsm_output(7)) AND (fsm_output(8)) AND
      (fsm_output(3)) AND (NOT (fsm_output(9))));
  mux_2123_nl <= MUX_s_1_2_2(mux_tmp_1610, or_tmp_1796, fsm_output(4));
  mux_tmp_2072 <= MUX_s_1_2_2(or_tmp_2183, mux_2123_nl, fsm_output(0));
  not_tmp_571 <= NOT((fsm_output(3)) AND (fsm_output(9)));
  or_tmp_2191 <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00")) OR
      not_tmp_571;
  or_tmp_2193 <= (NOT (fsm_output(4))) OR (fsm_output(7)) OR (fsm_output(8)) OR not_tmp_571;
  or_2302_nl <= (fsm_output(8)) OR not_tmp_571;
  mux_tmp_2081 <= MUX_s_1_2_2(or_2302_nl, or_2012_cse, fsm_output(7));
  mux_2134_nl <= MUX_s_1_2_2(mux_tmp_2081, or_tmp_2193, fsm_output(0));
  mux_2131_nl <= MUX_s_1_2_2(or_tmp_1793, or_tmp_1796, fsm_output(4));
  mux_2132_nl <= MUX_s_1_2_2(mux_2131_nl, mux_1583_cse, fsm_output(0));
  mux_tmp_2083 <= MUX_s_1_2_2(mux_2134_nl, mux_2132_nl, fsm_output(2));
  mux_tmp_2108 <= MUX_s_1_2_2(mux_tmp_1874, mux_tmp_1861, fsm_output(1));
  or_tmp_2223 <= (CONV_SL_1_1(fsm_output(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"))) OR
      CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"));
  mux_2163_nl <= MUX_s_1_2_2(or_tmp_2041, mux_1920_cse, fsm_output(1));
  mux_tmp_2112 <= MUX_s_1_2_2(or_tmp_2223, mux_2163_nl, fsm_output(7));
  or_tmp_2227 <= (NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000"))))
      OR CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"));
  mux_2169_nl <= MUX_s_1_2_2(or_tmp_2041, mux_1922_cse, fsm_output(1));
  mux_2170_nl <= MUX_s_1_2_2(or_tmp_2227, mux_2169_nl, fsm_output(7));
  mux_2166_nl <= MUX_s_1_2_2(nand_tmp_134, mux_tmp_1861, fsm_output(1));
  mux_2167_nl <= MUX_s_1_2_2(mux_2166_nl, or_tmp_2037, fsm_output(7));
  mux_tmp_2119 <= MUX_s_1_2_2(mux_2170_nl, mux_2167_nl, fsm_output(6));
  mux_2175_nl <= MUX_s_1_2_2(nand_tmp_134, mux_tmp_1874, fsm_output(1));
  mux_tmp_2124 <= MUX_s_1_2_2(mux_2175_nl, or_tmp_2037, fsm_output(7));
  mux_2179_nl <= MUX_s_1_2_2(mux_1938_cse, or_tmp_2041, fsm_output(1));
  mux_tmp_2128 <= MUX_s_1_2_2(mux_2179_nl, mux_tmp_1861, fsm_output(7));
  or_tmp_2236 <= CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_2150 <= MUX_s_1_2_2(or_tmp_2236, (fsm_output(8)), or_2146_cse);
  mux_tmp_2153 <= MUX_s_1_2_2((fsm_output(8)), or_2086_cse, fsm_output(2));
  mux_tmp_2154 <= MUX_s_1_2_2(mux_tmp_2153, or_tmp_2043, fsm_output(3));
  mux_tmp_2156 <= MUX_s_1_2_2(or_tmp_2236, (fsm_output(8)), fsm_output(3));
  mux_tmp_2159 <= MUX_s_1_2_2(mux_tmp_2154, or_tmp_2037, fsm_output(4));
  or_2346_nl <= and_357_cse OR CONV_SL_1_1(fsm_output(9 DOWNTO 8)/=STD_LOGIC_VECTOR'("01"));
  mux_2215_nl <= MUX_s_1_2_2(mux_tmp_1861, mux_tmp_2156, fsm_output(0));
  mux_tmp_2164 <= MUX_s_1_2_2(or_2346_nl, mux_2215_nl, fsm_output(4));
  mux_tmp_2165 <= MUX_s_1_2_2(mux_tmp_1861, mux_tmp_2154, fsm_output(4));
  mux_tmp_2167 <= MUX_s_1_2_2(mux_tmp_2153, or_tmp_2044, fsm_output(3));
  mux_2220_nl <= MUX_s_1_2_2(mux_tmp_2167, mux_tmp_2154, fsm_output(0));
  mux_tmp_2169 <= MUX_s_1_2_2(mux_2220_nl, or_212_cse, fsm_output(4));
  mux_tmp_2170 <= MUX_s_1_2_2(or_212_cse, mux_tmp_1861, fsm_output(4));
  mux_tmp_2179 <= MUX_s_1_2_2(or_tmp_2236, (fsm_output(8)), fsm_output(2));
  mux_tmp_2180 <= MUX_s_1_2_2(or_tmp_2035, mux_tmp_2179, fsm_output(3));
  or_tmp_2243 <= (fsm_output(5)) OR (fsm_output(1));
  or_tmp_2244 <= (fsm_output(5)) OR (NOT (fsm_output(1)));
  mux_tmp_2192 <= MUX_s_1_2_2(or_tmp_2244, or_tmp_2243, fsm_output(0));
  or_2350_nl <= (NOT((fsm_output(0)) OR (fsm_output(5)))) OR (fsm_output(1));
  mux_tmp_2193 <= MUX_s_1_2_2(mux_tmp_2192, or_2350_nl, fsm_output(4));
  or_tmp_2245 <= (fsm_output(0)) OR (NOT((fsm_output(5)) AND (fsm_output(1))));
  mux_tmp_2196 <= MUX_s_1_2_2(or_tmp_2245, or_tmp_2244, fsm_output(4));
  nand_399_nl <= NOT((fsm_output(0)) AND (fsm_output(5)) AND (fsm_output(1)));
  mux_2249_itm <= MUX_s_1_2_2(nand_399_nl, mux_tmp_2196, fsm_output(6));
  mux_tmp_2199 <= MUX_s_1_2_2(or_tmp_2243, or_2186_cse, fsm_output(4));
  or_2360_nl <= (NOT (fsm_output(0))) OR (NOT (fsm_output(5))) OR (fsm_output(1));
  mux_tmp_2204 <= MUX_s_1_2_2(or_2360_nl, mux_tmp_2192, fsm_output(4));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((and_dcpl_19 AND and_dcpl_15) OR STAGE_LOOP_i_3_0_sva_mx0c1) = '1' )
          THEN
        STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(STD_LOGIC_VECTOR'( "0001"), (z_out_7(3
            DOWNTO 0)), STAGE_LOOP_i_3_0_sva_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_121 = '0' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( not_tmp_121 = '0' ) THEN
        r_sva <= r_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        COMP_LOOP_nor_11_itm <= '0';
        COMP_LOOP_COMP_LOOP_nor_1_itm <= '0';
        COMP_LOOP_nor_12_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_139_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_140_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_141_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_143_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_144_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_145_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_146_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_147_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_148_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_149_itm <= '0';
        COMP_LOOP_nor_134_itm <= '0';
        COMP_LOOP_nor_137_itm <= '0';
      ELSE
        reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_18 AND and_dcpl_16 AND (fsm_output(1))
            AND (fsm_output(2)) AND (NOT (fsm_output(6))) AND (fsm_output(9)) AND
            (fsm_output(8)) AND (NOT (z_out_8_64_2(0)));
        reg_ensig_cgo_cse <= NOT mux_1581_itm;
        COMP_LOOP_nor_11_itm <= MUX_s_1_2_2((z_out_3(5)), COMP_LOOP_nor_11_nl, modExp_dev_while_or_2_cse);
        COMP_LOOP_COMP_LOOP_nor_1_itm <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_nor_12_itm <= NOT((z_out_6_10_1(3)) OR (z_out_6_10_1(2)) OR (z_out_6_10_1(0)));
        COMP_LOOP_COMP_LOOP_and_139_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_140_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_141_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_COMP_LOOP_and_143_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_144_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_145_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
        COMP_LOOP_COMP_LOOP_and_146_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_147_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_148_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_149_itm <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"));
        COMP_LOOP_nor_134_itm <= NOT((z_out_6_10_1(3)) OR (z_out_6_10_1(1)) OR (z_out_6_10_1(0)));
        COMP_LOOP_nor_137_itm <= NOT(CONV_SL_1_1(z_out_6_10_1(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_9, (operator_64_false_acc_mut_64
          & operator_64_false_acc_mut_63_0), and_dcpl_169);
      operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
          STAGE_LOOP_lshift_psp_sva, and_dcpl_169);
      modExp_dev_exp_1_sva_3_0 <= MUX_v_4_2_2(COMP_LOOP_and_nl, STD_LOGIC_VECTOR'("1111"),
          and_dcpl_221);
      COMP_LOOP_1_mul_itm <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED'( SIGNED(operator_64_false_acc_mut_63_0)
          * SIGNED(COMP_LOOP_mux1h_209_nl)), 64));
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(nor_271_nl, and_tmp_12, fsm_output(8))) = '1' ) THEN
        STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_2121_nl = '0' ) THEN
        operator_64_false_acc_mut_64 <= operator_64_false_operator_64_false_mux_rgt(64);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mux_2153_nl = '0' ) THEN
        operator_64_false_acc_mut_63_0 <= operator_64_false_operator_64_false_mux_rgt(63
            DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        VEC_LOOP_j_sva_9_0 <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( ((NOT(mux_tmp_1688 OR (fsm_output(5)) OR (fsm_output(7)) OR (fsm_output(3))
          OR (fsm_output(6)) OR (NOT nor_697_cse))) OR VEC_LOOP_j_sva_9_0_mx0c1)
          = '1' ) THEN
        VEC_LOOP_j_sva_9_0 <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"), (VEC_LOOP_acc_1_psp_1(9
            DOWNTO 0)), VEC_LOOP_j_sva_9_0_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(mux_2156_nl OR (fsm_output(3)))) = '1' ) THEN
        COMP_LOOP_k_9_4_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (z_out_3(4
            DOWNTO 0)), or_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_1749_nl OR and_195_rgt) = '1' ) THEN
        modExp_dev_result_sva <= MUX_v_64_2_2(STD_LOGIC_VECTOR'( "0000000000000000000000000000000000000000000000000000000000000001"),
            modulo_dev_cmp_return_rsc_z, and_195_rgt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_1754_nl OR CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("000"))
          OR (NOT nor_697_cse)) = '1' ) THEN
        modExp_dev_exp_sva <= MUX_v_64_2_2((operator_66_true_div_cmp_z(63 DOWNTO
            0)), (z_out_9(63 DOWNTO 0)), and_dcpl_183);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= '0';
      ELSIF ( (and_dcpl_183 OR not_tmp_402 OR and_dcpl_36 OR and_dcpl_44 OR and_dcpl_52
          OR and_dcpl_58 OR and_dcpl_63 OR and_dcpl_72 OR and_dcpl_78 OR and_dcpl_84
          OR and_dcpl_90 OR and_dcpl_93 OR and_dcpl_97 OR and_dcpl_102 OR and_dcpl_106
          OR and_dcpl_110 OR and_dcpl_115 OR and_dcpl_119) = '1' ) THEN
        COMP_LOOP_COMP_LOOP_and_137_itm <= MUX_s_1_2_2((NOT (z_out_7(64))), COMP_LOOP_COMP_LOOP_and_17_nl,
            modExp_dev_while_or_2_cse);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(or_tmp_74 OR (fsm_output(3)) OR (NOT (fsm_output(4))) OR (fsm_output(0))
          OR (fsm_output(1)) OR (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(9))
          OR (fsm_output(8)))) = '1' ) THEN
        COMP_LOOP_acc_psp_sva <= z_out_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_244_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_62_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_2_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_64_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_4_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_5_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_6_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_68_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_8_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_9_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_11_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_12_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_13_itm <= '0';
        COMP_LOOP_COMP_LOOP_and_14_itm <= '0';
      ELSIF ( mux_1832_itm = '1' ) THEN
        COMP_LOOP_COMP_LOOP_nor_itm <= NOT(CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)/=STD_LOGIC_VECTOR'("0000")));
        COMP_LOOP_COMP_LOOP_and_244_itm <= (COMP_LOOP_acc_13_psp_sva_1(0)) AND (VEC_LOOP_j_sva_9_0(0))
            AND (NOT((COMP_LOOP_acc_13_psp_sva_1(1)) OR (VEC_LOOP_j_sva_9_0(1))));
        COMP_LOOP_COMP_LOOP_and_62_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_COMP_LOOP_and_2_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0011"));
        COMP_LOOP_COMP_LOOP_and_64_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_4_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0101"));
        COMP_LOOP_COMP_LOOP_and_5_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0110"));
        COMP_LOOP_COMP_LOOP_and_6_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("0111"));
        COMP_LOOP_COMP_LOOP_and_68_itm <= CONV_SL_1_1(COMP_LOOP_acc_1_cse_2_sva_1(3
            DOWNTO 0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_8_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1001"));
        COMP_LOOP_COMP_LOOP_and_9_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1010"));
        COMP_LOOP_COMP_LOOP_and_11_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1100"));
        COMP_LOOP_COMP_LOOP_and_12_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1101"));
        COMP_LOOP_COMP_LOOP_and_13_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1110"));
        COMP_LOOP_COMP_LOOP_and_14_itm <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO
            0)=STD_LOGIC_VECTOR'("1111"));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_COMP_LOOP_and_10_itm <= '0';
      ELSIF ( mux_1842_nl = '0' ) THEN
        COMP_LOOP_COMP_LOOP_and_10_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_10_nl,
            (NOT (COMP_LOOP_1_acc_nl(9))), and_dcpl_119);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_13_psp_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (NOT(mux_1845_nl AND nor_697_cse)) = '1' ) THEN
        COMP_LOOP_acc_13_psp_sva <= COMP_LOOP_acc_13_psp_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_2_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( ((NOT mux_1848_nl) OR CONV_SL_1_1(fsm_output(9 DOWNTO 7)/=STD_LOGIC_VECTOR'("000")))
          = '1' ) THEN
        COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (NOT((NOT mux_1858_nl) AND nor_697_cse)) = '1' ) THEN
        COMP_LOOP_acc_11_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0(9
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "001")), 8), 9), 9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_4_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (NOT(mux_1862_nl AND nor_697_cse)) = '1' ) THEN
        COMP_LOOP_acc_1_cse_4_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "0011")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_6_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_1866_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_6_sva <= z_out_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (mux_1869_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_14_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0(9
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "011")), 8), 9), 9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_8_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_1872_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_8_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "0111")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_16_psp_sva <= STD_LOGIC_VECTOR'( "0000000");
      ELSIF ( (mux_1874_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_16_psp_sva <= z_out_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_10_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (mux_1875_nl OR (fsm_output(9))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_10_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1001")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_17_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (MUX_s_1_2_2(mux_1877_nl, (fsm_output(9)), fsm_output(8))) = '1' )
          THEN
        COMP_LOOP_acc_17_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0(9
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "101")), 8), 9), 9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_12_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_1880_nl, (fsm_output(9)), fsm_output(8))) = '1' )
          THEN
        COMP_LOOP_acc_1_cse_12_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1011")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_19_psp_sva <= STD_LOGIC_VECTOR'( "00000000");
      ELSIF ( (MUX_s_1_2_2(mux_1885_nl, (fsm_output(9)), or_110_nl)) = '1' ) THEN
        COMP_LOOP_acc_19_psp_sva <= z_out_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_14_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(mux_1888_nl, (fsm_output(9)), fsm_output(8))) = '1' )
          THEN
        COMP_LOOP_acc_1_cse_14_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1101")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_20_psp_sva <= STD_LOGIC_VECTOR'( "000000000");
      ELSIF ( (MUX_s_1_2_2(mux_1896_nl, (fsm_output(9)), fsm_output(8))) = '1' )
          THEN
        COMP_LOOP_acc_20_psp_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0(9
            DOWNTO 1)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
            & STD_LOGIC_VECTOR'( "111")), 8), 9), 9));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR'( "0000000000");
      ELSIF ( (MUX_s_1_2_2(nor_nl, and_nl, fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_1_cse_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0)
            + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & STD_LOGIC_VECTOR'(
            "1111")), 9), 10), 10));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_199 OR and_dcpl_200 OR and_dcpl_201 OR and_dcpl_202 OR and_dcpl_203
          OR and_dcpl_204 OR and_dcpl_206 OR and_dcpl_208 OR and_dcpl_210 OR and_dcpl_212
          OR and_dcpl_214 OR and_dcpl_215 OR and_dcpl_217 OR and_dcpl_219 OR and_dcpl_220
          OR and_dcpl_221) = '1' ) THEN
        tmp_10_lpi_4_dfm <= MUX1HOT_v_64_16_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
            vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
            vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
            vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
            vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_or_6_nl
            & COMP_LOOP_or_7_nl & COMP_LOOP_or_8_nl & COMP_LOOP_or_9_nl & COMP_LOOP_or_10_nl
            & COMP_LOOP_or_11_nl & COMP_LOOP_or_12_nl & COMP_LOOP_or_13_nl & COMP_LOOP_or_14_nl
            & COMP_LOOP_or_15_nl & COMP_LOOP_or_16_nl & COMP_LOOP_or_17_nl & COMP_LOOP_or_18_nl
            & COMP_LOOP_or_19_nl & COMP_LOOP_or_20_nl & COMP_LOOP_or_21_nl));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (MUX_s_1_2_2(mux_2196_nl, mux_2184_nl, fsm_output(4))) = '1' ) THEN
        modExp_dev_exp_1_sva_63_9 <= MUX_v_55_2_2(STD_LOGIC_VECTOR'("0000000000000000000000000000000000000000000000000000000"),
            (z_out_9(63 DOWNTO 9)), not_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva_9_5 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( mux_2243_nl = '0' ) THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva_9_5 <= COMP_LOOP_mux1h_192_rgt(9 DOWNTO 5);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
      ELSIF ( (MUX_s_1_2_2(mux_2262_nl, nor_800_nl, fsm_output(8))) = '1' ) THEN
        COMP_LOOP_acc_10_cse_10_1_1_sva_4_0 <= COMP_LOOP_mux1h_192_rgt(4 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_36 OR and_dcpl_44 OR and_dcpl_58 OR and_dcpl_63 OR and_dcpl_72
          OR and_dcpl_84 OR and_dcpl_90 OR and_dcpl_93 OR and_dcpl_102 OR and_dcpl_106
          OR and_dcpl_110) = '1' ) THEN
        COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm <= z_out_1(9);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (and_dcpl_52 OR and_dcpl_78 OR and_dcpl_97 OR and_dcpl_115) = '1' ) THEN
        COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= MUX1HOT_s_1_3_2((z_out_2(7)), (z_out_5(6)),
            (z_out_4(5)), STD_LOGIC_VECTOR'( COMP_LOOP_or_27_nl & and_dcpl_78 & and_dcpl_115));
      END IF;
    END IF;
  END PROCESS;
  COMP_LOOP_nor_11_nl <= NOT(CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  mux_1950_nl <= MUX_s_1_2_2(mux_1949_cse, mux_tmp_1874, fsm_output(7));
  mux_1951_nl <= MUX_s_1_2_2(mux_1950_nl, mux_tmp_1888, fsm_output(0));
  mux_1952_nl <= MUX_s_1_2_2(mux_tmp_1891, mux_1951_nl, fsm_output(5));
  mux_1948_nl <= MUX_s_1_2_2(mux_tmp_1876, mux_tmp_1883, fsm_output(5));
  mux_1953_nl <= MUX_s_1_2_2(mux_1952_nl, mux_1948_nl, fsm_output(6));
  mux_1944_nl <= MUX_s_1_2_2(nand_tmp_134, or_212_cse, fsm_output(7));
  mux_1945_nl <= MUX_s_1_2_2(mux_1944_nl, mux_tmp_1876, fsm_output(0));
  mux_1943_nl <= MUX_s_1_2_2(mux_tmp_1891, mux_tmp_1882, fsm_output(0));
  mux_1946_nl <= MUX_s_1_2_2(mux_1945_nl, mux_1943_nl, fsm_output(5));
  mux_1940_nl <= MUX_s_1_2_2(mux_tmp_1888, mux_tmp_1866, fsm_output(0));
  mux_1941_nl <= MUX_s_1_2_2(mux_1940_nl, mux_tmp_1877, fsm_output(5));
  mux_1947_nl <= MUX_s_1_2_2(mux_1946_nl, mux_1941_nl, fsm_output(6));
  mux_1954_nl <= MUX_s_1_2_2(mux_1953_nl, mux_1947_nl, fsm_output(4));
  mux_1935_nl <= MUX_s_1_2_2(mux_tmp_1883, mux_tmp_1866, fsm_output(5));
  mux_1931_nl <= MUX_s_1_2_2(mux_tmp_1875, mux_tmp_1863, fsm_output(0));
  mux_1932_nl <= MUX_s_1_2_2(mux_1931_nl, mux_tmp_1870, fsm_output(5));
  mux_1936_nl <= MUX_s_1_2_2(mux_1935_nl, mux_1932_nl, fsm_output(6));
  mux_1924_nl <= MUX_s_1_2_2(mux_tmp_1872, mux_tmp_1870, fsm_output(0));
  mux_1929_nl <= MUX_s_1_2_2(mux_tmp_1877, mux_1924_nl, fsm_output(5));
  mux_1916_nl <= MUX_s_1_2_2(or_tmp_2041, or_2336_cse, fsm_output(7));
  mux_1918_nl <= MUX_s_1_2_2(mux_tmp_1866, mux_1916_nl, fsm_output(0));
  mux_1913_nl <= MUX_s_1_2_2(mux_tmp_1861, or_1916_cse, fsm_output(7));
  mux_1915_nl <= MUX_s_1_2_2(mux_tmp_1863, mux_1913_nl, fsm_output(0));
  mux_1919_nl <= MUX_s_1_2_2(mux_1918_nl, mux_1915_nl, fsm_output(5));
  mux_1930_nl <= MUX_s_1_2_2(mux_1929_nl, mux_1919_nl, fsm_output(6));
  mux_1937_nl <= MUX_s_1_2_2(mux_1936_nl, mux_1930_nl, fsm_output(4));
  mux_1955_nl <= MUX_s_1_2_2(mux_1954_nl, mux_1937_nl, fsm_output(1));
  COMP_LOOP_mux1h_186_nl <= MUX1HOT_v_4_16_2((z_out_9(3 DOWNTO 0)), modExp_dev_exp_1_sva_3_0,
      STD_LOGIC_VECTOR'( "0001"), STD_LOGIC_VECTOR'( "0010"), STD_LOGIC_VECTOR'(
      "0011"), STD_LOGIC_VECTOR'( "0100"), STD_LOGIC_VECTOR'( "0101"), STD_LOGIC_VECTOR'(
      "0110"), STD_LOGIC_VECTOR'( "0111"), STD_LOGIC_VECTOR'( "1000"), STD_LOGIC_VECTOR'(
      "1001"), STD_LOGIC_VECTOR'( "1010"), STD_LOGIC_VECTOR'( "1011"), STD_LOGIC_VECTOR'(
      "1100"), STD_LOGIC_VECTOR'( "1101"), STD_LOGIC_VECTOR'( "1110"), STD_LOGIC_VECTOR'(
      not_tmp_402 & (NOT mux_1955_nl) & and_dcpl_200 & and_dcpl_201 & and_dcpl_202
      & and_dcpl_203 & and_dcpl_204 & and_dcpl_206 & and_dcpl_208 & and_dcpl_210
      & and_dcpl_212 & and_dcpl_214 & and_dcpl_215 & and_dcpl_217 & and_dcpl_219
      & and_dcpl_220));
  not_4628_nl <= NOT and_dcpl_199;
  COMP_LOOP_and_nl <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), COMP_LOOP_mux1h_186_nl,
      not_4628_nl);
  COMP_LOOP_COMP_LOOP_and_930_nl <= (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(0)) AND
      COMP_LOOP_nor_11_itm;
  COMP_LOOP_COMP_LOOP_and_932_nl <= (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(1)) AND
      COMP_LOOP_nor_12_itm;
  COMP_LOOP_COMP_LOOP_and_934_nl <= (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(2)) AND
      COMP_LOOP_nor_134_itm;
  COMP_LOOP_COMP_LOOP_and_936_nl <= (COMP_LOOP_acc_10_cse_10_1_1_sva_4_0(3)) AND
      COMP_LOOP_nor_137_itm;
  COMP_LOOP_mux1h_209_nl <= MUX1HOT_v_64_16_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
      vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
      vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
      vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
      vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, STD_LOGIC_VECTOR'( COMP_LOOP_COMP_LOOP_nor_1_itm
      & COMP_LOOP_COMP_LOOP_and_930_nl & COMP_LOOP_COMP_LOOP_and_932_nl & COMP_LOOP_COMP_LOOP_and_137_itm
      & COMP_LOOP_COMP_LOOP_and_934_nl & COMP_LOOP_COMP_LOOP_and_139_itm & COMP_LOOP_COMP_LOOP_and_140_itm
      & COMP_LOOP_COMP_LOOP_and_141_itm & COMP_LOOP_COMP_LOOP_and_936_nl & COMP_LOOP_COMP_LOOP_and_143_itm
      & COMP_LOOP_COMP_LOOP_and_144_itm & COMP_LOOP_COMP_LOOP_and_145_itm & COMP_LOOP_COMP_LOOP_and_146_itm
      & COMP_LOOP_COMP_LOOP_and_147_itm & COMP_LOOP_COMP_LOOP_and_148_itm & COMP_LOOP_COMP_LOOP_and_149_itm));
  nor_271_nl <= NOT((fsm_output(9)) OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(1))
      OR (fsm_output(4)) OR (fsm_output(3)) OR (fsm_output(7)) OR (fsm_output(5)));
  or_2286_nl <= (NOT((fsm_output(0)) OR (fsm_output(8)))) OR (fsm_output(9));
  or_2284_nl <= (fsm_output(0)) OR (NOT (fsm_output(8))) OR (fsm_output(9));
  mux_2116_nl <= MUX_s_1_2_2(or_2286_nl, or_2284_nl, fsm_output(4));
  or_2287_nl <= (fsm_output(3)) OR mux_2116_nl;
  mux_2117_nl <= MUX_s_1_2_2(or_2287_nl, or_tmp_2154, fsm_output(2));
  mux_2118_nl <= MUX_s_1_2_2(mux_2117_nl, mux_tmp_2058, fsm_output(7));
  or_2283_nl <= (NOT (fsm_output(4))) OR (fsm_output(0)) OR (NOT (fsm_output(8)))
      OR (fsm_output(9));
  mux_2113_nl <= MUX_s_1_2_2(or_2283_nl, or_tmp_2166, fsm_output(3));
  mux_2114_nl <= MUX_s_1_2_2(mux_2113_nl, or_tmp_2168, fsm_output(2));
  mux_2115_nl <= MUX_s_1_2_2(mux_2114_nl, mux_tmp_2046, fsm_output(7));
  mux_2119_nl <= MUX_s_1_2_2(mux_2118_nl, mux_2115_nl, fsm_output(5));
  or_2280_nl <= (fsm_output(3)) OR or_tmp_2171;
  mux_2109_nl <= MUX_s_1_2_2(or_tmp_2168, or_2280_nl, fsm_output(2));
  mux_2111_nl <= MUX_s_1_2_2(mux_tmp_2058, mux_2109_nl, fsm_output(7));
  mux_2112_nl <= MUX_s_1_2_2(mux_tmp_2052, mux_2111_nl, fsm_output(5));
  mux_2120_nl <= MUX_s_1_2_2(mux_2119_nl, mux_2112_nl, fsm_output(1));
  nand_390_nl <= NOT((fsm_output(3)) AND (NOT or_tmp_2171));
  mux_2105_nl <= MUX_s_1_2_2(nand_390_nl, or_tmp_2168, fsm_output(2));
  mux_2106_nl <= MUX_s_1_2_2(mux_2105_nl, mux_tmp_2041, fsm_output(7));
  mux_2107_nl <= MUX_s_1_2_2(mux_2106_nl, mux_tmp_2052, fsm_output(5));
  or_2265_nl <= (fsm_output(3)) OR or_tmp_2156;
  mux_2096_nl <= MUX_s_1_2_2(mux_tmp_2043, or_2265_nl, fsm_output(2));
  mux_2099_nl <= MUX_s_1_2_2(mux_tmp_2046, mux_2096_nl, fsm_output(7));
  or_2258_nl <= (fsm_output(3)) OR (fsm_output(4)) OR (fsm_output(0)) OR (fsm_output(8))
      OR (NOT (fsm_output(9)));
  mux_nl <= MUX_s_1_2_2(nand_tmp_139, or_2258_nl, fsm_output(2));
  mux_2094_nl <= MUX_s_1_2_2(mux_tmp_2041, mux_nl, fsm_output(7));
  mux_2100_nl <= MUX_s_1_2_2(mux_2099_nl, mux_2094_nl, fsm_output(5));
  mux_2108_nl <= MUX_s_1_2_2(mux_2107_nl, mux_2100_nl, fsm_output(1));
  mux_2121_nl <= MUX_s_1_2_2(mux_2120_nl, mux_2108_nl, fsm_output(6));
  or_2310_nl <= (fsm_output(4)) OR (fsm_output(7)) OR (NOT (fsm_output(8))) OR (fsm_output(3))
      OR (fsm_output(9));
  or_2309_nl <= (fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(9));
  mux_2149_nl <= MUX_s_1_2_2(or_2310_nl, or_2309_nl, fsm_output(0));
  mux_2150_nl <= MUX_s_1_2_2(mux_2149_nl, mux_tmp_2072, fsm_output(2));
  or_2308_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("01")) OR not_tmp_571;
  mux_2146_nl <= MUX_s_1_2_2(or_2308_nl, or_2306_cse, fsm_output(4));
  mux_2145_nl <= MUX_s_1_2_2(or_tmp_2191, mux_tmp_2081, fsm_output(4));
  mux_2147_nl <= MUX_s_1_2_2(mux_2146_nl, mux_2145_nl, fsm_output(0));
  mux_2144_nl <= MUX_s_1_2_2(mux_tmp_1610, or_tmp_2183, fsm_output(0));
  mux_2148_nl <= MUX_s_1_2_2(mux_2147_nl, mux_2144_nl, fsm_output(2));
  mux_2151_nl <= MUX_s_1_2_2(mux_2150_nl, mux_2148_nl, fsm_output(5));
  or_2305_nl <= (fsm_output(4)) OR (NOT (fsm_output(7))) OR (fsm_output(8)) OR (fsm_output(3))
      OR (fsm_output(9));
  nand_392_nl <= NOT((fsm_output(4)) AND (NOT mux_1583_cse));
  or_2304_nl <= (fsm_output(4)) OR mux_1583_cse;
  mux_2141_nl <= MUX_s_1_2_2(nand_392_nl, or_2304_nl, fsm_output(0));
  mux_2142_nl <= MUX_s_1_2_2(or_2305_nl, mux_2141_nl, fsm_output(2));
  mux_2143_nl <= MUX_s_1_2_2(mux_tmp_2083, mux_2142_nl, fsm_output(5));
  mux_2152_nl <= MUX_s_1_2_2(mux_2151_nl, mux_2143_nl, fsm_output(1));
  mux_2136_nl <= MUX_s_1_2_2(mux_tmp_2081, or_tmp_1788, fsm_output(4));
  mux_2137_nl <= MUX_s_1_2_2(or_tmp_2193, mux_2136_nl, fsm_output(0));
  or_2303_nl <= (fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(8)) OR (fsm_output(3))
      OR (fsm_output(9));
  mux_2138_nl <= MUX_s_1_2_2(mux_2137_nl, or_2303_nl, fsm_output(2));
  mux_2139_nl <= MUX_s_1_2_2(mux_2138_nl, mux_tmp_2083, fsm_output(5));
  mux_2127_nl <= MUX_s_1_2_2(or_tmp_2191, or_tmp_1788, fsm_output(4));
  mux_2126_nl <= MUX_s_1_2_2(or_tmp_1793, mux_tmp_1610, fsm_output(4));
  mux_2128_nl <= MUX_s_1_2_2(mux_2127_nl, mux_2126_nl, fsm_output(0));
  or_2367_nl <= nor_810_cse OR mux_1583_cse;
  mux_2129_nl <= MUX_s_1_2_2(mux_2128_nl, or_2367_nl, fsm_output(2));
  or_2292_nl <= (fsm_output(2)) OR mux_tmp_2072;
  mux_2130_nl <= MUX_s_1_2_2(mux_2129_nl, or_2292_nl, fsm_output(5));
  mux_2140_nl <= MUX_s_1_2_2(mux_2139_nl, mux_2130_nl, fsm_output(1));
  mux_2153_nl <= MUX_s_1_2_2(mux_2152_nl, mux_2140_nl, fsm_output(6));
  or_1923_nl <= (fsm_output(9)) OR mux_tmp_1688;
  or_1922_nl <= (NOT (fsm_output(9))) OR (NOT (fsm_output(2))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR (fsm_output(4));
  mux_1740_nl <= MUX_s_1_2_2(or_1923_nl, or_1922_nl, fsm_output(8));
  or_nl <= mux_1740_nl OR (NOT and_dcpl_17) OR (fsm_output(3)) OR (fsm_output(6));
  or_2316_nl <= (fsm_output(9)) OR (fsm_output(1)) OR (fsm_output(8)) OR (NOT (fsm_output(2)))
      OR (fsm_output(4));
  or_2315_nl <= (NOT (fsm_output(1))) OR (fsm_output(8)) OR (fsm_output(2)) OR (NOT
      (fsm_output(4)));
  or_2313_nl <= (fsm_output(1)) OR (NOT (fsm_output(8))) OR (NOT (fsm_output(2)))
      OR (fsm_output(4));
  mux_2154_nl <= MUX_s_1_2_2(or_2315_nl, or_2313_nl, fsm_output(9));
  mux_2155_nl <= MUX_s_1_2_2(or_2316_nl, mux_2154_nl, fsm_output(0));
  or_2365_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")) OR mux_2155_nl;
  or_2366_nl <= (NOT (fsm_output(7))) OR (NOT (fsm_output(6))) OR (fsm_output(0))
      OR (NOT (fsm_output(9))) OR (NOT (fsm_output(1))) OR (fsm_output(8)) OR (NOT
      (fsm_output(2))) OR (fsm_output(4));
  mux_2156_nl <= MUX_s_1_2_2(or_2365_nl, or_2366_nl, fsm_output(5));
  mux_1747_nl <= MUX_s_1_2_2(or_tmp_1899, or_103_cse, and_267_cse);
  mux_1748_nl <= MUX_s_1_2_2(mux_1747_nl, or_103_cse, fsm_output(2));
  nor_269_nl <= NOT((fsm_output(9)) OR (fsm_output(6)) OR mux_1748_nl);
  mux_1749_nl <= MUX_s_1_2_2(nor_269_nl, and_tmp_12, fsm_output(8));
  mux_1753_nl <= MUX_s_1_2_2((NOT (fsm_output(3))), (fsm_output(3)), fsm_output(4));
  or_1936_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("01"));
  mux_1752_nl <= MUX_s_1_2_2(or_1936_nl, (fsm_output(4)), fsm_output(1));
  mux_1754_nl <= MUX_s_1_2_2(mux_1753_nl, mux_1752_nl, fsm_output(2));
  COMP_LOOP_COMP_LOOP_and_17_nl <= CONV_SL_1_1(z_out_6_10_1(3 DOWNTO 0)=STD_LOGIC_VECTOR'("0011"));
  COMP_LOOP_COMP_LOOP_and_10_nl <= CONV_SL_1_1(VEC_LOOP_j_sva_9_0(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011"));
  COMP_LOOP_1_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(z_out_3 & STD_LOGIC_VECTOR'(
      "0000")) + SIGNED('1' & (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 1)))) + SIGNED'(
      "0000000001"), 10));
  mux_1836_nl <= MUX_s_1_2_2((NOT mux_1834_itm), or_tmp_1989, fsm_output(4));
  mux_1838_nl <= MUX_s_1_2_2(mux_tmp_1786, mux_1836_nl, fsm_output(1));
  or_2033_nl <= (fsm_output(4)) OR (NOT mux_1834_itm);
  mux_1835_nl <= MUX_s_1_2_2(or_2033_nl, mux_tmp_1782, fsm_output(1));
  mux_1839_nl <= MUX_s_1_2_2(mux_1838_nl, mux_1835_nl, fsm_output(0));
  mux_1840_nl <= MUX_s_1_2_2(mux_tmp_1786, mux_1839_nl, fsm_output(2));
  mux_1841_nl <= MUX_s_1_2_2(mux_1840_nl, mux_tmp_1782, fsm_output(3));
  nand_146_nl <= NOT((CONV_SL_1_1(fsm_output(7 DOWNTO 2)/=STD_LOGIC_VECTOR'("000000")))
      AND (fsm_output(9)));
  mux_1842_nl <= MUX_s_1_2_2(mux_1841_nl, nand_146_nl, fsm_output(8));
  nand_338_nl <= NOT((fsm_output(2)) AND or_2186_cse AND (fsm_output(4)) AND (fsm_output(3))
      AND (fsm_output(7)) AND (fsm_output(5)));
  mux_1845_nl <= MUX_s_1_2_2(mux_tmp_1793, nand_338_nl, fsm_output(6));
  or_23_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00"));
  mux_66_nl <= MUX_s_1_2_2(or_tmp_20, or_23_nl, or_2186_cse);
  mux_67_nl <= MUX_s_1_2_2(or_tmp_20, mux_66_nl, fsm_output(2));
  nand_145_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11")));
  mux_1848_nl <= MUX_s_1_2_2(mux_67_nl, nand_145_nl, fsm_output(6));
  mux_1855_nl <= MUX_s_1_2_2(mux_tmp_1803, mux_tmp_1801, fsm_output(0));
  mux_1849_nl <= MUX_s_1_2_2(nor_tmp_40, (fsm_output(7)), fsm_output(3));
  mux_1851_nl <= MUX_s_1_2_2(mux_tmp_1799, mux_1849_nl, fsm_output(4));
  mux_1853_nl <= MUX_s_1_2_2(mux_tmp_1801, mux_1851_nl, fsm_output(0));
  mux_1856_nl <= MUX_s_1_2_2(mux_1855_nl, mux_1853_nl, fsm_output(1));
  mux_1857_nl <= MUX_s_1_2_2(mux_tmp_1803, mux_1856_nl, fsm_output(2));
  mux_1858_nl <= MUX_s_1_2_2(mux_1857_nl, (fsm_output(7)), fsm_output(6));
  mux_1861_nl <= MUX_s_1_2_2(mux_tmp_1809, mux_tmp_1808, and_418_cse);
  mux_1862_nl <= MUX_s_1_2_2(mux_tmp_1793, (NOT mux_1861_nl), fsm_output(6));
  mux_1864_nl <= MUX_s_1_2_2((fsm_output(7)), or_tmp_74, fsm_output(4));
  mux_1863_nl <= MUX_s_1_2_2((fsm_output(7)), or_tmp_74, or_2040_cse);
  mux_1865_nl <= MUX_s_1_2_2(mux_1864_nl, mux_1863_nl, fsm_output(2));
  or_2041_nl <= (fsm_output(6)) OR mux_1865_nl;
  mux_1866_nl <= MUX_s_1_2_2(not_tmp_431, or_2041_nl, fsm_output(8));
  or_2043_nl <= ((fsm_output(1)) AND (fsm_output(0)) AND (fsm_output(4)) AND (fsm_output(3)))
      OR (fsm_output(7)) OR (fsm_output(5));
  mux_1867_nl <= MUX_s_1_2_2(or_2043_nl, or_tmp_1899, fsm_output(2));
  mux_1868_nl <= MUX_s_1_2_2((fsm_output(7)), mux_1867_nl, fsm_output(6));
  mux_1869_nl <= MUX_s_1_2_2(not_tmp_431, mux_1868_nl, fsm_output(8));
  or_2175_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  mux_1870_nl <= MUX_s_1_2_2(mux_tmp_1809, mux_tmp_1808, or_2175_nl);
  mux_1871_nl <= MUX_s_1_2_2(mux_1870_nl, (fsm_output(7)), fsm_output(6));
  mux_1872_nl <= MUX_s_1_2_2(not_tmp_431, mux_1871_nl, fsm_output(8));
  and_248_nl <= (CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))) AND
      (fsm_output(4)) AND (fsm_output(3)) AND (fsm_output(7)) AND (fsm_output(5));
  mux_1873_nl <= MUX_s_1_2_2(and_248_nl, (fsm_output(7)), fsm_output(6));
  mux_1874_nl <= MUX_s_1_2_2(not_tmp_431, mux_1873_nl, fsm_output(8));
  and_213_nl <= (fsm_output(6)) AND or_2040_cse AND (fsm_output(7)) AND (fsm_output(5));
  mux_1875_nl <= MUX_s_1_2_2(not_tmp_431, and_213_nl, fsm_output(8));
  mux_1876_nl <= MUX_s_1_2_2(or_tmp_1899, or_103_cse, and_247_cse);
  or_2047_nl <= (fsm_output(6)) OR mux_1876_nl;
  mux_1877_nl <= MUX_s_1_2_2(not_tmp_431, or_2047_nl, fsm_output(9));
  mux_1879_nl <= MUX_s_1_2_2((fsm_output(7)), or_tmp_1845, fsm_output(6));
  mux_1880_nl <= MUX_s_1_2_2(not_tmp_431, mux_1879_nl, fsm_output(9));
  mux_1882_nl <= MUX_s_1_2_2(not_tmp_439, nor_tmp_215, or_2186_cse);
  mux_1883_nl <= MUX_s_1_2_2(not_tmp_439, mux_1882_nl, fsm_output(2));
  mux_1884_nl <= MUX_s_1_2_2(mux_1883_nl, nor_tmp_215, fsm_output(3));
  mux_1885_nl <= MUX_s_1_2_2(not_tmp_439, mux_1884_nl, fsm_output(4));
  or_110_nl <= CONV_SL_1_1(fsm_output(8 DOWNTO 7)/=STD_LOGIC_VECTOR'("00"));
  and_245_nl <= (CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"))) AND
      (fsm_output(7)) AND (fsm_output(5));
  mux_1887_nl <= MUX_s_1_2_2(and_245_nl, (fsm_output(7)), fsm_output(6));
  mux_1888_nl <= MUX_s_1_2_2(not_tmp_431, mux_1887_nl, fsm_output(9));
  mux_1892_nl <= MUX_s_1_2_2(not_tmp_418, mux_tmp_1839, and_267_cse);
  mux_1891_nl <= MUX_s_1_2_2(mux_tmp_1839, nor_tmp_203, or_2186_cse);
  mux_1893_nl <= MUX_s_1_2_2(mux_1892_nl, mux_1891_nl, fsm_output(2));
  mux_1894_nl <= MUX_s_1_2_2(mux_1893_nl, nor_tmp_203, fsm_output(3));
  mux_1895_nl <= MUX_s_1_2_2(not_tmp_418, mux_1894_nl, fsm_output(4));
  mux_1896_nl <= MUX_s_1_2_2(mux_1895_nl, nor_tmp_203, fsm_output(5));
  nor_nl <= NOT((fsm_output(9)) OR (fsm_output(6)) OR mux_tmp_1793);
  and_nl <= (fsm_output(9)) AND (CONV_SL_1_1(fsm_output(7 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000000")));
  COMP_LOOP_or_6_nl <= (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_221);
  COMP_LOOP_or_7_nl <= (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_nor_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_221);
  COMP_LOOP_or_8_nl <= (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_dcpl_221);
  COMP_LOOP_or_9_nl <= (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_201) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_221);
  COMP_LOOP_or_10_nl <= (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_221);
  COMP_LOOP_or_11_nl <= (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_203) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_221);
  COMP_LOOP_or_12_nl <= (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_221);
  COMP_LOOP_or_13_nl <= (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_206) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_221);
  COMP_LOOP_or_14_nl <= (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_221);
  COMP_LOOP_or_15_nl <= (COMP_LOOP_COMP_LOOP_and_8_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_210) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_221);
  COMP_LOOP_or_16_nl <= (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_221);
  COMP_LOOP_or_17_nl <= (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_214) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_221);
  COMP_LOOP_or_18_nl <= (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_221);
  COMP_LOOP_or_19_nl <= (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_217) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_221);
  COMP_LOOP_or_20_nl <= (COMP_LOOP_COMP_LOOP_and_13_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_12_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_11_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_10_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_9_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_8_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_68_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_6_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_5_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_4_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_64_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_2_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_62_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_244_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_220) OR (COMP_LOOP_COMP_LOOP_and_14_itm
      AND and_dcpl_221);
  COMP_LOOP_or_21_nl <= (COMP_LOOP_COMP_LOOP_and_14_itm AND and_dcpl_199) OR (COMP_LOOP_COMP_LOOP_and_13_itm
      AND and_dcpl_200) OR (COMP_LOOP_COMP_LOOP_and_12_itm AND and_dcpl_201) OR (COMP_LOOP_COMP_LOOP_and_11_itm
      AND and_dcpl_202) OR (COMP_LOOP_COMP_LOOP_and_10_itm AND and_dcpl_203) OR (COMP_LOOP_COMP_LOOP_and_9_itm
      AND and_dcpl_204) OR (COMP_LOOP_COMP_LOOP_and_8_itm AND and_dcpl_206) OR (COMP_LOOP_COMP_LOOP_and_68_itm
      AND and_dcpl_208) OR (COMP_LOOP_COMP_LOOP_and_6_itm AND and_dcpl_210) OR (COMP_LOOP_COMP_LOOP_and_5_itm
      AND and_dcpl_212) OR (COMP_LOOP_COMP_LOOP_and_4_itm AND and_dcpl_214) OR (COMP_LOOP_COMP_LOOP_and_64_itm
      AND and_dcpl_215) OR (COMP_LOOP_COMP_LOOP_and_2_itm AND and_dcpl_217) OR (COMP_LOOP_COMP_LOOP_and_62_itm
      AND and_dcpl_219) OR (COMP_LOOP_COMP_LOOP_and_244_itm AND and_dcpl_220) OR
      (COMP_LOOP_COMP_LOOP_nor_itm AND and_dcpl_221);
  not_nl <= NOT mux_1911_cse;
  mux_2193_nl <= MUX_s_1_2_2(or_tmp_2227, or_tmp_2041, fsm_output(7));
  mux_2194_nl <= MUX_s_1_2_2(mux_2193_nl, mux_tmp_2124, fsm_output(6));
  mux_2195_nl <= MUX_s_1_2_2(mux_2194_nl, mux_tmp_2119, fsm_output(0));
  mux_2189_nl <= MUX_s_1_2_2(mux_1949_cse, or_tmp_2041, fsm_output(1));
  mux_2190_nl <= MUX_s_1_2_2(mux_2189_nl, mux_tmp_2108, fsm_output(7));
  mux_2191_nl <= MUX_s_1_2_2(mux_2190_nl, mux_tmp_2112, fsm_output(6));
  mux_2185_nl <= MUX_s_1_2_2(mux_1922_cse, mux_1920_cse, fsm_output(1));
  mux_2186_nl <= MUX_s_1_2_2(or_tmp_2223, mux_2185_nl, fsm_output(7));
  mux_2187_nl <= MUX_s_1_2_2(mux_tmp_2128, mux_2186_nl, fsm_output(6));
  mux_2192_nl <= MUX_s_1_2_2(mux_2191_nl, mux_2187_nl, fsm_output(0));
  mux_2196_nl <= MUX_s_1_2_2(mux_2195_nl, mux_2192_nl, fsm_output(5));
  mux_2181_nl <= MUX_s_1_2_2(nand_tmp_134, or_tmp_2223, fsm_output(7));
  mux_2182_nl <= MUX_s_1_2_2(mux_2181_nl, mux_tmp_2128, fsm_output(6));
  mux_2173_nl <= MUX_s_1_2_2(mux_tmp_1861, or_2336_cse, fsm_output(1));
  mux_2174_nl <= MUX_s_1_2_2(or_tmp_2041, mux_2173_nl, fsm_output(7));
  mux_2177_nl <= MUX_s_1_2_2(mux_tmp_2124, mux_2174_nl, fsm_output(6));
  mux_2183_nl <= MUX_s_1_2_2(mux_2182_nl, mux_2177_nl, fsm_output(0));
  mux_2157_nl <= MUX_s_1_2_2(or_tmp_2037, or_1916_cse, fsm_output(1));
  mux_2161_nl <= MUX_s_1_2_2(mux_tmp_2108, mux_2157_nl, fsm_output(7));
  mux_2165_nl <= MUX_s_1_2_2(mux_tmp_2112, mux_2161_nl, fsm_output(6));
  mux_2172_nl <= MUX_s_1_2_2(mux_tmp_2119, mux_2165_nl, fsm_output(0));
  mux_2184_nl <= MUX_s_1_2_2(mux_2183_nl, mux_2172_nl, fsm_output(5));
  or_2347_nl <= (fsm_output(2)) OR (NOT (fsm_output(8))) OR (fsm_output(9));
  mux_2237_nl <= MUX_s_1_2_2(or_2347_nl, mux_tmp_2179, fsm_output(3));
  mux_2238_nl <= MUX_s_1_2_2(mux_2237_nl, mux_tmp_2180, fsm_output(0));
  mux_2239_nl <= MUX_s_1_2_2(or_212_cse, mux_2238_nl, fsm_output(4));
  mux_2236_nl <= MUX_s_1_2_2(mux_1949_cse, or_212_cse, fsm_output(4));
  mux_2240_nl <= MUX_s_1_2_2(mux_2239_nl, mux_2236_nl, fsm_output(5));
  mux_2233_nl <= MUX_s_1_2_2(mux_tmp_2180, mux_tmp_1861, fsm_output(0));
  mux_2230_nl <= MUX_s_1_2_2(mux_1949_cse, mux_tmp_2167, fsm_output(0));
  mux_2234_nl <= MUX_s_1_2_2(mux_2233_nl, mux_2230_nl, fsm_output(4));
  mux_2235_nl <= MUX_s_1_2_2(mux_2234_nl, mux_tmp_2170, fsm_output(5));
  mux_2241_nl <= MUX_s_1_2_2(mux_2240_nl, mux_2235_nl, fsm_output(6));
  mux_2227_nl <= MUX_s_1_2_2(mux_tmp_2169, mux_tmp_2165, fsm_output(5));
  mux_2226_nl <= MUX_s_1_2_2(mux_tmp_2164, mux_tmp_2159, fsm_output(5));
  mux_2228_nl <= MUX_s_1_2_2(mux_2227_nl, mux_2226_nl, fsm_output(6));
  mux_2242_nl <= MUX_s_1_2_2(mux_2241_nl, mux_2228_nl, fsm_output(7));
  mux_2223_nl <= MUX_s_1_2_2(mux_tmp_2170, mux_tmp_2169, fsm_output(5));
  mux_2218_nl <= MUX_s_1_2_2(mux_tmp_2165, mux_tmp_2164, fsm_output(5));
  mux_2224_nl <= MUX_s_1_2_2(mux_2223_nl, mux_2218_nl, fsm_output(6));
  mux_2209_nl <= MUX_s_1_2_2(mux_tmp_2156, mux_tmp_2150, fsm_output(0));
  mux_2207_nl <= MUX_s_1_2_2(mux_tmp_2154, mux_1922_cse, fsm_output(0));
  mux_2210_nl <= MUX_s_1_2_2(mux_2209_nl, mux_2207_nl, fsm_output(4));
  mux_2212_nl <= MUX_s_1_2_2(mux_tmp_2159, mux_2210_nl, fsm_output(5));
  mux_2203_nl <= MUX_s_1_2_2(or_tmp_2037, mux_tmp_2150, fsm_output(4));
  mux_2198_nl <= MUX_s_1_2_2(or_tmp_2044, or_212_cse, fsm_output(3));
  mux_2200_nl <= MUX_s_1_2_2(mux_1922_cse, mux_2198_nl, fsm_output(0));
  mux_2201_nl <= MUX_s_1_2_2(mux_2200_nl, or_tmp_2037, fsm_output(4));
  mux_2204_nl <= MUX_s_1_2_2(mux_2203_nl, mux_2201_nl, fsm_output(5));
  mux_2213_nl <= MUX_s_1_2_2(mux_2212_nl, mux_2204_nl, fsm_output(6));
  mux_2225_nl <= MUX_s_1_2_2(mux_2224_nl, mux_2213_nl, fsm_output(7));
  mux_2243_nl <= MUX_s_1_2_2(mux_2242_nl, mux_2225_nl, fsm_output(1));
  nand_396_nl <= NOT((fsm_output(6)) AND (fsm_output(4)) AND (fsm_output(0)) AND
      (fsm_output(5)) AND (fsm_output(1)));
  mux_2259_nl <= MUX_s_1_2_2(mux_tmp_2204, mux_tmp_2199, fsm_output(6));
  mux_2260_nl <= MUX_s_1_2_2(nand_396_nl, mux_2259_nl, fsm_output(2));
  nand_397_nl <= NOT(((fsm_output(0)) OR (fsm_output(5))) AND (fsm_output(1)));
  mux_2257_nl <= MUX_s_1_2_2(nand_397_nl, or_tmp_2245, fsm_output(4));
  mux_2258_nl <= MUX_s_1_2_2(mux_2257_nl, mux_tmp_2204, fsm_output(6));
  or_2362_nl <= (fsm_output(2)) OR mux_2258_nl;
  mux_2261_nl <= MUX_s_1_2_2(mux_2260_nl, or_2362_nl, fsm_output(7));
  nor_797_nl <= NOT((fsm_output(3)) OR mux_2261_nl);
  and_700_nl <= (fsm_output(7)) AND (fsm_output(2)) AND (NOT mux_2249_itm);
  mux_2253_nl <= MUX_s_1_2_2(mux_tmp_2196, mux_tmp_2193, fsm_output(6));
  nor_798_nl <= NOT((fsm_output(2)) OR mux_2253_nl);
  nor_799_nl <= NOT((fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(0))
      OR (fsm_output(1)));
  mux_2254_nl <= MUX_s_1_2_2(nor_798_nl, nor_799_nl, fsm_output(7));
  mux_2255_nl <= MUX_s_1_2_2(and_700_nl, mux_2254_nl, fsm_output(3));
  mux_2262_nl <= MUX_s_1_2_2(nor_797_nl, mux_2255_nl, fsm_output(9));
  or_2356_nl <= (fsm_output(7)) OR (fsm_output(2)) OR (fsm_output(6)) OR mux_tmp_2199;
  nand_394_nl <= NOT((fsm_output(2)) AND (NOT mux_2249_itm));
  nand_398_nl <= NOT((fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(5)) AND
      (fsm_output(1)));
  mux_2246_nl <= MUX_s_1_2_2(mux_tmp_2193, or_2348_cse, fsm_output(6));
  mux_2247_nl <= MUX_s_1_2_2(nand_398_nl, mux_2246_nl, fsm_output(2));
  mux_2250_nl <= MUX_s_1_2_2(nand_394_nl, mux_2247_nl, fsm_output(7));
  mux_2252_nl <= MUX_s_1_2_2(or_2356_nl, mux_2250_nl, fsm_output(3));
  nor_800_nl <= NOT((fsm_output(9)) OR mux_2252_nl);
  COMP_LOOP_or_27_nl <= and_dcpl_52 OR and_dcpl_97;
  COMP_LOOP_COMP_LOOP_or_3_nl <= (VEC_LOOP_j_sva_9_0(9)) OR and_dcpl_242 OR and_dcpl_246
      OR and_dcpl_252 OR and_dcpl_255 OR and_dcpl_260 OR and_dcpl_267 OR and_dcpl_272
      OR and_dcpl_274 OR and_dcpl_279 OR and_dcpl_281 OR and_dcpl_284;
  COMP_LOOP_or_52_nl <= and_dcpl_242 OR and_dcpl_246 OR and_dcpl_252 OR and_dcpl_255
      OR and_dcpl_260 OR and_dcpl_267 OR and_dcpl_272 OR and_dcpl_274 OR and_dcpl_279
      OR and_dcpl_281 OR and_dcpl_284;
  COMP_LOOP_COMP_LOOP_mux_15_nl <= MUX_v_9_2_2((VEC_LOOP_j_sva_9_0(8 DOWNTO 0)),
      (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 1))), COMP_LOOP_or_52_nl);
  COMP_LOOP_or_53_nl <= (NOT and_dcpl_238) OR and_dcpl_242 OR and_dcpl_246 OR and_dcpl_252
      OR and_dcpl_255 OR and_dcpl_260 OR and_dcpl_267 OR and_dcpl_272 OR and_dcpl_274
      OR and_dcpl_279 OR and_dcpl_281 OR and_dcpl_284;
  COMP_LOOP_or_54_nl <= and_dcpl_238 OR and_dcpl_255;
  COMP_LOOP_mux1h_271_nl <= MUX1HOT_v_4_11_2(STD_LOGIC_VECTOR'( "0101"), STD_LOGIC_VECTOR'(
      "0001"), STD_LOGIC_VECTOR'( "0010"), STD_LOGIC_VECTOR'( "0100"), STD_LOGIC_VECTOR'(
      "0110"), STD_LOGIC_VECTOR'( "1000"), STD_LOGIC_VECTOR'( "1001"), STD_LOGIC_VECTOR'(
      "1010"), STD_LOGIC_VECTOR'( "1100"), STD_LOGIC_VECTOR'( "1101"), STD_LOGIC_VECTOR'(
      "1110"), STD_LOGIC_VECTOR'( COMP_LOOP_or_54_nl & and_dcpl_242 & and_dcpl_246
      & and_dcpl_252 & and_dcpl_260 & and_dcpl_267 & and_dcpl_272 & and_dcpl_274
      & and_dcpl_279 & and_dcpl_281 & and_dcpl_284));
  acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_3_nl &
      COMP_LOOP_COMP_LOOP_mux_15_nl & COMP_LOOP_or_53_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
      & COMP_LOOP_mux1h_271_nl & '1'), 10), 11), 11));
  z_out_1 <= acc_nl(10 DOWNTO 1);
  COMP_LOOP_COMP_LOOP_or_4_nl <= (VEC_LOOP_j_sva_9_0(9)) OR and_dcpl_300 OR and_dcpl_308;
  COMP_LOOP_or_55_nl <= and_dcpl_300 OR and_dcpl_308;
  COMP_LOOP_COMP_LOOP_mux_16_nl <= MUX_v_7_2_2((VEC_LOOP_j_sva_9_0(8 DOWNTO 2)),
      (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 3))), COMP_LOOP_or_55_nl);
  COMP_LOOP_or_56_nl <= (NOT and_dcpl_293) OR and_dcpl_300 OR and_dcpl_308;
  COMP_LOOP_COMP_LOOP_or_5_nl <= (NOT and_dcpl_300) OR and_dcpl_293;
  acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_COMP_LOOP_or_4_nl
      & COMP_LOOP_COMP_LOOP_mux_16_nl & COMP_LOOP_or_56_nl) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
      & COMP_LOOP_COMP_LOOP_or_5_nl & and_dcpl_293 & '1'), 8), 9), 9));
  z_out_2 <= acc_1_nl(8 DOWNTO 1);
  operator_64_false_1_mux_1_nl <= MUX_v_5_2_2((NOT COMP_LOOP_k_9_4_sva_4_0), COMP_LOOP_k_9_4_sva_4_0,
      and_551_ssc);
  z_out_3 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED((NOT and_551_ssc) & operator_64_false_1_mux_1_nl)
      + UNSIGNED'( "000001"), 6));
  COMP_LOOP_mux_35_nl <= MUX_v_6_2_2(('1' & (NOT (STAGE_LOOP_lshift_psp_sva(9 DOWNTO
      5)))), (VEC_LOOP_j_sva_9_0(9 DOWNTO 4)), and_dcpl_344);
  COMP_LOOP_COMP_LOOP_nand_1_nl <= NOT(and_dcpl_344 AND (NOT(CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("1010110111")))));
  acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_35_nl & COMP_LOOP_COMP_LOOP_nand_1_nl)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & '1'), 6),
      7), 7));
  z_out_4 <= acc_3_nl(6 DOWNTO 1);
  COMP_LOOP_mux_36_nl <= MUX_v_7_2_2((VEC_LOOP_j_sva_9_0(9 DOWNTO 3)), ('1' & (NOT
      (STAGE_LOOP_lshift_psp_sva(9 DOWNTO 4)))), and_dcpl_361);
  COMP_LOOP_or_57_nl <= (NOT(and_dcpl_236 AND and_dcpl_234 AND nor_761_cse AND (NOT
      (fsm_output(0))) AND (fsm_output(4)))) OR and_dcpl_361;
  acc_4_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_mux_36_nl & COMP_LOOP_or_57_nl)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0 & (NOT and_dcpl_361)
      & '1'), 7), 8), 8));
  z_out_5 <= acc_4_nl(7 DOWNTO 1);
  and_706_nl <= and_dcpl_251 AND and_dcpl_376 AND (NOT (fsm_output(5))) AND and_dcpl_32;
  and_707_nl <= and_dcpl_251 AND and_dcpl_382 AND and_dcpl_29;
  and_708_nl <= and_dcpl_70 AND (NOT (fsm_output(3))) AND and_dcpl_256 AND and_dcpl_232
      AND and_dcpl_29;
  and_709_nl <= and_dcpl_398 AND and_dcpl_396;
  and_710_nl <= and_dcpl_398 AND and_dcpl_403;
  and_711_nl <= and_dcpl_407 AND and_dcpl_232 AND and_dcpl_66;
  and_712_nl <= and_dcpl_407 AND and_dcpl_244 AND and_dcpl_16;
  and_713_nl <= and_dcpl_265 AND and_dcpl_250 AND and_dcpl_402 AND and_dcpl_66;
  and_714_nl <= and_dcpl_417 AND and_dcpl_382 AND and_dcpl_16;
  and_715_nl <= and_dcpl_417 AND and_dcpl_244 AND and_dcpl_66;
  and_716_nl <= and_dcpl_416 AND and_dcpl_250 AND and_dcpl_232 AND and_dcpl_16;
  and_717_nl <= and_dcpl_425 AND and_dcpl_396;
  COMP_LOOP_mux1h_272_nl <= MUX1HOT_v_4_14_2(STD_LOGIC_VECTOR'( "1110"), STD_LOGIC_VECTOR'(
      "1101"), STD_LOGIC_VECTOR'( "1100"), STD_LOGIC_VECTOR'( "1011"), STD_LOGIC_VECTOR'(
      "1010"), STD_LOGIC_VECTOR'( "1001"), STD_LOGIC_VECTOR'( "1000"), STD_LOGIC_VECTOR'(
      "0111"), STD_LOGIC_VECTOR'( "0110"), STD_LOGIC_VECTOR'( "0101"), STD_LOGIC_VECTOR'(
      "0100"), STD_LOGIC_VECTOR'( "0011"), STD_LOGIC_VECTOR'( "0010"), STD_LOGIC_VECTOR'(
      "0001"), STD_LOGIC_VECTOR'( and_dcpl_246 & and_706_nl & and_707_nl & and_dcpl_255
      & and_708_nl & and_709_nl & and_710_nl & and_711_nl & and_712_nl & and_713_nl
      & and_714_nl & and_715_nl & and_716_nl & and_717_nl));
  COMP_LOOP_COMP_LOOP_nor_63_nl <= NOT(MUX_v_4_2_2(COMP_LOOP_mux1h_272_nl, STD_LOGIC_VECTOR'("1111"),
      and_dcpl_242));
  and_718_nl <= and_dcpl_425 AND and_dcpl_403;
  COMP_LOOP_or_58_nl <= MUX_v_4_2_2(COMP_LOOP_COMP_LOOP_nor_63_nl, STD_LOGIC_VECTOR'("1111"),
      and_718_nl);
  acc_5_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(COMP_LOOP_k_9_4_sva_4_0
      & COMP_LOOP_or_58_nl), 9), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(VEC_LOOP_j_sva_9_0),
      10), 11) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_lshift_psp_sva),
      10), 11), 11));
  z_out_6_10_1 <= acc_5_nl(10 DOWNTO 1);
  STAGE_LOOP_STAGE_LOOP_or_1_nl <= (NOT((fsm_output(9)) AND (fsm_output(8)) AND (NOT
      (fsm_output(3))) AND and_dcpl_234 AND (fsm_output(1)) AND (NOT (fsm_output(6)))
      AND (NOT (fsm_output(5))) AND (NOT (fsm_output(0))) AND (NOT (fsm_output(4)))))
      OR (NOT mux_2066_cse) OR and_dcpl_444;
  STAGE_LOOP_or_2_nl <= (NOT mux_2066_cse) OR and_dcpl_444;
  STAGE_LOOP_STAGE_LOOP_mux_2_nl <= MUX_v_64_2_2((STD_LOGIC_VECTOR'( "000000000000000000000000000000000000000000000000000000000000")
      & STAGE_LOOP_i_3_0_sva), (NOT (z_out_9(63 DOWNTO 0))), STAGE_LOOP_or_2_nl);
  z_out_7 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(STAGE_LOOP_STAGE_LOOP_or_1_nl
      & STAGE_LOOP_STAGE_LOOP_mux_2_nl) + UNSIGNED'( "00000000000000000000000000000000000000000000000000000000000000001"),
      65));
  operator_64_false_operator_64_false_operator_64_false_nor_1_nl <= NOT(MUX_v_61_2_2((operator_66_true_div_cmp_z(63
      DOWNTO 3)), STD_LOGIC_VECTOR'("1111111111111111111111111111111111111111111111111111111111111"),
      and_dcpl_460));
  operator_64_false_mux_1_nl <= MUX_v_3_2_2((NOT (operator_66_true_div_cmp_z(2 DOWNTO
      0))), (z_out_7(3 DOWNTO 1)), and_dcpl_460);
  operator_64_false_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED((NOT and_dcpl_460)
      & operator_64_false_operator_64_false_operator_64_false_nor_1_nl & operator_64_false_mux_1_nl)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( and_dcpl_460 & '1'), 2), 65), 65));
  z_out_8_64_2 <= operator_64_false_acc_nl(64 DOWNTO 2);
  and_719_nl <= and_dcpl_236 AND and_dcpl_256 AND and_dcpl_464;
  and_720_nl <= and_dcpl_236 AND (NOT (fsm_output(7))) AND (fsm_output(2)) AND and_dcpl_464;
  operator_64_false_mux1h_1_nl <= MUX1HOT_v_64_3_2(p_sva, modExp_dev_exp_sva, (modExp_dev_exp_1_sva_63_9
      & COMP_LOOP_acc_10_cse_10_1_1_sva_4_0 & modExp_dev_exp_1_sva_3_0), STD_LOGIC_VECTOR'(
      and_719_nl & and_720_nl & (NOT mux_2066_cse)));
  z_out_9 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(operator_64_false_mux1h_1_nl),
      65) + UNSIGNED'( "11111111111111111111111111111111111111111111111111111111111111111"),
      65));
END v11;

-- ------------------------------------------------------------------
--  Design Unit:    inPlaceNTT_DIT
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;


ENTITY inPlaceNTT_DIT IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    vec_rsc_0_0_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_0_we : OUT STD_LOGIC;
    vec_rsc_0_0_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_0_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    vec_rsc_0_1_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_1_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_1_we : OUT STD_LOGIC;
    vec_rsc_0_1_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_1_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    vec_rsc_0_2_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_2_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_2_we : OUT STD_LOGIC;
    vec_rsc_0_2_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_2_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    vec_rsc_0_3_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_3_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_3_we : OUT STD_LOGIC;
    vec_rsc_0_3_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_3_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    vec_rsc_0_4_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_4_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_4_we : OUT STD_LOGIC;
    vec_rsc_0_4_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_4_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    vec_rsc_0_5_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_5_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_5_we : OUT STD_LOGIC;
    vec_rsc_0_5_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_5_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    vec_rsc_0_6_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_6_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_6_we : OUT STD_LOGIC;
    vec_rsc_0_6_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_6_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    vec_rsc_0_7_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_7_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_7_we : OUT STD_LOGIC;
    vec_rsc_0_7_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_7_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    vec_rsc_0_8_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_8_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_8_we : OUT STD_LOGIC;
    vec_rsc_0_8_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_8_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    vec_rsc_0_9_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_9_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_9_we : OUT STD_LOGIC;
    vec_rsc_0_9_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_9_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    vec_rsc_0_10_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_10_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_10_we : OUT STD_LOGIC;
    vec_rsc_0_10_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_10_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    vec_rsc_0_11_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_11_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_11_we : OUT STD_LOGIC;
    vec_rsc_0_11_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_11_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    vec_rsc_0_12_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_12_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_12_we : OUT STD_LOGIC;
    vec_rsc_0_12_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_12_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    vec_rsc_0_13_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_13_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_13_we : OUT STD_LOGIC;
    vec_rsc_0_13_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_13_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    vec_rsc_0_14_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_14_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_14_we : OUT STD_LOGIC;
    vec_rsc_0_14_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_14_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    vec_rsc_0_15_wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_15_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_0_15_we : OUT STD_LOGIC;
    vec_rsc_0_15_radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    vec_rsc_0_15_q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC
  );
END inPlaceNTT_DIT;

ARCHITECTURE v11 OF inPlaceNTT_DIT IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL vec_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL vec_rsc_0_0_i_d_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr_d_iff : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_1_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_2_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_3_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_4_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_5_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_6_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_7_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_8_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_9_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_10_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_11_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_12_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_13_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_14_i_we_d_iff : STD_LOGIC;
  SIGNAL vec_rsc_0_15_i_we_d_iff : STD_LOGIC;

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_0_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_0_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_1_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_1_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_2_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_2_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_3_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_3_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_4_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_4_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_5_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_5_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_6_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_6_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_7_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_7_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_8_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_8_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_9_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_9_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_10_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_10_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_11_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_11_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_12_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_12_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_13_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_13_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_14_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_14_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      d_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL vec_rsc_0_15_i_q : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_radr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_wadr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_d_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_q_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_radr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL vec_rsc_0_15_i_wadr_d : STD_LOGIC_VECTOR (5 DOWNTO 0);

  COMPONENT inPlaceNTT_DIT_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      vec_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      vec_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_dat : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      r_rsc_triosy_lz : OUT STD_LOGIC;
      vec_rsc_0_0_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_1_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_2_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_3_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_4_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_5_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_6_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_7_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_8_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_9_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_10_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_11_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_12_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_13_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_14_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_15_i_q_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      vec_rsc_0_0_i_d_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      vec_rsc_0_0_i_radr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      vec_rsc_0_0_i_wadr_d_pff : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      vec_rsc_0_0_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_1_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_2_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_3_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_4_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_5_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_6_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_7_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_8_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_9_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_10_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_11_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_12_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_13_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_14_i_we_d_pff : OUT STD_LOGIC;
      vec_rsc_0_15_i_we_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL inPlaceNTT_DIT_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_r_rsc_dat : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_q_d : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_d_d_pff : STD_LOGIC_VECTOR (63 DOWNTO
      0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_radr_d_pff : STD_LOGIC_VECTOR (5
      DOWNTO 0);
  SIGNAL inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_wadr_d_pff : STD_LOGIC_VECTOR (5
      DOWNTO 0);

BEGIN
  vec_rsc_0_0_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_8_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_0_i_q,
      radr => vec_rsc_0_0_i_radr,
      we => vec_rsc_0_0_we,
      d => vec_rsc_0_0_i_d,
      wadr => vec_rsc_0_0_i_wadr,
      d_d => vec_rsc_0_0_i_d_d,
      q_d => vec_rsc_0_0_i_q_d_1,
      radr_d => vec_rsc_0_0_i_radr_d,
      wadr_d => vec_rsc_0_0_i_wadr_d,
      we_d => vec_rsc_0_0_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_0_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_0_i_q <= vec_rsc_0_0_q;
  vec_rsc_0_0_radr <= vec_rsc_0_0_i_radr;
  vec_rsc_0_0_d <= vec_rsc_0_0_i_d;
  vec_rsc_0_0_wadr <= vec_rsc_0_0_i_wadr;
  vec_rsc_0_0_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_0_i_q_d <= vec_rsc_0_0_i_q_d_1;
  vec_rsc_0_0_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_0_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_1_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_1_i_q,
      radr => vec_rsc_0_1_i_radr,
      we => vec_rsc_0_1_we,
      d => vec_rsc_0_1_i_d,
      wadr => vec_rsc_0_1_i_wadr,
      d_d => vec_rsc_0_1_i_d_d,
      q_d => vec_rsc_0_1_i_q_d_1,
      radr_d => vec_rsc_0_1_i_radr_d,
      wadr_d => vec_rsc_0_1_i_wadr_d,
      we_d => vec_rsc_0_1_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_1_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_1_i_q <= vec_rsc_0_1_q;
  vec_rsc_0_1_radr <= vec_rsc_0_1_i_radr;
  vec_rsc_0_1_d <= vec_rsc_0_1_i_d;
  vec_rsc_0_1_wadr <= vec_rsc_0_1_i_wadr;
  vec_rsc_0_1_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_1_i_q_d <= vec_rsc_0_1_i_q_d_1;
  vec_rsc_0_1_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_1_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_2_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_2_i_q,
      radr => vec_rsc_0_2_i_radr,
      we => vec_rsc_0_2_we,
      d => vec_rsc_0_2_i_d,
      wadr => vec_rsc_0_2_i_wadr,
      d_d => vec_rsc_0_2_i_d_d,
      q_d => vec_rsc_0_2_i_q_d_1,
      radr_d => vec_rsc_0_2_i_radr_d,
      wadr_d => vec_rsc_0_2_i_wadr_d,
      we_d => vec_rsc_0_2_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_2_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_2_i_q <= vec_rsc_0_2_q;
  vec_rsc_0_2_radr <= vec_rsc_0_2_i_radr;
  vec_rsc_0_2_d <= vec_rsc_0_2_i_d;
  vec_rsc_0_2_wadr <= vec_rsc_0_2_i_wadr;
  vec_rsc_0_2_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_2_i_q_d <= vec_rsc_0_2_i_q_d_1;
  vec_rsc_0_2_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_2_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_3_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_3_i_q,
      radr => vec_rsc_0_3_i_radr,
      we => vec_rsc_0_3_we,
      d => vec_rsc_0_3_i_d,
      wadr => vec_rsc_0_3_i_wadr,
      d_d => vec_rsc_0_3_i_d_d,
      q_d => vec_rsc_0_3_i_q_d_1,
      radr_d => vec_rsc_0_3_i_radr_d,
      wadr_d => vec_rsc_0_3_i_wadr_d,
      we_d => vec_rsc_0_3_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_3_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_3_i_q <= vec_rsc_0_3_q;
  vec_rsc_0_3_radr <= vec_rsc_0_3_i_radr;
  vec_rsc_0_3_d <= vec_rsc_0_3_i_d;
  vec_rsc_0_3_wadr <= vec_rsc_0_3_i_wadr;
  vec_rsc_0_3_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_3_i_q_d <= vec_rsc_0_3_i_q_d_1;
  vec_rsc_0_3_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_3_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_4_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_4_i_q,
      radr => vec_rsc_0_4_i_radr,
      we => vec_rsc_0_4_we,
      d => vec_rsc_0_4_i_d,
      wadr => vec_rsc_0_4_i_wadr,
      d_d => vec_rsc_0_4_i_d_d,
      q_d => vec_rsc_0_4_i_q_d_1,
      radr_d => vec_rsc_0_4_i_radr_d,
      wadr_d => vec_rsc_0_4_i_wadr_d,
      we_d => vec_rsc_0_4_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_4_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_4_i_q <= vec_rsc_0_4_q;
  vec_rsc_0_4_radr <= vec_rsc_0_4_i_radr;
  vec_rsc_0_4_d <= vec_rsc_0_4_i_d;
  vec_rsc_0_4_wadr <= vec_rsc_0_4_i_wadr;
  vec_rsc_0_4_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_4_i_q_d <= vec_rsc_0_4_i_q_d_1;
  vec_rsc_0_4_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_4_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_5_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_5_i_q,
      radr => vec_rsc_0_5_i_radr,
      we => vec_rsc_0_5_we,
      d => vec_rsc_0_5_i_d,
      wadr => vec_rsc_0_5_i_wadr,
      d_d => vec_rsc_0_5_i_d_d,
      q_d => vec_rsc_0_5_i_q_d_1,
      radr_d => vec_rsc_0_5_i_radr_d,
      wadr_d => vec_rsc_0_5_i_wadr_d,
      we_d => vec_rsc_0_5_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_5_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_5_i_q <= vec_rsc_0_5_q;
  vec_rsc_0_5_radr <= vec_rsc_0_5_i_radr;
  vec_rsc_0_5_d <= vec_rsc_0_5_i_d;
  vec_rsc_0_5_wadr <= vec_rsc_0_5_i_wadr;
  vec_rsc_0_5_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_5_i_q_d <= vec_rsc_0_5_i_q_d_1;
  vec_rsc_0_5_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_5_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_6_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_6_i_q,
      radr => vec_rsc_0_6_i_radr,
      we => vec_rsc_0_6_we,
      d => vec_rsc_0_6_i_d,
      wadr => vec_rsc_0_6_i_wadr,
      d_d => vec_rsc_0_6_i_d_d,
      q_d => vec_rsc_0_6_i_q_d_1,
      radr_d => vec_rsc_0_6_i_radr_d,
      wadr_d => vec_rsc_0_6_i_wadr_d,
      we_d => vec_rsc_0_6_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_6_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_6_i_q <= vec_rsc_0_6_q;
  vec_rsc_0_6_radr <= vec_rsc_0_6_i_radr;
  vec_rsc_0_6_d <= vec_rsc_0_6_i_d;
  vec_rsc_0_6_wadr <= vec_rsc_0_6_i_wadr;
  vec_rsc_0_6_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_6_i_q_d <= vec_rsc_0_6_i_q_d_1;
  vec_rsc_0_6_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_6_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_7_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_7_i_q,
      radr => vec_rsc_0_7_i_radr,
      we => vec_rsc_0_7_we,
      d => vec_rsc_0_7_i_d,
      wadr => vec_rsc_0_7_i_wadr,
      d_d => vec_rsc_0_7_i_d_d,
      q_d => vec_rsc_0_7_i_q_d_1,
      radr_d => vec_rsc_0_7_i_radr_d,
      wadr_d => vec_rsc_0_7_i_wadr_d,
      we_d => vec_rsc_0_7_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_7_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_7_i_q <= vec_rsc_0_7_q;
  vec_rsc_0_7_radr <= vec_rsc_0_7_i_radr;
  vec_rsc_0_7_d <= vec_rsc_0_7_i_d;
  vec_rsc_0_7_wadr <= vec_rsc_0_7_i_wadr;
  vec_rsc_0_7_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_7_i_q_d <= vec_rsc_0_7_i_q_d_1;
  vec_rsc_0_7_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_7_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_8_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_8_i_q,
      radr => vec_rsc_0_8_i_radr,
      we => vec_rsc_0_8_we,
      d => vec_rsc_0_8_i_d,
      wadr => vec_rsc_0_8_i_wadr,
      d_d => vec_rsc_0_8_i_d_d,
      q_d => vec_rsc_0_8_i_q_d_1,
      radr_d => vec_rsc_0_8_i_radr_d,
      wadr_d => vec_rsc_0_8_i_wadr_d,
      we_d => vec_rsc_0_8_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_8_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_8_i_q <= vec_rsc_0_8_q;
  vec_rsc_0_8_radr <= vec_rsc_0_8_i_radr;
  vec_rsc_0_8_d <= vec_rsc_0_8_i_d;
  vec_rsc_0_8_wadr <= vec_rsc_0_8_i_wadr;
  vec_rsc_0_8_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_8_i_q_d <= vec_rsc_0_8_i_q_d_1;
  vec_rsc_0_8_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_8_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_9_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_9_i_q,
      radr => vec_rsc_0_9_i_radr,
      we => vec_rsc_0_9_we,
      d => vec_rsc_0_9_i_d,
      wadr => vec_rsc_0_9_i_wadr,
      d_d => vec_rsc_0_9_i_d_d,
      q_d => vec_rsc_0_9_i_q_d_1,
      radr_d => vec_rsc_0_9_i_radr_d,
      wadr_d => vec_rsc_0_9_i_wadr_d,
      we_d => vec_rsc_0_9_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_9_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_9_i_q <= vec_rsc_0_9_q;
  vec_rsc_0_9_radr <= vec_rsc_0_9_i_radr;
  vec_rsc_0_9_d <= vec_rsc_0_9_i_d;
  vec_rsc_0_9_wadr <= vec_rsc_0_9_i_wadr;
  vec_rsc_0_9_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_9_i_q_d <= vec_rsc_0_9_i_q_d_1;
  vec_rsc_0_9_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_9_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_10_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_10_i_q,
      radr => vec_rsc_0_10_i_radr,
      we => vec_rsc_0_10_we,
      d => vec_rsc_0_10_i_d,
      wadr => vec_rsc_0_10_i_wadr,
      d_d => vec_rsc_0_10_i_d_d,
      q_d => vec_rsc_0_10_i_q_d_1,
      radr_d => vec_rsc_0_10_i_radr_d,
      wadr_d => vec_rsc_0_10_i_wadr_d,
      we_d => vec_rsc_0_10_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_10_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_10_i_q <= vec_rsc_0_10_q;
  vec_rsc_0_10_radr <= vec_rsc_0_10_i_radr;
  vec_rsc_0_10_d <= vec_rsc_0_10_i_d;
  vec_rsc_0_10_wadr <= vec_rsc_0_10_i_wadr;
  vec_rsc_0_10_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_10_i_q_d <= vec_rsc_0_10_i_q_d_1;
  vec_rsc_0_10_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_10_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_11_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_11_i_q,
      radr => vec_rsc_0_11_i_radr,
      we => vec_rsc_0_11_we,
      d => vec_rsc_0_11_i_d,
      wadr => vec_rsc_0_11_i_wadr,
      d_d => vec_rsc_0_11_i_d_d,
      q_d => vec_rsc_0_11_i_q_d_1,
      radr_d => vec_rsc_0_11_i_radr_d,
      wadr_d => vec_rsc_0_11_i_wadr_d,
      we_d => vec_rsc_0_11_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_11_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_11_i_q <= vec_rsc_0_11_q;
  vec_rsc_0_11_radr <= vec_rsc_0_11_i_radr;
  vec_rsc_0_11_d <= vec_rsc_0_11_i_d;
  vec_rsc_0_11_wadr <= vec_rsc_0_11_i_wadr;
  vec_rsc_0_11_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_11_i_q_d <= vec_rsc_0_11_i_q_d_1;
  vec_rsc_0_11_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_11_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_12_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_12_i_q,
      radr => vec_rsc_0_12_i_radr,
      we => vec_rsc_0_12_we,
      d => vec_rsc_0_12_i_d,
      wadr => vec_rsc_0_12_i_wadr,
      d_d => vec_rsc_0_12_i_d_d,
      q_d => vec_rsc_0_12_i_q_d_1,
      radr_d => vec_rsc_0_12_i_radr_d,
      wadr_d => vec_rsc_0_12_i_wadr_d,
      we_d => vec_rsc_0_12_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_12_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_12_i_q <= vec_rsc_0_12_q;
  vec_rsc_0_12_radr <= vec_rsc_0_12_i_radr;
  vec_rsc_0_12_d <= vec_rsc_0_12_i_d;
  vec_rsc_0_12_wadr <= vec_rsc_0_12_i_wadr;
  vec_rsc_0_12_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_12_i_q_d <= vec_rsc_0_12_i_q_d_1;
  vec_rsc_0_12_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_12_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_13_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_13_i_q,
      radr => vec_rsc_0_13_i_radr,
      we => vec_rsc_0_13_we,
      d => vec_rsc_0_13_i_d,
      wadr => vec_rsc_0_13_i_wadr,
      d_d => vec_rsc_0_13_i_d_d,
      q_d => vec_rsc_0_13_i_q_d_1,
      radr_d => vec_rsc_0_13_i_radr_d,
      wadr_d => vec_rsc_0_13_i_wadr_d,
      we_d => vec_rsc_0_13_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_13_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_13_i_q <= vec_rsc_0_13_q;
  vec_rsc_0_13_radr <= vec_rsc_0_13_i_radr;
  vec_rsc_0_13_d <= vec_rsc_0_13_i_d;
  vec_rsc_0_13_wadr <= vec_rsc_0_13_i_wadr;
  vec_rsc_0_13_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_13_i_q_d <= vec_rsc_0_13_i_q_d_1;
  vec_rsc_0_13_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_13_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_14_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_14_i_q,
      radr => vec_rsc_0_14_i_radr,
      we => vec_rsc_0_14_we,
      d => vec_rsc_0_14_i_d,
      wadr => vec_rsc_0_14_i_wadr,
      d_d => vec_rsc_0_14_i_d_d,
      q_d => vec_rsc_0_14_i_q_d_1,
      radr_d => vec_rsc_0_14_i_radr_d,
      wadr_d => vec_rsc_0_14_i_wadr_d,
      we_d => vec_rsc_0_14_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_14_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_14_i_q <= vec_rsc_0_14_q;
  vec_rsc_0_14_radr <= vec_rsc_0_14_i_radr;
  vec_rsc_0_14_d <= vec_rsc_0_14_i_d;
  vec_rsc_0_14_wadr <= vec_rsc_0_14_i_wadr;
  vec_rsc_0_14_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_14_i_q_d <= vec_rsc_0_14_i_q_d_1;
  vec_rsc_0_14_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_14_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  vec_rsc_0_15_i : inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_6_64_64_64_64_1_gen
    PORT MAP(
      q => vec_rsc_0_15_i_q,
      radr => vec_rsc_0_15_i_radr,
      we => vec_rsc_0_15_we,
      d => vec_rsc_0_15_i_d,
      wadr => vec_rsc_0_15_i_wadr,
      d_d => vec_rsc_0_15_i_d_d,
      q_d => vec_rsc_0_15_i_q_d_1,
      radr_d => vec_rsc_0_15_i_radr_d,
      wadr_d => vec_rsc_0_15_i_wadr_d,
      we_d => vec_rsc_0_15_i_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => vec_rsc_0_15_i_we_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d
    );
  vec_rsc_0_15_i_q <= vec_rsc_0_15_q;
  vec_rsc_0_15_radr <= vec_rsc_0_15_i_radr;
  vec_rsc_0_15_d <= vec_rsc_0_15_i_d;
  vec_rsc_0_15_wadr <= vec_rsc_0_15_i_wadr;
  vec_rsc_0_15_i_d_d <= vec_rsc_0_0_i_d_d_iff;
  vec_rsc_0_15_i_q_d <= vec_rsc_0_15_i_q_d_1;
  vec_rsc_0_15_i_radr_d <= vec_rsc_0_0_i_radr_d_iff;
  vec_rsc_0_15_i_wadr_d <= vec_rsc_0_0_i_wadr_d_iff;

  inPlaceNTT_DIT_core_inst : inPlaceNTT_DIT_core
    PORT MAP(
      clk => clk,
      rst => rst,
      vec_rsc_triosy_0_0_lz => vec_rsc_triosy_0_0_lz,
      vec_rsc_triosy_0_1_lz => vec_rsc_triosy_0_1_lz,
      vec_rsc_triosy_0_2_lz => vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz => vec_rsc_triosy_0_3_lz,
      vec_rsc_triosy_0_4_lz => vec_rsc_triosy_0_4_lz,
      vec_rsc_triosy_0_5_lz => vec_rsc_triosy_0_5_lz,
      vec_rsc_triosy_0_6_lz => vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz => vec_rsc_triosy_0_7_lz,
      vec_rsc_triosy_0_8_lz => vec_rsc_triosy_0_8_lz,
      vec_rsc_triosy_0_9_lz => vec_rsc_triosy_0_9_lz,
      vec_rsc_triosy_0_10_lz => vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz => vec_rsc_triosy_0_11_lz,
      vec_rsc_triosy_0_12_lz => vec_rsc_triosy_0_12_lz,
      vec_rsc_triosy_0_13_lz => vec_rsc_triosy_0_13_lz,
      vec_rsc_triosy_0_14_lz => vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz => vec_rsc_triosy_0_15_lz,
      p_rsc_dat => inPlaceNTT_DIT_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_dat => inPlaceNTT_DIT_core_inst_r_rsc_dat,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      vec_rsc_0_0_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_q_d,
      vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_q_d,
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_2_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_q_d,
      vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_q_d,
      vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_4_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_q_d,
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_5_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_q_d,
      vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_q_d,
      vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_7_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_q_d,
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_8_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_q_d,
      vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_q_d,
      vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_10_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_q_d,
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_11_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_q_d,
      vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_q_d,
      vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_13_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_q_d,
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_14_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_q_d,
      vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_q_d => inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_q_d,
      vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d => vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_0_i_d_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_d_d_pff,
      vec_rsc_0_0_i_radr_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_radr_d_pff,
      vec_rsc_0_0_i_wadr_d_pff => inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_wadr_d_pff,
      vec_rsc_0_0_i_we_d_pff => vec_rsc_0_0_i_we_d_iff,
      vec_rsc_0_1_i_we_d_pff => vec_rsc_0_1_i_we_d_iff,
      vec_rsc_0_2_i_we_d_pff => vec_rsc_0_2_i_we_d_iff,
      vec_rsc_0_3_i_we_d_pff => vec_rsc_0_3_i_we_d_iff,
      vec_rsc_0_4_i_we_d_pff => vec_rsc_0_4_i_we_d_iff,
      vec_rsc_0_5_i_we_d_pff => vec_rsc_0_5_i_we_d_iff,
      vec_rsc_0_6_i_we_d_pff => vec_rsc_0_6_i_we_d_iff,
      vec_rsc_0_7_i_we_d_pff => vec_rsc_0_7_i_we_d_iff,
      vec_rsc_0_8_i_we_d_pff => vec_rsc_0_8_i_we_d_iff,
      vec_rsc_0_9_i_we_d_pff => vec_rsc_0_9_i_we_d_iff,
      vec_rsc_0_10_i_we_d_pff => vec_rsc_0_10_i_we_d_iff,
      vec_rsc_0_11_i_we_d_pff => vec_rsc_0_11_i_we_d_iff,
      vec_rsc_0_12_i_we_d_pff => vec_rsc_0_12_i_we_d_iff,
      vec_rsc_0_13_i_we_d_pff => vec_rsc_0_13_i_we_d_iff,
      vec_rsc_0_14_i_we_d_pff => vec_rsc_0_14_i_we_d_iff,
      vec_rsc_0_15_i_we_d_pff => vec_rsc_0_15_i_we_d_iff
    );
  inPlaceNTT_DIT_core_inst_p_rsc_dat <= p_rsc_dat;
  inPlaceNTT_DIT_core_inst_r_rsc_dat <= r_rsc_dat;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_q_d <= vec_rsc_0_0_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_1_i_q_d <= vec_rsc_0_1_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_2_i_q_d <= vec_rsc_0_2_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_3_i_q_d <= vec_rsc_0_3_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_4_i_q_d <= vec_rsc_0_4_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_5_i_q_d <= vec_rsc_0_5_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_6_i_q_d <= vec_rsc_0_6_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_7_i_q_d <= vec_rsc_0_7_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_8_i_q_d <= vec_rsc_0_8_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_9_i_q_d <= vec_rsc_0_9_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_10_i_q_d <= vec_rsc_0_10_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_11_i_q_d <= vec_rsc_0_11_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_12_i_q_d <= vec_rsc_0_12_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_13_i_q_d <= vec_rsc_0_13_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_14_i_q_d <= vec_rsc_0_14_i_q_d;
  inPlaceNTT_DIT_core_inst_vec_rsc_0_15_i_q_d <= vec_rsc_0_15_i_q_d;
  vec_rsc_0_0_i_d_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_d_d_pff;
  vec_rsc_0_0_i_radr_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_radr_d_pff;
  vec_rsc_0_0_i_wadr_d_iff <= inPlaceNTT_DIT_core_inst_vec_rsc_0_0_i_wadr_d_pff;

END v11;



