
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Mon May 17 21:44:25 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_11_64_2048_2048_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_11_64_2048_2048_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [10:0] adra;
  input [10:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_11_64_2048_2048_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_11_64_2048_2048_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [10:0] adra;
  input [10:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_10_tr0, modExp_while_C_47_tr0, VEC_LOOP_1_COMP_LOOP_C_1_tr0,
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_47_tr0, VEC_LOOP_1_COMP_LOOP_C_76_tr0,
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47_tr0, VEC_LOOP_1_COMP_LOOP_C_152_tr0,
      VEC_LOOP_C_0_tr0, VEC_LOOP_2_COMP_LOOP_C_1_tr0, VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_47_tr0,
      VEC_LOOP_2_COMP_LOOP_C_76_tr0, VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47_tr0,
      VEC_LOOP_2_COMP_LOOP_C_152_tr0, VEC_LOOP_C_1_tr0, STAGE_LOOP_C_11_tr0
);
  input clk;
  input rst;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;
  input STAGE_LOOP_C_10_tr0;
  input modExp_while_C_47_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_1_tr0;
  input VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_47_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_76_tr0;
  input VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_152_tr0;
  input VEC_LOOP_C_0_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_1_tr0;
  input VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_47_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_76_tr0;
  input VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_152_tr0;
  input VEC_LOOP_C_1_tr0;
  input STAGE_LOOP_C_11_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 10'd0,
    STAGE_LOOP_C_0 = 10'd1,
    STAGE_LOOP_C_1 = 10'd2,
    STAGE_LOOP_C_2 = 10'd3,
    STAGE_LOOP_C_3 = 10'd4,
    STAGE_LOOP_C_4 = 10'd5,
    STAGE_LOOP_C_5 = 10'd6,
    STAGE_LOOP_C_6 = 10'd7,
    STAGE_LOOP_C_7 = 10'd8,
    STAGE_LOOP_C_8 = 10'd9,
    STAGE_LOOP_C_9 = 10'd10,
    STAGE_LOOP_C_10 = 10'd11,
    modExp_while_C_0 = 10'd12,
    modExp_while_C_1 = 10'd13,
    modExp_while_C_2 = 10'd14,
    modExp_while_C_3 = 10'd15,
    modExp_while_C_4 = 10'd16,
    modExp_while_C_5 = 10'd17,
    modExp_while_C_6 = 10'd18,
    modExp_while_C_7 = 10'd19,
    modExp_while_C_8 = 10'd20,
    modExp_while_C_9 = 10'd21,
    modExp_while_C_10 = 10'd22,
    modExp_while_C_11 = 10'd23,
    modExp_while_C_12 = 10'd24,
    modExp_while_C_13 = 10'd25,
    modExp_while_C_14 = 10'd26,
    modExp_while_C_15 = 10'd27,
    modExp_while_C_16 = 10'd28,
    modExp_while_C_17 = 10'd29,
    modExp_while_C_18 = 10'd30,
    modExp_while_C_19 = 10'd31,
    modExp_while_C_20 = 10'd32,
    modExp_while_C_21 = 10'd33,
    modExp_while_C_22 = 10'd34,
    modExp_while_C_23 = 10'd35,
    modExp_while_C_24 = 10'd36,
    modExp_while_C_25 = 10'd37,
    modExp_while_C_26 = 10'd38,
    modExp_while_C_27 = 10'd39,
    modExp_while_C_28 = 10'd40,
    modExp_while_C_29 = 10'd41,
    modExp_while_C_30 = 10'd42,
    modExp_while_C_31 = 10'd43,
    modExp_while_C_32 = 10'd44,
    modExp_while_C_33 = 10'd45,
    modExp_while_C_34 = 10'd46,
    modExp_while_C_35 = 10'd47,
    modExp_while_C_36 = 10'd48,
    modExp_while_C_37 = 10'd49,
    modExp_while_C_38 = 10'd50,
    modExp_while_C_39 = 10'd51,
    modExp_while_C_40 = 10'd52,
    modExp_while_C_41 = 10'd53,
    modExp_while_C_42 = 10'd54,
    modExp_while_C_43 = 10'd55,
    modExp_while_C_44 = 10'd56,
    modExp_while_C_45 = 10'd57,
    modExp_while_C_46 = 10'd58,
    modExp_while_C_47 = 10'd59,
    VEC_LOOP_1_COMP_LOOP_C_0 = 10'd60,
    VEC_LOOP_1_COMP_LOOP_C_1 = 10'd61,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0 = 10'd62,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1 = 10'd63,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2 = 10'd64,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3 = 10'd65,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4 = 10'd66,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5 = 10'd67,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6 = 10'd68,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7 = 10'd69,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8 = 10'd70,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9 = 10'd71,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10 = 10'd72,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11 = 10'd73,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12 = 10'd74,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13 = 10'd75,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14 = 10'd76,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15 = 10'd77,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16 = 10'd78,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17 = 10'd79,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18 = 10'd80,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19 = 10'd81,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20 = 10'd82,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21 = 10'd83,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22 = 10'd84,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23 = 10'd85,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24 = 10'd86,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_25 = 10'd87,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_26 = 10'd88,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_27 = 10'd89,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_28 = 10'd90,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_29 = 10'd91,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_30 = 10'd92,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_31 = 10'd93,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_32 = 10'd94,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_33 = 10'd95,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_34 = 10'd96,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_35 = 10'd97,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_36 = 10'd98,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_37 = 10'd99,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38 = 10'd100,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_39 = 10'd101,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_40 = 10'd102,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_41 = 10'd103,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_42 = 10'd104,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_43 = 10'd105,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_44 = 10'd106,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_45 = 10'd107,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_46 = 10'd108,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_47 = 10'd109,
    VEC_LOOP_1_COMP_LOOP_C_2 = 10'd110,
    VEC_LOOP_1_COMP_LOOP_C_3 = 10'd111,
    VEC_LOOP_1_COMP_LOOP_C_4 = 10'd112,
    VEC_LOOP_1_COMP_LOOP_C_5 = 10'd113,
    VEC_LOOP_1_COMP_LOOP_C_6 = 10'd114,
    VEC_LOOP_1_COMP_LOOP_C_7 = 10'd115,
    VEC_LOOP_1_COMP_LOOP_C_8 = 10'd116,
    VEC_LOOP_1_COMP_LOOP_C_9 = 10'd117,
    VEC_LOOP_1_COMP_LOOP_C_10 = 10'd118,
    VEC_LOOP_1_COMP_LOOP_C_11 = 10'd119,
    VEC_LOOP_1_COMP_LOOP_C_12 = 10'd120,
    VEC_LOOP_1_COMP_LOOP_C_13 = 10'd121,
    VEC_LOOP_1_COMP_LOOP_C_14 = 10'd122,
    VEC_LOOP_1_COMP_LOOP_C_15 = 10'd123,
    VEC_LOOP_1_COMP_LOOP_C_16 = 10'd124,
    VEC_LOOP_1_COMP_LOOP_C_17 = 10'd125,
    VEC_LOOP_1_COMP_LOOP_C_18 = 10'd126,
    VEC_LOOP_1_COMP_LOOP_C_19 = 10'd127,
    VEC_LOOP_1_COMP_LOOP_C_20 = 10'd128,
    VEC_LOOP_1_COMP_LOOP_C_21 = 10'd129,
    VEC_LOOP_1_COMP_LOOP_C_22 = 10'd130,
    VEC_LOOP_1_COMP_LOOP_C_23 = 10'd131,
    VEC_LOOP_1_COMP_LOOP_C_24 = 10'd132,
    VEC_LOOP_1_COMP_LOOP_C_25 = 10'd133,
    VEC_LOOP_1_COMP_LOOP_C_26 = 10'd134,
    VEC_LOOP_1_COMP_LOOP_C_27 = 10'd135,
    VEC_LOOP_1_COMP_LOOP_C_28 = 10'd136,
    VEC_LOOP_1_COMP_LOOP_C_29 = 10'd137,
    VEC_LOOP_1_COMP_LOOP_C_30 = 10'd138,
    VEC_LOOP_1_COMP_LOOP_C_31 = 10'd139,
    VEC_LOOP_1_COMP_LOOP_C_32 = 10'd140,
    VEC_LOOP_1_COMP_LOOP_C_33 = 10'd141,
    VEC_LOOP_1_COMP_LOOP_C_34 = 10'd142,
    VEC_LOOP_1_COMP_LOOP_C_35 = 10'd143,
    VEC_LOOP_1_COMP_LOOP_C_36 = 10'd144,
    VEC_LOOP_1_COMP_LOOP_C_37 = 10'd145,
    VEC_LOOP_1_COMP_LOOP_C_38 = 10'd146,
    VEC_LOOP_1_COMP_LOOP_C_39 = 10'd147,
    VEC_LOOP_1_COMP_LOOP_C_40 = 10'd148,
    VEC_LOOP_1_COMP_LOOP_C_41 = 10'd149,
    VEC_LOOP_1_COMP_LOOP_C_42 = 10'd150,
    VEC_LOOP_1_COMP_LOOP_C_43 = 10'd151,
    VEC_LOOP_1_COMP_LOOP_C_44 = 10'd152,
    VEC_LOOP_1_COMP_LOOP_C_45 = 10'd153,
    VEC_LOOP_1_COMP_LOOP_C_46 = 10'd154,
    VEC_LOOP_1_COMP_LOOP_C_47 = 10'd155,
    VEC_LOOP_1_COMP_LOOP_C_48 = 10'd156,
    VEC_LOOP_1_COMP_LOOP_C_49 = 10'd157,
    VEC_LOOP_1_COMP_LOOP_C_50 = 10'd158,
    VEC_LOOP_1_COMP_LOOP_C_51 = 10'd159,
    VEC_LOOP_1_COMP_LOOP_C_52 = 10'd160,
    VEC_LOOP_1_COMP_LOOP_C_53 = 10'd161,
    VEC_LOOP_1_COMP_LOOP_C_54 = 10'd162,
    VEC_LOOP_1_COMP_LOOP_C_55 = 10'd163,
    VEC_LOOP_1_COMP_LOOP_C_56 = 10'd164,
    VEC_LOOP_1_COMP_LOOP_C_57 = 10'd165,
    VEC_LOOP_1_COMP_LOOP_C_58 = 10'd166,
    VEC_LOOP_1_COMP_LOOP_C_59 = 10'd167,
    VEC_LOOP_1_COMP_LOOP_C_60 = 10'd168,
    VEC_LOOP_1_COMP_LOOP_C_61 = 10'd169,
    VEC_LOOP_1_COMP_LOOP_C_62 = 10'd170,
    VEC_LOOP_1_COMP_LOOP_C_63 = 10'd171,
    VEC_LOOP_1_COMP_LOOP_C_64 = 10'd172,
    VEC_LOOP_1_COMP_LOOP_C_65 = 10'd173,
    VEC_LOOP_1_COMP_LOOP_C_66 = 10'd174,
    VEC_LOOP_1_COMP_LOOP_C_67 = 10'd175,
    VEC_LOOP_1_COMP_LOOP_C_68 = 10'd176,
    VEC_LOOP_1_COMP_LOOP_C_69 = 10'd177,
    VEC_LOOP_1_COMP_LOOP_C_70 = 10'd178,
    VEC_LOOP_1_COMP_LOOP_C_71 = 10'd179,
    VEC_LOOP_1_COMP_LOOP_C_72 = 10'd180,
    VEC_LOOP_1_COMP_LOOP_C_73 = 10'd181,
    VEC_LOOP_1_COMP_LOOP_C_74 = 10'd182,
    VEC_LOOP_1_COMP_LOOP_C_75 = 10'd183,
    VEC_LOOP_1_COMP_LOOP_C_76 = 10'd184,
    VEC_LOOP_1_COMP_LOOP_C_77 = 10'd185,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0 = 10'd186,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1 = 10'd187,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2 = 10'd188,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3 = 10'd189,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4 = 10'd190,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5 = 10'd191,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6 = 10'd192,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7 = 10'd193,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8 = 10'd194,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9 = 10'd195,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10 = 10'd196,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11 = 10'd197,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12 = 10'd198,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13 = 10'd199,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14 = 10'd200,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15 = 10'd201,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16 = 10'd202,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17 = 10'd203,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18 = 10'd204,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19 = 10'd205,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20 = 10'd206,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21 = 10'd207,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22 = 10'd208,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23 = 10'd209,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24 = 10'd210,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_25 = 10'd211,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_26 = 10'd212,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_27 = 10'd213,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_28 = 10'd214,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_29 = 10'd215,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_30 = 10'd216,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_31 = 10'd217,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_32 = 10'd218,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_33 = 10'd219,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_34 = 10'd220,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_35 = 10'd221,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_36 = 10'd222,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_37 = 10'd223,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38 = 10'd224,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_39 = 10'd225,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_40 = 10'd226,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_41 = 10'd227,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_42 = 10'd228,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_43 = 10'd229,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_44 = 10'd230,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_45 = 10'd231,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_46 = 10'd232,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47 = 10'd233,
    VEC_LOOP_1_COMP_LOOP_C_78 = 10'd234,
    VEC_LOOP_1_COMP_LOOP_C_79 = 10'd235,
    VEC_LOOP_1_COMP_LOOP_C_80 = 10'd236,
    VEC_LOOP_1_COMP_LOOP_C_81 = 10'd237,
    VEC_LOOP_1_COMP_LOOP_C_82 = 10'd238,
    VEC_LOOP_1_COMP_LOOP_C_83 = 10'd239,
    VEC_LOOP_1_COMP_LOOP_C_84 = 10'd240,
    VEC_LOOP_1_COMP_LOOP_C_85 = 10'd241,
    VEC_LOOP_1_COMP_LOOP_C_86 = 10'd242,
    VEC_LOOP_1_COMP_LOOP_C_87 = 10'd243,
    VEC_LOOP_1_COMP_LOOP_C_88 = 10'd244,
    VEC_LOOP_1_COMP_LOOP_C_89 = 10'd245,
    VEC_LOOP_1_COMP_LOOP_C_90 = 10'd246,
    VEC_LOOP_1_COMP_LOOP_C_91 = 10'd247,
    VEC_LOOP_1_COMP_LOOP_C_92 = 10'd248,
    VEC_LOOP_1_COMP_LOOP_C_93 = 10'd249,
    VEC_LOOP_1_COMP_LOOP_C_94 = 10'd250,
    VEC_LOOP_1_COMP_LOOP_C_95 = 10'd251,
    VEC_LOOP_1_COMP_LOOP_C_96 = 10'd252,
    VEC_LOOP_1_COMP_LOOP_C_97 = 10'd253,
    VEC_LOOP_1_COMP_LOOP_C_98 = 10'd254,
    VEC_LOOP_1_COMP_LOOP_C_99 = 10'd255,
    VEC_LOOP_1_COMP_LOOP_C_100 = 10'd256,
    VEC_LOOP_1_COMP_LOOP_C_101 = 10'd257,
    VEC_LOOP_1_COMP_LOOP_C_102 = 10'd258,
    VEC_LOOP_1_COMP_LOOP_C_103 = 10'd259,
    VEC_LOOP_1_COMP_LOOP_C_104 = 10'd260,
    VEC_LOOP_1_COMP_LOOP_C_105 = 10'd261,
    VEC_LOOP_1_COMP_LOOP_C_106 = 10'd262,
    VEC_LOOP_1_COMP_LOOP_C_107 = 10'd263,
    VEC_LOOP_1_COMP_LOOP_C_108 = 10'd264,
    VEC_LOOP_1_COMP_LOOP_C_109 = 10'd265,
    VEC_LOOP_1_COMP_LOOP_C_110 = 10'd266,
    VEC_LOOP_1_COMP_LOOP_C_111 = 10'd267,
    VEC_LOOP_1_COMP_LOOP_C_112 = 10'd268,
    VEC_LOOP_1_COMP_LOOP_C_113 = 10'd269,
    VEC_LOOP_1_COMP_LOOP_C_114 = 10'd270,
    VEC_LOOP_1_COMP_LOOP_C_115 = 10'd271,
    VEC_LOOP_1_COMP_LOOP_C_116 = 10'd272,
    VEC_LOOP_1_COMP_LOOP_C_117 = 10'd273,
    VEC_LOOP_1_COMP_LOOP_C_118 = 10'd274,
    VEC_LOOP_1_COMP_LOOP_C_119 = 10'd275,
    VEC_LOOP_1_COMP_LOOP_C_120 = 10'd276,
    VEC_LOOP_1_COMP_LOOP_C_121 = 10'd277,
    VEC_LOOP_1_COMP_LOOP_C_122 = 10'd278,
    VEC_LOOP_1_COMP_LOOP_C_123 = 10'd279,
    VEC_LOOP_1_COMP_LOOP_C_124 = 10'd280,
    VEC_LOOP_1_COMP_LOOP_C_125 = 10'd281,
    VEC_LOOP_1_COMP_LOOP_C_126 = 10'd282,
    VEC_LOOP_1_COMP_LOOP_C_127 = 10'd283,
    VEC_LOOP_1_COMP_LOOP_C_128 = 10'd284,
    VEC_LOOP_1_COMP_LOOP_C_129 = 10'd285,
    VEC_LOOP_1_COMP_LOOP_C_130 = 10'd286,
    VEC_LOOP_1_COMP_LOOP_C_131 = 10'd287,
    VEC_LOOP_1_COMP_LOOP_C_132 = 10'd288,
    VEC_LOOP_1_COMP_LOOP_C_133 = 10'd289,
    VEC_LOOP_1_COMP_LOOP_C_134 = 10'd290,
    VEC_LOOP_1_COMP_LOOP_C_135 = 10'd291,
    VEC_LOOP_1_COMP_LOOP_C_136 = 10'd292,
    VEC_LOOP_1_COMP_LOOP_C_137 = 10'd293,
    VEC_LOOP_1_COMP_LOOP_C_138 = 10'd294,
    VEC_LOOP_1_COMP_LOOP_C_139 = 10'd295,
    VEC_LOOP_1_COMP_LOOP_C_140 = 10'd296,
    VEC_LOOP_1_COMP_LOOP_C_141 = 10'd297,
    VEC_LOOP_1_COMP_LOOP_C_142 = 10'd298,
    VEC_LOOP_1_COMP_LOOP_C_143 = 10'd299,
    VEC_LOOP_1_COMP_LOOP_C_144 = 10'd300,
    VEC_LOOP_1_COMP_LOOP_C_145 = 10'd301,
    VEC_LOOP_1_COMP_LOOP_C_146 = 10'd302,
    VEC_LOOP_1_COMP_LOOP_C_147 = 10'd303,
    VEC_LOOP_1_COMP_LOOP_C_148 = 10'd304,
    VEC_LOOP_1_COMP_LOOP_C_149 = 10'd305,
    VEC_LOOP_1_COMP_LOOP_C_150 = 10'd306,
    VEC_LOOP_1_COMP_LOOP_C_151 = 10'd307,
    VEC_LOOP_1_COMP_LOOP_C_152 = 10'd308,
    VEC_LOOP_C_0 = 10'd309,
    VEC_LOOP_2_COMP_LOOP_C_0 = 10'd310,
    VEC_LOOP_2_COMP_LOOP_C_1 = 10'd311,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0 = 10'd312,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1 = 10'd313,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2 = 10'd314,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3 = 10'd315,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4 = 10'd316,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5 = 10'd317,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6 = 10'd318,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7 = 10'd319,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8 = 10'd320,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9 = 10'd321,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10 = 10'd322,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11 = 10'd323,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12 = 10'd324,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13 = 10'd325,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14 = 10'd326,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15 = 10'd327,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16 = 10'd328,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17 = 10'd329,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18 = 10'd330,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19 = 10'd331,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20 = 10'd332,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21 = 10'd333,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22 = 10'd334,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23 = 10'd335,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24 = 10'd336,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_25 = 10'd337,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_26 = 10'd338,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_27 = 10'd339,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_28 = 10'd340,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_29 = 10'd341,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_30 = 10'd342,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_31 = 10'd343,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_32 = 10'd344,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_33 = 10'd345,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_34 = 10'd346,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_35 = 10'd347,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_36 = 10'd348,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_37 = 10'd349,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38 = 10'd350,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_39 = 10'd351,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_40 = 10'd352,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_41 = 10'd353,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_42 = 10'd354,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_43 = 10'd355,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_44 = 10'd356,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_45 = 10'd357,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_46 = 10'd358,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_47 = 10'd359,
    VEC_LOOP_2_COMP_LOOP_C_2 = 10'd360,
    VEC_LOOP_2_COMP_LOOP_C_3 = 10'd361,
    VEC_LOOP_2_COMP_LOOP_C_4 = 10'd362,
    VEC_LOOP_2_COMP_LOOP_C_5 = 10'd363,
    VEC_LOOP_2_COMP_LOOP_C_6 = 10'd364,
    VEC_LOOP_2_COMP_LOOP_C_7 = 10'd365,
    VEC_LOOP_2_COMP_LOOP_C_8 = 10'd366,
    VEC_LOOP_2_COMP_LOOP_C_9 = 10'd367,
    VEC_LOOP_2_COMP_LOOP_C_10 = 10'd368,
    VEC_LOOP_2_COMP_LOOP_C_11 = 10'd369,
    VEC_LOOP_2_COMP_LOOP_C_12 = 10'd370,
    VEC_LOOP_2_COMP_LOOP_C_13 = 10'd371,
    VEC_LOOP_2_COMP_LOOP_C_14 = 10'd372,
    VEC_LOOP_2_COMP_LOOP_C_15 = 10'd373,
    VEC_LOOP_2_COMP_LOOP_C_16 = 10'd374,
    VEC_LOOP_2_COMP_LOOP_C_17 = 10'd375,
    VEC_LOOP_2_COMP_LOOP_C_18 = 10'd376,
    VEC_LOOP_2_COMP_LOOP_C_19 = 10'd377,
    VEC_LOOP_2_COMP_LOOP_C_20 = 10'd378,
    VEC_LOOP_2_COMP_LOOP_C_21 = 10'd379,
    VEC_LOOP_2_COMP_LOOP_C_22 = 10'd380,
    VEC_LOOP_2_COMP_LOOP_C_23 = 10'd381,
    VEC_LOOP_2_COMP_LOOP_C_24 = 10'd382,
    VEC_LOOP_2_COMP_LOOP_C_25 = 10'd383,
    VEC_LOOP_2_COMP_LOOP_C_26 = 10'd384,
    VEC_LOOP_2_COMP_LOOP_C_27 = 10'd385,
    VEC_LOOP_2_COMP_LOOP_C_28 = 10'd386,
    VEC_LOOP_2_COMP_LOOP_C_29 = 10'd387,
    VEC_LOOP_2_COMP_LOOP_C_30 = 10'd388,
    VEC_LOOP_2_COMP_LOOP_C_31 = 10'd389,
    VEC_LOOP_2_COMP_LOOP_C_32 = 10'd390,
    VEC_LOOP_2_COMP_LOOP_C_33 = 10'd391,
    VEC_LOOP_2_COMP_LOOP_C_34 = 10'd392,
    VEC_LOOP_2_COMP_LOOP_C_35 = 10'd393,
    VEC_LOOP_2_COMP_LOOP_C_36 = 10'd394,
    VEC_LOOP_2_COMP_LOOP_C_37 = 10'd395,
    VEC_LOOP_2_COMP_LOOP_C_38 = 10'd396,
    VEC_LOOP_2_COMP_LOOP_C_39 = 10'd397,
    VEC_LOOP_2_COMP_LOOP_C_40 = 10'd398,
    VEC_LOOP_2_COMP_LOOP_C_41 = 10'd399,
    VEC_LOOP_2_COMP_LOOP_C_42 = 10'd400,
    VEC_LOOP_2_COMP_LOOP_C_43 = 10'd401,
    VEC_LOOP_2_COMP_LOOP_C_44 = 10'd402,
    VEC_LOOP_2_COMP_LOOP_C_45 = 10'd403,
    VEC_LOOP_2_COMP_LOOP_C_46 = 10'd404,
    VEC_LOOP_2_COMP_LOOP_C_47 = 10'd405,
    VEC_LOOP_2_COMP_LOOP_C_48 = 10'd406,
    VEC_LOOP_2_COMP_LOOP_C_49 = 10'd407,
    VEC_LOOP_2_COMP_LOOP_C_50 = 10'd408,
    VEC_LOOP_2_COMP_LOOP_C_51 = 10'd409,
    VEC_LOOP_2_COMP_LOOP_C_52 = 10'd410,
    VEC_LOOP_2_COMP_LOOP_C_53 = 10'd411,
    VEC_LOOP_2_COMP_LOOP_C_54 = 10'd412,
    VEC_LOOP_2_COMP_LOOP_C_55 = 10'd413,
    VEC_LOOP_2_COMP_LOOP_C_56 = 10'd414,
    VEC_LOOP_2_COMP_LOOP_C_57 = 10'd415,
    VEC_LOOP_2_COMP_LOOP_C_58 = 10'd416,
    VEC_LOOP_2_COMP_LOOP_C_59 = 10'd417,
    VEC_LOOP_2_COMP_LOOP_C_60 = 10'd418,
    VEC_LOOP_2_COMP_LOOP_C_61 = 10'd419,
    VEC_LOOP_2_COMP_LOOP_C_62 = 10'd420,
    VEC_LOOP_2_COMP_LOOP_C_63 = 10'd421,
    VEC_LOOP_2_COMP_LOOP_C_64 = 10'd422,
    VEC_LOOP_2_COMP_LOOP_C_65 = 10'd423,
    VEC_LOOP_2_COMP_LOOP_C_66 = 10'd424,
    VEC_LOOP_2_COMP_LOOP_C_67 = 10'd425,
    VEC_LOOP_2_COMP_LOOP_C_68 = 10'd426,
    VEC_LOOP_2_COMP_LOOP_C_69 = 10'd427,
    VEC_LOOP_2_COMP_LOOP_C_70 = 10'd428,
    VEC_LOOP_2_COMP_LOOP_C_71 = 10'd429,
    VEC_LOOP_2_COMP_LOOP_C_72 = 10'd430,
    VEC_LOOP_2_COMP_LOOP_C_73 = 10'd431,
    VEC_LOOP_2_COMP_LOOP_C_74 = 10'd432,
    VEC_LOOP_2_COMP_LOOP_C_75 = 10'd433,
    VEC_LOOP_2_COMP_LOOP_C_76 = 10'd434,
    VEC_LOOP_2_COMP_LOOP_C_77 = 10'd435,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0 = 10'd436,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1 = 10'd437,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2 = 10'd438,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3 = 10'd439,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4 = 10'd440,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5 = 10'd441,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6 = 10'd442,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7 = 10'd443,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8 = 10'd444,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9 = 10'd445,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10 = 10'd446,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11 = 10'd447,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12 = 10'd448,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13 = 10'd449,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14 = 10'd450,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15 = 10'd451,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16 = 10'd452,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17 = 10'd453,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18 = 10'd454,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19 = 10'd455,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20 = 10'd456,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21 = 10'd457,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22 = 10'd458,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23 = 10'd459,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24 = 10'd460,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_25 = 10'd461,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_26 = 10'd462,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_27 = 10'd463,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_28 = 10'd464,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_29 = 10'd465,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_30 = 10'd466,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_31 = 10'd467,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_32 = 10'd468,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_33 = 10'd469,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_34 = 10'd470,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_35 = 10'd471,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_36 = 10'd472,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_37 = 10'd473,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38 = 10'd474,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_39 = 10'd475,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_40 = 10'd476,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_41 = 10'd477,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_42 = 10'd478,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_43 = 10'd479,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_44 = 10'd480,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_45 = 10'd481,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_46 = 10'd482,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47 = 10'd483,
    VEC_LOOP_2_COMP_LOOP_C_78 = 10'd484,
    VEC_LOOP_2_COMP_LOOP_C_79 = 10'd485,
    VEC_LOOP_2_COMP_LOOP_C_80 = 10'd486,
    VEC_LOOP_2_COMP_LOOP_C_81 = 10'd487,
    VEC_LOOP_2_COMP_LOOP_C_82 = 10'd488,
    VEC_LOOP_2_COMP_LOOP_C_83 = 10'd489,
    VEC_LOOP_2_COMP_LOOP_C_84 = 10'd490,
    VEC_LOOP_2_COMP_LOOP_C_85 = 10'd491,
    VEC_LOOP_2_COMP_LOOP_C_86 = 10'd492,
    VEC_LOOP_2_COMP_LOOP_C_87 = 10'd493,
    VEC_LOOP_2_COMP_LOOP_C_88 = 10'd494,
    VEC_LOOP_2_COMP_LOOP_C_89 = 10'd495,
    VEC_LOOP_2_COMP_LOOP_C_90 = 10'd496,
    VEC_LOOP_2_COMP_LOOP_C_91 = 10'd497,
    VEC_LOOP_2_COMP_LOOP_C_92 = 10'd498,
    VEC_LOOP_2_COMP_LOOP_C_93 = 10'd499,
    VEC_LOOP_2_COMP_LOOP_C_94 = 10'd500,
    VEC_LOOP_2_COMP_LOOP_C_95 = 10'd501,
    VEC_LOOP_2_COMP_LOOP_C_96 = 10'd502,
    VEC_LOOP_2_COMP_LOOP_C_97 = 10'd503,
    VEC_LOOP_2_COMP_LOOP_C_98 = 10'd504,
    VEC_LOOP_2_COMP_LOOP_C_99 = 10'd505,
    VEC_LOOP_2_COMP_LOOP_C_100 = 10'd506,
    VEC_LOOP_2_COMP_LOOP_C_101 = 10'd507,
    VEC_LOOP_2_COMP_LOOP_C_102 = 10'd508,
    VEC_LOOP_2_COMP_LOOP_C_103 = 10'd509,
    VEC_LOOP_2_COMP_LOOP_C_104 = 10'd510,
    VEC_LOOP_2_COMP_LOOP_C_105 = 10'd511,
    VEC_LOOP_2_COMP_LOOP_C_106 = 10'd512,
    VEC_LOOP_2_COMP_LOOP_C_107 = 10'd513,
    VEC_LOOP_2_COMP_LOOP_C_108 = 10'd514,
    VEC_LOOP_2_COMP_LOOP_C_109 = 10'd515,
    VEC_LOOP_2_COMP_LOOP_C_110 = 10'd516,
    VEC_LOOP_2_COMP_LOOP_C_111 = 10'd517,
    VEC_LOOP_2_COMP_LOOP_C_112 = 10'd518,
    VEC_LOOP_2_COMP_LOOP_C_113 = 10'd519,
    VEC_LOOP_2_COMP_LOOP_C_114 = 10'd520,
    VEC_LOOP_2_COMP_LOOP_C_115 = 10'd521,
    VEC_LOOP_2_COMP_LOOP_C_116 = 10'd522,
    VEC_LOOP_2_COMP_LOOP_C_117 = 10'd523,
    VEC_LOOP_2_COMP_LOOP_C_118 = 10'd524,
    VEC_LOOP_2_COMP_LOOP_C_119 = 10'd525,
    VEC_LOOP_2_COMP_LOOP_C_120 = 10'd526,
    VEC_LOOP_2_COMP_LOOP_C_121 = 10'd527,
    VEC_LOOP_2_COMP_LOOP_C_122 = 10'd528,
    VEC_LOOP_2_COMP_LOOP_C_123 = 10'd529,
    VEC_LOOP_2_COMP_LOOP_C_124 = 10'd530,
    VEC_LOOP_2_COMP_LOOP_C_125 = 10'd531,
    VEC_LOOP_2_COMP_LOOP_C_126 = 10'd532,
    VEC_LOOP_2_COMP_LOOP_C_127 = 10'd533,
    VEC_LOOP_2_COMP_LOOP_C_128 = 10'd534,
    VEC_LOOP_2_COMP_LOOP_C_129 = 10'd535,
    VEC_LOOP_2_COMP_LOOP_C_130 = 10'd536,
    VEC_LOOP_2_COMP_LOOP_C_131 = 10'd537,
    VEC_LOOP_2_COMP_LOOP_C_132 = 10'd538,
    VEC_LOOP_2_COMP_LOOP_C_133 = 10'd539,
    VEC_LOOP_2_COMP_LOOP_C_134 = 10'd540,
    VEC_LOOP_2_COMP_LOOP_C_135 = 10'd541,
    VEC_LOOP_2_COMP_LOOP_C_136 = 10'd542,
    VEC_LOOP_2_COMP_LOOP_C_137 = 10'd543,
    VEC_LOOP_2_COMP_LOOP_C_138 = 10'd544,
    VEC_LOOP_2_COMP_LOOP_C_139 = 10'd545,
    VEC_LOOP_2_COMP_LOOP_C_140 = 10'd546,
    VEC_LOOP_2_COMP_LOOP_C_141 = 10'd547,
    VEC_LOOP_2_COMP_LOOP_C_142 = 10'd548,
    VEC_LOOP_2_COMP_LOOP_C_143 = 10'd549,
    VEC_LOOP_2_COMP_LOOP_C_144 = 10'd550,
    VEC_LOOP_2_COMP_LOOP_C_145 = 10'd551,
    VEC_LOOP_2_COMP_LOOP_C_146 = 10'd552,
    VEC_LOOP_2_COMP_LOOP_C_147 = 10'd553,
    VEC_LOOP_2_COMP_LOOP_C_148 = 10'd554,
    VEC_LOOP_2_COMP_LOOP_C_149 = 10'd555,
    VEC_LOOP_2_COMP_LOOP_C_150 = 10'd556,
    VEC_LOOP_2_COMP_LOOP_C_151 = 10'd557,
    VEC_LOOP_2_COMP_LOOP_C_152 = 10'd558,
    VEC_LOOP_C_1 = 10'd559,
    STAGE_LOOP_C_11 = 10'd560,
    main_C_1 = 10'd561;

  reg [9:0] state_var;
  reg [9:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 10'b0000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 10'b0000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 10'b0000000100;
        state_var_NS = STAGE_LOOP_C_4;
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 10'b0000000101;
        state_var_NS = STAGE_LOOP_C_5;
      end
      STAGE_LOOP_C_5 : begin
        fsm_output = 10'b0000000110;
        state_var_NS = STAGE_LOOP_C_6;
      end
      STAGE_LOOP_C_6 : begin
        fsm_output = 10'b0000000111;
        state_var_NS = STAGE_LOOP_C_7;
      end
      STAGE_LOOP_C_7 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = STAGE_LOOP_C_8;
      end
      STAGE_LOOP_C_8 : begin
        fsm_output = 10'b0000001001;
        state_var_NS = STAGE_LOOP_C_9;
      end
      STAGE_LOOP_C_9 : begin
        fsm_output = 10'b0000001010;
        state_var_NS = STAGE_LOOP_C_10;
      end
      STAGE_LOOP_C_10 : begin
        fsm_output = 10'b0000001011;
        if ( STAGE_LOOP_C_10_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      modExp_while_C_0 : begin
        fsm_output = 10'b0000001100;
        state_var_NS = modExp_while_C_1;
      end
      modExp_while_C_1 : begin
        fsm_output = 10'b0000001101;
        state_var_NS = modExp_while_C_2;
      end
      modExp_while_C_2 : begin
        fsm_output = 10'b0000001110;
        state_var_NS = modExp_while_C_3;
      end
      modExp_while_C_3 : begin
        fsm_output = 10'b0000001111;
        state_var_NS = modExp_while_C_4;
      end
      modExp_while_C_4 : begin
        fsm_output = 10'b0000010000;
        state_var_NS = modExp_while_C_5;
      end
      modExp_while_C_5 : begin
        fsm_output = 10'b0000010001;
        state_var_NS = modExp_while_C_6;
      end
      modExp_while_C_6 : begin
        fsm_output = 10'b0000010010;
        state_var_NS = modExp_while_C_7;
      end
      modExp_while_C_7 : begin
        fsm_output = 10'b0000010011;
        state_var_NS = modExp_while_C_8;
      end
      modExp_while_C_8 : begin
        fsm_output = 10'b0000010100;
        state_var_NS = modExp_while_C_9;
      end
      modExp_while_C_9 : begin
        fsm_output = 10'b0000010101;
        state_var_NS = modExp_while_C_10;
      end
      modExp_while_C_10 : begin
        fsm_output = 10'b0000010110;
        state_var_NS = modExp_while_C_11;
      end
      modExp_while_C_11 : begin
        fsm_output = 10'b0000010111;
        state_var_NS = modExp_while_C_12;
      end
      modExp_while_C_12 : begin
        fsm_output = 10'b0000011000;
        state_var_NS = modExp_while_C_13;
      end
      modExp_while_C_13 : begin
        fsm_output = 10'b0000011001;
        state_var_NS = modExp_while_C_14;
      end
      modExp_while_C_14 : begin
        fsm_output = 10'b0000011010;
        state_var_NS = modExp_while_C_15;
      end
      modExp_while_C_15 : begin
        fsm_output = 10'b0000011011;
        state_var_NS = modExp_while_C_16;
      end
      modExp_while_C_16 : begin
        fsm_output = 10'b0000011100;
        state_var_NS = modExp_while_C_17;
      end
      modExp_while_C_17 : begin
        fsm_output = 10'b0000011101;
        state_var_NS = modExp_while_C_18;
      end
      modExp_while_C_18 : begin
        fsm_output = 10'b0000011110;
        state_var_NS = modExp_while_C_19;
      end
      modExp_while_C_19 : begin
        fsm_output = 10'b0000011111;
        state_var_NS = modExp_while_C_20;
      end
      modExp_while_C_20 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = modExp_while_C_21;
      end
      modExp_while_C_21 : begin
        fsm_output = 10'b0000100001;
        state_var_NS = modExp_while_C_22;
      end
      modExp_while_C_22 : begin
        fsm_output = 10'b0000100010;
        state_var_NS = modExp_while_C_23;
      end
      modExp_while_C_23 : begin
        fsm_output = 10'b0000100011;
        state_var_NS = modExp_while_C_24;
      end
      modExp_while_C_24 : begin
        fsm_output = 10'b0000100100;
        state_var_NS = modExp_while_C_25;
      end
      modExp_while_C_25 : begin
        fsm_output = 10'b0000100101;
        state_var_NS = modExp_while_C_26;
      end
      modExp_while_C_26 : begin
        fsm_output = 10'b0000100110;
        state_var_NS = modExp_while_C_27;
      end
      modExp_while_C_27 : begin
        fsm_output = 10'b0000100111;
        state_var_NS = modExp_while_C_28;
      end
      modExp_while_C_28 : begin
        fsm_output = 10'b0000101000;
        state_var_NS = modExp_while_C_29;
      end
      modExp_while_C_29 : begin
        fsm_output = 10'b0000101001;
        state_var_NS = modExp_while_C_30;
      end
      modExp_while_C_30 : begin
        fsm_output = 10'b0000101010;
        state_var_NS = modExp_while_C_31;
      end
      modExp_while_C_31 : begin
        fsm_output = 10'b0000101011;
        state_var_NS = modExp_while_C_32;
      end
      modExp_while_C_32 : begin
        fsm_output = 10'b0000101100;
        state_var_NS = modExp_while_C_33;
      end
      modExp_while_C_33 : begin
        fsm_output = 10'b0000101101;
        state_var_NS = modExp_while_C_34;
      end
      modExp_while_C_34 : begin
        fsm_output = 10'b0000101110;
        state_var_NS = modExp_while_C_35;
      end
      modExp_while_C_35 : begin
        fsm_output = 10'b0000101111;
        state_var_NS = modExp_while_C_36;
      end
      modExp_while_C_36 : begin
        fsm_output = 10'b0000110000;
        state_var_NS = modExp_while_C_37;
      end
      modExp_while_C_37 : begin
        fsm_output = 10'b0000110001;
        state_var_NS = modExp_while_C_38;
      end
      modExp_while_C_38 : begin
        fsm_output = 10'b0000110010;
        state_var_NS = modExp_while_C_39;
      end
      modExp_while_C_39 : begin
        fsm_output = 10'b0000110011;
        state_var_NS = modExp_while_C_40;
      end
      modExp_while_C_40 : begin
        fsm_output = 10'b0000110100;
        state_var_NS = modExp_while_C_41;
      end
      modExp_while_C_41 : begin
        fsm_output = 10'b0000110101;
        state_var_NS = modExp_while_C_42;
      end
      modExp_while_C_42 : begin
        fsm_output = 10'b0000110110;
        state_var_NS = modExp_while_C_43;
      end
      modExp_while_C_43 : begin
        fsm_output = 10'b0000110111;
        state_var_NS = modExp_while_C_44;
      end
      modExp_while_C_44 : begin
        fsm_output = 10'b0000111000;
        state_var_NS = modExp_while_C_45;
      end
      modExp_while_C_45 : begin
        fsm_output = 10'b0000111001;
        state_var_NS = modExp_while_C_46;
      end
      modExp_while_C_46 : begin
        fsm_output = 10'b0000111010;
        state_var_NS = modExp_while_C_47;
      end
      modExp_while_C_47 : begin
        fsm_output = 10'b0000111011;
        if ( modExp_while_C_47_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_0 : begin
        fsm_output = 10'b0000111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_C_1 : begin
        fsm_output = 10'b0000111101;
        if ( VEC_LOOP_1_COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 10'b0000111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 10'b0000111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 10'b0001000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 10'b0001000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 10'b0001000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 10'b0001000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 10'b0001000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 10'b0001000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 10'b0001000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 10'b0001001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 10'b0001001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 10'b0001001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 10'b0001001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 10'b0001001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 10'b0001001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 10'b0001001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 10'b0001001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 10'b0001010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 10'b0001010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 10'b0001010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 10'b0001010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 10'b0001010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 10'b0001010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 10'b0001010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_25;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 10'b0001010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_26;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 10'b0001011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_27;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 10'b0001011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_28;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 10'b0001011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_29;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 10'b0001011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_30;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 10'b0001011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_31;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 10'b0001011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_32;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 10'b0001011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_33;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 10'b0001011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_34;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 10'b0001100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_35;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 10'b0001100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_36;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 10'b0001100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_37;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 10'b0001100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 10'b0001100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_39;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_39 : begin
        fsm_output = 10'b0001100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_40;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_40 : begin
        fsm_output = 10'b0001100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_41;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_41 : begin
        fsm_output = 10'b0001100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_42;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_42 : begin
        fsm_output = 10'b0001101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_43;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_43 : begin
        fsm_output = 10'b0001101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_44;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_44 : begin
        fsm_output = 10'b0001101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_45;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_45 : begin
        fsm_output = 10'b0001101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_46;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_46 : begin
        fsm_output = 10'b0001101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_47;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_47 : begin
        fsm_output = 10'b0001101101;
        if ( VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_47_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_2 : begin
        fsm_output = 10'b0001101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_C_3 : begin
        fsm_output = 10'b0001101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_C_4 : begin
        fsm_output = 10'b0001110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_C_5 : begin
        fsm_output = 10'b0001110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_C_6 : begin
        fsm_output = 10'b0001110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_C_7 : begin
        fsm_output = 10'b0001110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_C_8 : begin
        fsm_output = 10'b0001110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_C_9 : begin
        fsm_output = 10'b0001110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_C_10 : begin
        fsm_output = 10'b0001110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_C_11 : begin
        fsm_output = 10'b0001110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_C_12 : begin
        fsm_output = 10'b0001111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_C_13 : begin
        fsm_output = 10'b0001111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_C_14 : begin
        fsm_output = 10'b0001111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_C_15 : begin
        fsm_output = 10'b0001111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_C_16 : begin
        fsm_output = 10'b0001111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_C_17 : begin
        fsm_output = 10'b0001111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_C_18 : begin
        fsm_output = 10'b0001111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_C_19 : begin
        fsm_output = 10'b0001111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_C_20 : begin
        fsm_output = 10'b0010000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_C_21 : begin
        fsm_output = 10'b0010000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_C_22 : begin
        fsm_output = 10'b0010000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_C_23 : begin
        fsm_output = 10'b0010000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_C_24 : begin
        fsm_output = 10'b0010000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_25;
      end
      VEC_LOOP_1_COMP_LOOP_C_25 : begin
        fsm_output = 10'b0010000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_26;
      end
      VEC_LOOP_1_COMP_LOOP_C_26 : begin
        fsm_output = 10'b0010000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_27;
      end
      VEC_LOOP_1_COMP_LOOP_C_27 : begin
        fsm_output = 10'b0010000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_28;
      end
      VEC_LOOP_1_COMP_LOOP_C_28 : begin
        fsm_output = 10'b0010001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_29;
      end
      VEC_LOOP_1_COMP_LOOP_C_29 : begin
        fsm_output = 10'b0010001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_30;
      end
      VEC_LOOP_1_COMP_LOOP_C_30 : begin
        fsm_output = 10'b0010001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_31;
      end
      VEC_LOOP_1_COMP_LOOP_C_31 : begin
        fsm_output = 10'b0010001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_32;
      end
      VEC_LOOP_1_COMP_LOOP_C_32 : begin
        fsm_output = 10'b0010001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_33;
      end
      VEC_LOOP_1_COMP_LOOP_C_33 : begin
        fsm_output = 10'b0010001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_34;
      end
      VEC_LOOP_1_COMP_LOOP_C_34 : begin
        fsm_output = 10'b0010001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_35;
      end
      VEC_LOOP_1_COMP_LOOP_C_35 : begin
        fsm_output = 10'b0010001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_36;
      end
      VEC_LOOP_1_COMP_LOOP_C_36 : begin
        fsm_output = 10'b0010010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_37;
      end
      VEC_LOOP_1_COMP_LOOP_C_37 : begin
        fsm_output = 10'b0010010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_38;
      end
      VEC_LOOP_1_COMP_LOOP_C_38 : begin
        fsm_output = 10'b0010010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_39;
      end
      VEC_LOOP_1_COMP_LOOP_C_39 : begin
        fsm_output = 10'b0010010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_40;
      end
      VEC_LOOP_1_COMP_LOOP_C_40 : begin
        fsm_output = 10'b0010010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_41;
      end
      VEC_LOOP_1_COMP_LOOP_C_41 : begin
        fsm_output = 10'b0010010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_42;
      end
      VEC_LOOP_1_COMP_LOOP_C_42 : begin
        fsm_output = 10'b0010010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_43;
      end
      VEC_LOOP_1_COMP_LOOP_C_43 : begin
        fsm_output = 10'b0010010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_44;
      end
      VEC_LOOP_1_COMP_LOOP_C_44 : begin
        fsm_output = 10'b0010011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_45;
      end
      VEC_LOOP_1_COMP_LOOP_C_45 : begin
        fsm_output = 10'b0010011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_46;
      end
      VEC_LOOP_1_COMP_LOOP_C_46 : begin
        fsm_output = 10'b0010011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_47;
      end
      VEC_LOOP_1_COMP_LOOP_C_47 : begin
        fsm_output = 10'b0010011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_48;
      end
      VEC_LOOP_1_COMP_LOOP_C_48 : begin
        fsm_output = 10'b0010011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_49;
      end
      VEC_LOOP_1_COMP_LOOP_C_49 : begin
        fsm_output = 10'b0010011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_50;
      end
      VEC_LOOP_1_COMP_LOOP_C_50 : begin
        fsm_output = 10'b0010011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_51;
      end
      VEC_LOOP_1_COMP_LOOP_C_51 : begin
        fsm_output = 10'b0010011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_52;
      end
      VEC_LOOP_1_COMP_LOOP_C_52 : begin
        fsm_output = 10'b0010100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_53;
      end
      VEC_LOOP_1_COMP_LOOP_C_53 : begin
        fsm_output = 10'b0010100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_54;
      end
      VEC_LOOP_1_COMP_LOOP_C_54 : begin
        fsm_output = 10'b0010100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_55;
      end
      VEC_LOOP_1_COMP_LOOP_C_55 : begin
        fsm_output = 10'b0010100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_56;
      end
      VEC_LOOP_1_COMP_LOOP_C_56 : begin
        fsm_output = 10'b0010100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_57;
      end
      VEC_LOOP_1_COMP_LOOP_C_57 : begin
        fsm_output = 10'b0010100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_58;
      end
      VEC_LOOP_1_COMP_LOOP_C_58 : begin
        fsm_output = 10'b0010100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_59;
      end
      VEC_LOOP_1_COMP_LOOP_C_59 : begin
        fsm_output = 10'b0010100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_60;
      end
      VEC_LOOP_1_COMP_LOOP_C_60 : begin
        fsm_output = 10'b0010101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_61;
      end
      VEC_LOOP_1_COMP_LOOP_C_61 : begin
        fsm_output = 10'b0010101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_62;
      end
      VEC_LOOP_1_COMP_LOOP_C_62 : begin
        fsm_output = 10'b0010101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_63;
      end
      VEC_LOOP_1_COMP_LOOP_C_63 : begin
        fsm_output = 10'b0010101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_64;
      end
      VEC_LOOP_1_COMP_LOOP_C_64 : begin
        fsm_output = 10'b0010101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_65;
      end
      VEC_LOOP_1_COMP_LOOP_C_65 : begin
        fsm_output = 10'b0010101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_66;
      end
      VEC_LOOP_1_COMP_LOOP_C_66 : begin
        fsm_output = 10'b0010101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_67;
      end
      VEC_LOOP_1_COMP_LOOP_C_67 : begin
        fsm_output = 10'b0010101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_68;
      end
      VEC_LOOP_1_COMP_LOOP_C_68 : begin
        fsm_output = 10'b0010110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_69;
      end
      VEC_LOOP_1_COMP_LOOP_C_69 : begin
        fsm_output = 10'b0010110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_70;
      end
      VEC_LOOP_1_COMP_LOOP_C_70 : begin
        fsm_output = 10'b0010110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_71;
      end
      VEC_LOOP_1_COMP_LOOP_C_71 : begin
        fsm_output = 10'b0010110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_72;
      end
      VEC_LOOP_1_COMP_LOOP_C_72 : begin
        fsm_output = 10'b0010110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_73;
      end
      VEC_LOOP_1_COMP_LOOP_C_73 : begin
        fsm_output = 10'b0010110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_74;
      end
      VEC_LOOP_1_COMP_LOOP_C_74 : begin
        fsm_output = 10'b0010110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_75;
      end
      VEC_LOOP_1_COMP_LOOP_C_75 : begin
        fsm_output = 10'b0010110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_76;
      end
      VEC_LOOP_1_COMP_LOOP_C_76 : begin
        fsm_output = 10'b0010111000;
        if ( VEC_LOOP_1_COMP_LOOP_C_76_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_77;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_77 : begin
        fsm_output = 10'b0010111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 10'b0010111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 10'b0010111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 10'b0010111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 10'b0010111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 10'b0010111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 10'b0010111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 10'b0011000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 10'b0011000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 10'b0011000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 10'b0011000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 10'b0011000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 10'b0011000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 10'b0011000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 10'b0011000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 10'b0011001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 10'b0011001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 10'b0011001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 10'b0011001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 10'b0011001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 10'b0011001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 10'b0011001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 10'b0011001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 10'b0011010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 10'b0011010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 10'b0011010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_25;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 10'b0011010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_26;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 10'b0011010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_27;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 10'b0011010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_28;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 10'b0011010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_29;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 10'b0011010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_30;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 10'b0011011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_31;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 10'b0011011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_32;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 10'b0011011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_33;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 10'b0011011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_34;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 10'b0011011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_35;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 10'b0011011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_36;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 10'b0011011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_37;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 10'b0011011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 10'b0011100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_39;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_39 : begin
        fsm_output = 10'b0011100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_40;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_40 : begin
        fsm_output = 10'b0011100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_41;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_41 : begin
        fsm_output = 10'b0011100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_42;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_42 : begin
        fsm_output = 10'b0011100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_43;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_43 : begin
        fsm_output = 10'b0011100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_44;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_44 : begin
        fsm_output = 10'b0011100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_45;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_45 : begin
        fsm_output = 10'b0011100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_46;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_46 : begin
        fsm_output = 10'b0011101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47 : begin
        fsm_output = 10'b0011101001;
        if ( VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_78;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_78 : begin
        fsm_output = 10'b0011101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_79;
      end
      VEC_LOOP_1_COMP_LOOP_C_79 : begin
        fsm_output = 10'b0011101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_80;
      end
      VEC_LOOP_1_COMP_LOOP_C_80 : begin
        fsm_output = 10'b0011101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_81;
      end
      VEC_LOOP_1_COMP_LOOP_C_81 : begin
        fsm_output = 10'b0011101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_82;
      end
      VEC_LOOP_1_COMP_LOOP_C_82 : begin
        fsm_output = 10'b0011101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_83;
      end
      VEC_LOOP_1_COMP_LOOP_C_83 : begin
        fsm_output = 10'b0011101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_84;
      end
      VEC_LOOP_1_COMP_LOOP_C_84 : begin
        fsm_output = 10'b0011110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_85;
      end
      VEC_LOOP_1_COMP_LOOP_C_85 : begin
        fsm_output = 10'b0011110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_86;
      end
      VEC_LOOP_1_COMP_LOOP_C_86 : begin
        fsm_output = 10'b0011110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_87;
      end
      VEC_LOOP_1_COMP_LOOP_C_87 : begin
        fsm_output = 10'b0011110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_88;
      end
      VEC_LOOP_1_COMP_LOOP_C_88 : begin
        fsm_output = 10'b0011110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_89;
      end
      VEC_LOOP_1_COMP_LOOP_C_89 : begin
        fsm_output = 10'b0011110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_90;
      end
      VEC_LOOP_1_COMP_LOOP_C_90 : begin
        fsm_output = 10'b0011110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_91;
      end
      VEC_LOOP_1_COMP_LOOP_C_91 : begin
        fsm_output = 10'b0011110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_92;
      end
      VEC_LOOP_1_COMP_LOOP_C_92 : begin
        fsm_output = 10'b0011111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_93;
      end
      VEC_LOOP_1_COMP_LOOP_C_93 : begin
        fsm_output = 10'b0011111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_94;
      end
      VEC_LOOP_1_COMP_LOOP_C_94 : begin
        fsm_output = 10'b0011111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_95;
      end
      VEC_LOOP_1_COMP_LOOP_C_95 : begin
        fsm_output = 10'b0011111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_96;
      end
      VEC_LOOP_1_COMP_LOOP_C_96 : begin
        fsm_output = 10'b0011111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_97;
      end
      VEC_LOOP_1_COMP_LOOP_C_97 : begin
        fsm_output = 10'b0011111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_98;
      end
      VEC_LOOP_1_COMP_LOOP_C_98 : begin
        fsm_output = 10'b0011111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_99;
      end
      VEC_LOOP_1_COMP_LOOP_C_99 : begin
        fsm_output = 10'b0011111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_100;
      end
      VEC_LOOP_1_COMP_LOOP_C_100 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_101;
      end
      VEC_LOOP_1_COMP_LOOP_C_101 : begin
        fsm_output = 10'b0100000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_102;
      end
      VEC_LOOP_1_COMP_LOOP_C_102 : begin
        fsm_output = 10'b0100000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_103;
      end
      VEC_LOOP_1_COMP_LOOP_C_103 : begin
        fsm_output = 10'b0100000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_104;
      end
      VEC_LOOP_1_COMP_LOOP_C_104 : begin
        fsm_output = 10'b0100000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_105;
      end
      VEC_LOOP_1_COMP_LOOP_C_105 : begin
        fsm_output = 10'b0100000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_106;
      end
      VEC_LOOP_1_COMP_LOOP_C_106 : begin
        fsm_output = 10'b0100000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_107;
      end
      VEC_LOOP_1_COMP_LOOP_C_107 : begin
        fsm_output = 10'b0100000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_108;
      end
      VEC_LOOP_1_COMP_LOOP_C_108 : begin
        fsm_output = 10'b0100001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_109;
      end
      VEC_LOOP_1_COMP_LOOP_C_109 : begin
        fsm_output = 10'b0100001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_110;
      end
      VEC_LOOP_1_COMP_LOOP_C_110 : begin
        fsm_output = 10'b0100001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_111;
      end
      VEC_LOOP_1_COMP_LOOP_C_111 : begin
        fsm_output = 10'b0100001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_112;
      end
      VEC_LOOP_1_COMP_LOOP_C_112 : begin
        fsm_output = 10'b0100001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_113;
      end
      VEC_LOOP_1_COMP_LOOP_C_113 : begin
        fsm_output = 10'b0100001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_114;
      end
      VEC_LOOP_1_COMP_LOOP_C_114 : begin
        fsm_output = 10'b0100001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_115;
      end
      VEC_LOOP_1_COMP_LOOP_C_115 : begin
        fsm_output = 10'b0100001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_116;
      end
      VEC_LOOP_1_COMP_LOOP_C_116 : begin
        fsm_output = 10'b0100010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_117;
      end
      VEC_LOOP_1_COMP_LOOP_C_117 : begin
        fsm_output = 10'b0100010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_118;
      end
      VEC_LOOP_1_COMP_LOOP_C_118 : begin
        fsm_output = 10'b0100010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_119;
      end
      VEC_LOOP_1_COMP_LOOP_C_119 : begin
        fsm_output = 10'b0100010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_120;
      end
      VEC_LOOP_1_COMP_LOOP_C_120 : begin
        fsm_output = 10'b0100010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_121;
      end
      VEC_LOOP_1_COMP_LOOP_C_121 : begin
        fsm_output = 10'b0100010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_122;
      end
      VEC_LOOP_1_COMP_LOOP_C_122 : begin
        fsm_output = 10'b0100010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_123;
      end
      VEC_LOOP_1_COMP_LOOP_C_123 : begin
        fsm_output = 10'b0100010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_124;
      end
      VEC_LOOP_1_COMP_LOOP_C_124 : begin
        fsm_output = 10'b0100011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_125;
      end
      VEC_LOOP_1_COMP_LOOP_C_125 : begin
        fsm_output = 10'b0100011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_126;
      end
      VEC_LOOP_1_COMP_LOOP_C_126 : begin
        fsm_output = 10'b0100011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_127;
      end
      VEC_LOOP_1_COMP_LOOP_C_127 : begin
        fsm_output = 10'b0100011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_128;
      end
      VEC_LOOP_1_COMP_LOOP_C_128 : begin
        fsm_output = 10'b0100011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_129;
      end
      VEC_LOOP_1_COMP_LOOP_C_129 : begin
        fsm_output = 10'b0100011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_130;
      end
      VEC_LOOP_1_COMP_LOOP_C_130 : begin
        fsm_output = 10'b0100011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_131;
      end
      VEC_LOOP_1_COMP_LOOP_C_131 : begin
        fsm_output = 10'b0100011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_132;
      end
      VEC_LOOP_1_COMP_LOOP_C_132 : begin
        fsm_output = 10'b0100100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_133;
      end
      VEC_LOOP_1_COMP_LOOP_C_133 : begin
        fsm_output = 10'b0100100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_134;
      end
      VEC_LOOP_1_COMP_LOOP_C_134 : begin
        fsm_output = 10'b0100100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_135;
      end
      VEC_LOOP_1_COMP_LOOP_C_135 : begin
        fsm_output = 10'b0100100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_136;
      end
      VEC_LOOP_1_COMP_LOOP_C_136 : begin
        fsm_output = 10'b0100100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_137;
      end
      VEC_LOOP_1_COMP_LOOP_C_137 : begin
        fsm_output = 10'b0100100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_138;
      end
      VEC_LOOP_1_COMP_LOOP_C_138 : begin
        fsm_output = 10'b0100100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_139;
      end
      VEC_LOOP_1_COMP_LOOP_C_139 : begin
        fsm_output = 10'b0100100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_140;
      end
      VEC_LOOP_1_COMP_LOOP_C_140 : begin
        fsm_output = 10'b0100101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_141;
      end
      VEC_LOOP_1_COMP_LOOP_C_141 : begin
        fsm_output = 10'b0100101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_142;
      end
      VEC_LOOP_1_COMP_LOOP_C_142 : begin
        fsm_output = 10'b0100101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_143;
      end
      VEC_LOOP_1_COMP_LOOP_C_143 : begin
        fsm_output = 10'b0100101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_144;
      end
      VEC_LOOP_1_COMP_LOOP_C_144 : begin
        fsm_output = 10'b0100101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_145;
      end
      VEC_LOOP_1_COMP_LOOP_C_145 : begin
        fsm_output = 10'b0100101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_146;
      end
      VEC_LOOP_1_COMP_LOOP_C_146 : begin
        fsm_output = 10'b0100101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_147;
      end
      VEC_LOOP_1_COMP_LOOP_C_147 : begin
        fsm_output = 10'b0100101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_148;
      end
      VEC_LOOP_1_COMP_LOOP_C_148 : begin
        fsm_output = 10'b0100110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_149;
      end
      VEC_LOOP_1_COMP_LOOP_C_149 : begin
        fsm_output = 10'b0100110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_150;
      end
      VEC_LOOP_1_COMP_LOOP_C_150 : begin
        fsm_output = 10'b0100110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_151;
      end
      VEC_LOOP_1_COMP_LOOP_C_151 : begin
        fsm_output = 10'b0100110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_152;
      end
      VEC_LOOP_1_COMP_LOOP_C_152 : begin
        fsm_output = 10'b0100110100;
        if ( VEC_LOOP_1_COMP_LOOP_C_152_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 10'b0100110101;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_11;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_0 : begin
        fsm_output = 10'b0100110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_C_1 : begin
        fsm_output = 10'b0100110111;
        if ( VEC_LOOP_2_COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 10'b0100111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 10'b0100111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 10'b0100111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 10'b0100111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 10'b0100111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 10'b0100111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 10'b0100111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 10'b0100111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 10'b0101000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 10'b0101000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 10'b0101000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 10'b0101000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 10'b0101000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 10'b0101000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 10'b0101000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 10'b0101000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 10'b0101001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 10'b0101001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 10'b0101001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 10'b0101001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 10'b0101001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 10'b0101001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 10'b0101001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 10'b0101001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 10'b0101010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_25;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 10'b0101010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_26;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 10'b0101010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_27;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 10'b0101010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_28;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 10'b0101010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_29;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 10'b0101010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_30;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 10'b0101010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_31;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 10'b0101010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_32;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 10'b0101011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_33;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 10'b0101011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_34;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 10'b0101011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_35;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 10'b0101011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_36;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 10'b0101011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_37;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 10'b0101011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 10'b0101011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_39;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_39 : begin
        fsm_output = 10'b0101011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_40;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_40 : begin
        fsm_output = 10'b0101100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_41;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_41 : begin
        fsm_output = 10'b0101100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_42;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_42 : begin
        fsm_output = 10'b0101100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_43;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_43 : begin
        fsm_output = 10'b0101100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_44;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_44 : begin
        fsm_output = 10'b0101100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_45;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_45 : begin
        fsm_output = 10'b0101100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_46;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_46 : begin
        fsm_output = 10'b0101100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_47;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_47 : begin
        fsm_output = 10'b0101100111;
        if ( VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_47_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_2 : begin
        fsm_output = 10'b0101101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_C_3 : begin
        fsm_output = 10'b0101101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_C_4 : begin
        fsm_output = 10'b0101101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_C_5 : begin
        fsm_output = 10'b0101101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_C_6 : begin
        fsm_output = 10'b0101101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_C_7 : begin
        fsm_output = 10'b0101101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_C_8 : begin
        fsm_output = 10'b0101101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_C_9 : begin
        fsm_output = 10'b0101101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_C_10 : begin
        fsm_output = 10'b0101110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_C_11 : begin
        fsm_output = 10'b0101110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_C_12 : begin
        fsm_output = 10'b0101110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_C_13 : begin
        fsm_output = 10'b0101110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_C_14 : begin
        fsm_output = 10'b0101110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_C_15 : begin
        fsm_output = 10'b0101110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_C_16 : begin
        fsm_output = 10'b0101110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_C_17 : begin
        fsm_output = 10'b0101110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_C_18 : begin
        fsm_output = 10'b0101111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_C_19 : begin
        fsm_output = 10'b0101111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_C_20 : begin
        fsm_output = 10'b0101111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_C_21 : begin
        fsm_output = 10'b0101111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_C_22 : begin
        fsm_output = 10'b0101111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_C_23 : begin
        fsm_output = 10'b0101111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_C_24 : begin
        fsm_output = 10'b0101111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_25;
      end
      VEC_LOOP_2_COMP_LOOP_C_25 : begin
        fsm_output = 10'b0101111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_26;
      end
      VEC_LOOP_2_COMP_LOOP_C_26 : begin
        fsm_output = 10'b0110000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_27;
      end
      VEC_LOOP_2_COMP_LOOP_C_27 : begin
        fsm_output = 10'b0110000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_28;
      end
      VEC_LOOP_2_COMP_LOOP_C_28 : begin
        fsm_output = 10'b0110000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_29;
      end
      VEC_LOOP_2_COMP_LOOP_C_29 : begin
        fsm_output = 10'b0110000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_30;
      end
      VEC_LOOP_2_COMP_LOOP_C_30 : begin
        fsm_output = 10'b0110000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_31;
      end
      VEC_LOOP_2_COMP_LOOP_C_31 : begin
        fsm_output = 10'b0110000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_32;
      end
      VEC_LOOP_2_COMP_LOOP_C_32 : begin
        fsm_output = 10'b0110000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_33;
      end
      VEC_LOOP_2_COMP_LOOP_C_33 : begin
        fsm_output = 10'b0110000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_34;
      end
      VEC_LOOP_2_COMP_LOOP_C_34 : begin
        fsm_output = 10'b0110001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_35;
      end
      VEC_LOOP_2_COMP_LOOP_C_35 : begin
        fsm_output = 10'b0110001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_36;
      end
      VEC_LOOP_2_COMP_LOOP_C_36 : begin
        fsm_output = 10'b0110001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_37;
      end
      VEC_LOOP_2_COMP_LOOP_C_37 : begin
        fsm_output = 10'b0110001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_38;
      end
      VEC_LOOP_2_COMP_LOOP_C_38 : begin
        fsm_output = 10'b0110001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_39;
      end
      VEC_LOOP_2_COMP_LOOP_C_39 : begin
        fsm_output = 10'b0110001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_40;
      end
      VEC_LOOP_2_COMP_LOOP_C_40 : begin
        fsm_output = 10'b0110001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_41;
      end
      VEC_LOOP_2_COMP_LOOP_C_41 : begin
        fsm_output = 10'b0110001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_42;
      end
      VEC_LOOP_2_COMP_LOOP_C_42 : begin
        fsm_output = 10'b0110010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_43;
      end
      VEC_LOOP_2_COMP_LOOP_C_43 : begin
        fsm_output = 10'b0110010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_44;
      end
      VEC_LOOP_2_COMP_LOOP_C_44 : begin
        fsm_output = 10'b0110010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_45;
      end
      VEC_LOOP_2_COMP_LOOP_C_45 : begin
        fsm_output = 10'b0110010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_46;
      end
      VEC_LOOP_2_COMP_LOOP_C_46 : begin
        fsm_output = 10'b0110010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_47;
      end
      VEC_LOOP_2_COMP_LOOP_C_47 : begin
        fsm_output = 10'b0110010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_48;
      end
      VEC_LOOP_2_COMP_LOOP_C_48 : begin
        fsm_output = 10'b0110010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_49;
      end
      VEC_LOOP_2_COMP_LOOP_C_49 : begin
        fsm_output = 10'b0110010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_50;
      end
      VEC_LOOP_2_COMP_LOOP_C_50 : begin
        fsm_output = 10'b0110011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_51;
      end
      VEC_LOOP_2_COMP_LOOP_C_51 : begin
        fsm_output = 10'b0110011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_52;
      end
      VEC_LOOP_2_COMP_LOOP_C_52 : begin
        fsm_output = 10'b0110011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_53;
      end
      VEC_LOOP_2_COMP_LOOP_C_53 : begin
        fsm_output = 10'b0110011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_54;
      end
      VEC_LOOP_2_COMP_LOOP_C_54 : begin
        fsm_output = 10'b0110011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_55;
      end
      VEC_LOOP_2_COMP_LOOP_C_55 : begin
        fsm_output = 10'b0110011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_56;
      end
      VEC_LOOP_2_COMP_LOOP_C_56 : begin
        fsm_output = 10'b0110011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_57;
      end
      VEC_LOOP_2_COMP_LOOP_C_57 : begin
        fsm_output = 10'b0110011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_58;
      end
      VEC_LOOP_2_COMP_LOOP_C_58 : begin
        fsm_output = 10'b0110100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_59;
      end
      VEC_LOOP_2_COMP_LOOP_C_59 : begin
        fsm_output = 10'b0110100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_60;
      end
      VEC_LOOP_2_COMP_LOOP_C_60 : begin
        fsm_output = 10'b0110100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_61;
      end
      VEC_LOOP_2_COMP_LOOP_C_61 : begin
        fsm_output = 10'b0110100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_62;
      end
      VEC_LOOP_2_COMP_LOOP_C_62 : begin
        fsm_output = 10'b0110100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_63;
      end
      VEC_LOOP_2_COMP_LOOP_C_63 : begin
        fsm_output = 10'b0110100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_64;
      end
      VEC_LOOP_2_COMP_LOOP_C_64 : begin
        fsm_output = 10'b0110100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_65;
      end
      VEC_LOOP_2_COMP_LOOP_C_65 : begin
        fsm_output = 10'b0110100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_66;
      end
      VEC_LOOP_2_COMP_LOOP_C_66 : begin
        fsm_output = 10'b0110101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_67;
      end
      VEC_LOOP_2_COMP_LOOP_C_67 : begin
        fsm_output = 10'b0110101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_68;
      end
      VEC_LOOP_2_COMP_LOOP_C_68 : begin
        fsm_output = 10'b0110101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_69;
      end
      VEC_LOOP_2_COMP_LOOP_C_69 : begin
        fsm_output = 10'b0110101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_70;
      end
      VEC_LOOP_2_COMP_LOOP_C_70 : begin
        fsm_output = 10'b0110101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_71;
      end
      VEC_LOOP_2_COMP_LOOP_C_71 : begin
        fsm_output = 10'b0110101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_72;
      end
      VEC_LOOP_2_COMP_LOOP_C_72 : begin
        fsm_output = 10'b0110101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_73;
      end
      VEC_LOOP_2_COMP_LOOP_C_73 : begin
        fsm_output = 10'b0110101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_74;
      end
      VEC_LOOP_2_COMP_LOOP_C_74 : begin
        fsm_output = 10'b0110110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_75;
      end
      VEC_LOOP_2_COMP_LOOP_C_75 : begin
        fsm_output = 10'b0110110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_76;
      end
      VEC_LOOP_2_COMP_LOOP_C_76 : begin
        fsm_output = 10'b0110110010;
        if ( VEC_LOOP_2_COMP_LOOP_C_76_tr0 ) begin
          state_var_NS = VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_77;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_77 : begin
        fsm_output = 10'b0110110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 10'b0110110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 10'b0110110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 10'b0110110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 10'b0110110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 10'b0110111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 10'b0110111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 10'b0110111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 10'b0110111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 10'b0110111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 10'b0110111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 10'b0110111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 10'b0110111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 10'b0111000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 10'b0111000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 10'b0111000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 10'b0111000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 10'b0111000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 10'b0111000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 10'b0111000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 10'b0111000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 10'b0111001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 10'b0111001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 10'b0111001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 10'b0111001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 10'b0111001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_25;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 10'b0111001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_26;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 10'b0111001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_27;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 10'b0111001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_28;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 10'b0111010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_29;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 10'b0111010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_30;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 10'b0111010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_31;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 10'b0111010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_32;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 10'b0111010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_33;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 10'b0111010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_34;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 10'b0111010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_35;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 10'b0111010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_36;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 10'b0111011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_37;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 10'b0111011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 10'b0111011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_39;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_39 : begin
        fsm_output = 10'b0111011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_40;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_40 : begin
        fsm_output = 10'b0111011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_41;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_41 : begin
        fsm_output = 10'b0111011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_42;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_42 : begin
        fsm_output = 10'b0111011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_43;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_43 : begin
        fsm_output = 10'b0111011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_44;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_44 : begin
        fsm_output = 10'b0111100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_45;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_45 : begin
        fsm_output = 10'b0111100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_46;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_46 : begin
        fsm_output = 10'b0111100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47 : begin
        fsm_output = 10'b0111100011;
        if ( VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_78;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_78 : begin
        fsm_output = 10'b0111100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_79;
      end
      VEC_LOOP_2_COMP_LOOP_C_79 : begin
        fsm_output = 10'b0111100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_80;
      end
      VEC_LOOP_2_COMP_LOOP_C_80 : begin
        fsm_output = 10'b0111100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_81;
      end
      VEC_LOOP_2_COMP_LOOP_C_81 : begin
        fsm_output = 10'b0111100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_82;
      end
      VEC_LOOP_2_COMP_LOOP_C_82 : begin
        fsm_output = 10'b0111101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_83;
      end
      VEC_LOOP_2_COMP_LOOP_C_83 : begin
        fsm_output = 10'b0111101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_84;
      end
      VEC_LOOP_2_COMP_LOOP_C_84 : begin
        fsm_output = 10'b0111101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_85;
      end
      VEC_LOOP_2_COMP_LOOP_C_85 : begin
        fsm_output = 10'b0111101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_86;
      end
      VEC_LOOP_2_COMP_LOOP_C_86 : begin
        fsm_output = 10'b0111101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_87;
      end
      VEC_LOOP_2_COMP_LOOP_C_87 : begin
        fsm_output = 10'b0111101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_88;
      end
      VEC_LOOP_2_COMP_LOOP_C_88 : begin
        fsm_output = 10'b0111101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_89;
      end
      VEC_LOOP_2_COMP_LOOP_C_89 : begin
        fsm_output = 10'b0111101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_90;
      end
      VEC_LOOP_2_COMP_LOOP_C_90 : begin
        fsm_output = 10'b0111110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_91;
      end
      VEC_LOOP_2_COMP_LOOP_C_91 : begin
        fsm_output = 10'b0111110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_92;
      end
      VEC_LOOP_2_COMP_LOOP_C_92 : begin
        fsm_output = 10'b0111110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_93;
      end
      VEC_LOOP_2_COMP_LOOP_C_93 : begin
        fsm_output = 10'b0111110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_94;
      end
      VEC_LOOP_2_COMP_LOOP_C_94 : begin
        fsm_output = 10'b0111110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_95;
      end
      VEC_LOOP_2_COMP_LOOP_C_95 : begin
        fsm_output = 10'b0111110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_96;
      end
      VEC_LOOP_2_COMP_LOOP_C_96 : begin
        fsm_output = 10'b0111110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_97;
      end
      VEC_LOOP_2_COMP_LOOP_C_97 : begin
        fsm_output = 10'b0111110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_98;
      end
      VEC_LOOP_2_COMP_LOOP_C_98 : begin
        fsm_output = 10'b0111111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_99;
      end
      VEC_LOOP_2_COMP_LOOP_C_99 : begin
        fsm_output = 10'b0111111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_100;
      end
      VEC_LOOP_2_COMP_LOOP_C_100 : begin
        fsm_output = 10'b0111111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_101;
      end
      VEC_LOOP_2_COMP_LOOP_C_101 : begin
        fsm_output = 10'b0111111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_102;
      end
      VEC_LOOP_2_COMP_LOOP_C_102 : begin
        fsm_output = 10'b0111111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_103;
      end
      VEC_LOOP_2_COMP_LOOP_C_103 : begin
        fsm_output = 10'b0111111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_104;
      end
      VEC_LOOP_2_COMP_LOOP_C_104 : begin
        fsm_output = 10'b0111111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_105;
      end
      VEC_LOOP_2_COMP_LOOP_C_105 : begin
        fsm_output = 10'b0111111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_106;
      end
      VEC_LOOP_2_COMP_LOOP_C_106 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_107;
      end
      VEC_LOOP_2_COMP_LOOP_C_107 : begin
        fsm_output = 10'b1000000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_108;
      end
      VEC_LOOP_2_COMP_LOOP_C_108 : begin
        fsm_output = 10'b1000000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_109;
      end
      VEC_LOOP_2_COMP_LOOP_C_109 : begin
        fsm_output = 10'b1000000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_110;
      end
      VEC_LOOP_2_COMP_LOOP_C_110 : begin
        fsm_output = 10'b1000000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_111;
      end
      VEC_LOOP_2_COMP_LOOP_C_111 : begin
        fsm_output = 10'b1000000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_112;
      end
      VEC_LOOP_2_COMP_LOOP_C_112 : begin
        fsm_output = 10'b1000000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_113;
      end
      VEC_LOOP_2_COMP_LOOP_C_113 : begin
        fsm_output = 10'b1000000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_114;
      end
      VEC_LOOP_2_COMP_LOOP_C_114 : begin
        fsm_output = 10'b1000001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_115;
      end
      VEC_LOOP_2_COMP_LOOP_C_115 : begin
        fsm_output = 10'b1000001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_116;
      end
      VEC_LOOP_2_COMP_LOOP_C_116 : begin
        fsm_output = 10'b1000001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_117;
      end
      VEC_LOOP_2_COMP_LOOP_C_117 : begin
        fsm_output = 10'b1000001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_118;
      end
      VEC_LOOP_2_COMP_LOOP_C_118 : begin
        fsm_output = 10'b1000001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_119;
      end
      VEC_LOOP_2_COMP_LOOP_C_119 : begin
        fsm_output = 10'b1000001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_120;
      end
      VEC_LOOP_2_COMP_LOOP_C_120 : begin
        fsm_output = 10'b1000001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_121;
      end
      VEC_LOOP_2_COMP_LOOP_C_121 : begin
        fsm_output = 10'b1000001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_122;
      end
      VEC_LOOP_2_COMP_LOOP_C_122 : begin
        fsm_output = 10'b1000010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_123;
      end
      VEC_LOOP_2_COMP_LOOP_C_123 : begin
        fsm_output = 10'b1000010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_124;
      end
      VEC_LOOP_2_COMP_LOOP_C_124 : begin
        fsm_output = 10'b1000010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_125;
      end
      VEC_LOOP_2_COMP_LOOP_C_125 : begin
        fsm_output = 10'b1000010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_126;
      end
      VEC_LOOP_2_COMP_LOOP_C_126 : begin
        fsm_output = 10'b1000010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_127;
      end
      VEC_LOOP_2_COMP_LOOP_C_127 : begin
        fsm_output = 10'b1000010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_128;
      end
      VEC_LOOP_2_COMP_LOOP_C_128 : begin
        fsm_output = 10'b1000010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_129;
      end
      VEC_LOOP_2_COMP_LOOP_C_129 : begin
        fsm_output = 10'b1000010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_130;
      end
      VEC_LOOP_2_COMP_LOOP_C_130 : begin
        fsm_output = 10'b1000011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_131;
      end
      VEC_LOOP_2_COMP_LOOP_C_131 : begin
        fsm_output = 10'b1000011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_132;
      end
      VEC_LOOP_2_COMP_LOOP_C_132 : begin
        fsm_output = 10'b1000011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_133;
      end
      VEC_LOOP_2_COMP_LOOP_C_133 : begin
        fsm_output = 10'b1000011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_134;
      end
      VEC_LOOP_2_COMP_LOOP_C_134 : begin
        fsm_output = 10'b1000011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_135;
      end
      VEC_LOOP_2_COMP_LOOP_C_135 : begin
        fsm_output = 10'b1000011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_136;
      end
      VEC_LOOP_2_COMP_LOOP_C_136 : begin
        fsm_output = 10'b1000011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_137;
      end
      VEC_LOOP_2_COMP_LOOP_C_137 : begin
        fsm_output = 10'b1000011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_138;
      end
      VEC_LOOP_2_COMP_LOOP_C_138 : begin
        fsm_output = 10'b1000100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_139;
      end
      VEC_LOOP_2_COMP_LOOP_C_139 : begin
        fsm_output = 10'b1000100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_140;
      end
      VEC_LOOP_2_COMP_LOOP_C_140 : begin
        fsm_output = 10'b1000100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_141;
      end
      VEC_LOOP_2_COMP_LOOP_C_141 : begin
        fsm_output = 10'b1000100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_142;
      end
      VEC_LOOP_2_COMP_LOOP_C_142 : begin
        fsm_output = 10'b1000100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_143;
      end
      VEC_LOOP_2_COMP_LOOP_C_143 : begin
        fsm_output = 10'b1000100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_144;
      end
      VEC_LOOP_2_COMP_LOOP_C_144 : begin
        fsm_output = 10'b1000100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_145;
      end
      VEC_LOOP_2_COMP_LOOP_C_145 : begin
        fsm_output = 10'b1000100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_146;
      end
      VEC_LOOP_2_COMP_LOOP_C_146 : begin
        fsm_output = 10'b1000101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_147;
      end
      VEC_LOOP_2_COMP_LOOP_C_147 : begin
        fsm_output = 10'b1000101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_148;
      end
      VEC_LOOP_2_COMP_LOOP_C_148 : begin
        fsm_output = 10'b1000101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_149;
      end
      VEC_LOOP_2_COMP_LOOP_C_149 : begin
        fsm_output = 10'b1000101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_150;
      end
      VEC_LOOP_2_COMP_LOOP_C_150 : begin
        fsm_output = 10'b1000101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_151;
      end
      VEC_LOOP_2_COMP_LOOP_C_151 : begin
        fsm_output = 10'b1000101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_152;
      end
      VEC_LOOP_2_COMP_LOOP_C_152 : begin
        fsm_output = 10'b1000101110;
        if ( VEC_LOOP_2_COMP_LOOP_C_152_tr0 ) begin
          state_var_NS = VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_1 : begin
        fsm_output = 10'b1000101111;
        if ( VEC_LOOP_C_1_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_11;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_11 : begin
        fsm_output = 10'b1000110000;
        if ( STAGE_LOOP_C_11_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 10'b1000110001;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 10'b0000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_wait_dp
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_wait_dp (
  clk, operator_66_true_div_cmp_z, operator_66_true_div_cmp_z_oreg
);
  input clk;
  input [64:0] operator_66_true_div_cmp_z;
  output [63:0] operator_66_true_div_cmp_z_oreg;


  // Interconnect Declarations
  reg [63:0] operator_66_true_div_cmp_z_oreg_pconst_63_0;


  // Interconnect Declarations for Component Instantiations 
  assign operator_66_true_div_cmp_z_oreg = operator_66_true_div_cmp_z_oreg_pconst_63_0;
  always @(posedge clk) begin
    operator_66_true_div_cmp_z_oreg_pconst_63_0 <= operator_66_true_div_cmp_z[63:0];
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, p_rsc_dat, p_rsc_triosy_lz,
      r_rsc_dat, r_rsc_triosy_lz, vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_1_i_qa_d, vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, operator_66_true_div_cmp_a,
      operator_66_true_div_cmp_b, operator_66_true_div_cmp_z, vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff, vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [64:0] operator_66_true_div_cmp_a;
  reg [64:0] operator_66_true_div_cmp_a;
  output [10:0] operator_66_true_div_cmp_b;
  input [64:0] operator_66_true_div_cmp_z;
  output [10:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  reg [63:0] modulo_result_rem_cmp_a;
  reg [63:0] modulo_result_rem_cmp_b;
  wire [63:0] modulo_result_rem_cmp_z;
  wire [63:0] operator_66_true_div_cmp_z_oreg;
  wire [9:0] fsm_output;
  wire or_tmp_1;
  wire nor_tmp_1;
  wire nor_tmp_2;
  wire or_tmp_11;
  wire or_tmp_19;
  wire or_tmp_29;
  wire and_dcpl;
  wire or_tmp_52;
  wire and_tmp_10;
  wire not_tmp_63;
  wire and_dcpl_20;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_25;
  wire and_dcpl_26;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_36;
  wire and_dcpl_37;
  wire and_dcpl_38;
  wire and_dcpl_41;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire and_dcpl_52;
  wire mux_tmp_106;
  wire and_dcpl_58;
  wire and_dcpl_61;
  wire and_dcpl_68;
  wire and_dcpl_73;
  wire and_dcpl_75;
  wire and_dcpl_79;
  wire not_tmp_94;
  wire and_dcpl_91;
  wire and_dcpl_93;
  wire mux_tmp_137;
  wire mux_tmp_138;
  wire or_tmp_154;
  wire and_dcpl_98;
  wire mux_tmp_146;
  wire and_tmp_11;
  wire not_tmp_111;
  wire and_dcpl_100;
  wire or_tmp_167;
  wire and_dcpl_106;
  wire nor_tmp_38;
  wire mux_tmp_157;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire or_tmp_189;
  wire mux_tmp_171;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_113;
  wire and_dcpl_119;
  wire not_tmp_141;
  wire and_dcpl_121;
  wire or_tmp_201;
  wire and_dcpl_127;
  wire or_tmp_204;
  wire and_dcpl_136;
  wire or_tmp_207;
  wire and_dcpl_137;
  wire and_dcpl_144;
  wire mux_tmp_185;
  wire mux_tmp_187;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_155;
  wire and_dcpl_157;
  wire or_tmp_263;
  wire and_dcpl_164;
  wire or_tmp_267;
  wire mux_tmp_236;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_171;
  wire and_tmp_17;
  wire or_tmp_271;
  wire or_tmp_273;
  wire or_tmp_279;
  wire and_dcpl_179;
  wire and_dcpl_181;
  wire or_tmp_283;
  wire mux_tmp_256;
  wire or_tmp_284;
  wire nor_tmp_56;
  wire nor_tmp_57;
  wire mux_tmp_263;
  wire nor_tmp_59;
  wire mux_tmp_269;
  wire mux_tmp_272;
  wire and_tmp_19;
  wire or_tmp_295;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_189;
  wire and_dcpl_190;
  wire mux_tmp_296;
  wire and_dcpl_193;
  wire and_dcpl_194;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire or_dcpl_39;
  wire or_dcpl_44;
  wire and_dcpl_202;
  wire or_tmp_335;
  wire mux_tmp_314;
  wire or_tmp_337;
  wire mux_tmp_320;
  wire or_tmp_341;
  wire mux_tmp_326;
  wire or_dcpl_58;
  wire and_dcpl_211;
  wire nor_tmp_77;
  wire nor_tmp_79;
  wire nor_tmp_81;
  wire and_dcpl_214;
  wire or_dcpl_62;
  wire or_dcpl_63;
  wire or_dcpl_68;
  wire or_dcpl_72;
  wire or_dcpl_82;
  wire or_dcpl_83;
  wire or_dcpl_84;
  wire or_dcpl_89;
  reg exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva;
  reg VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  reg [11:0] VEC_LOOP_j_1_12_0_sva_11_0;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg modExp_exp_1_0_1_sva;
  reg [11:0] COMP_LOOP_acc_10_cse_12_1_1_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_2_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_2_sva;
  reg [64:0] operator_64_false_acc_mut;
  reg [7:0] COMP_LOOP_k_9_1_1_sva_7_0;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_1_acc_8_itm;
  reg [11:0] reg_VEC_LOOP_1_acc_1_psp_ftd_1;
  wire and_171_m1c;
  wire and_178_m1c;
  reg reg_vec_rsc_triosy_0_1_obj_ld_cse;
  wire and_271_cse;
  wire or_492_cse;
  wire or_71_cse;
  wire and_282_cse;
  wire or_96_cse;
  wire or_100_cse;
  wire and_259_cse;
  wire or_89_cse;
  wire or_25_cse;
  wire and_334_cse;
  wire or_74_cse;
  wire nand_51_cse;
  wire or_52_cse;
  wire and_273_cse;
  wire or_210_cse;
  reg modExp_while_and_itm;
  reg modExp_while_and_1_itm;
  reg [9:0] reg_operator_66_true_div_cmp_b_reg;
  wire or_252_cse;
  reg [10:0] COMP_LOOP_acc_psp_1_sva;
  wire [63:0] COMP_LOOP_mux_1_itm_mx1;
  wire and_dcpl_232;
  wire [9:0] z_out;
  wire and_dcpl_234;
  wire and_dcpl_239;
  wire and_dcpl_241;
  wire and_dcpl_242;
  wire and_dcpl_244;
  wire and_dcpl_247;
  wire and_dcpl_249;
  wire and_dcpl_250;
  wire and_dcpl_253;
  wire and_dcpl_255;
  wire and_dcpl_256;
  wire and_dcpl_261;
  wire and_dcpl_262;
  wire and_dcpl_266;
  wire and_dcpl_267;
  wire and_dcpl_270;
  wire and_dcpl_272;
  wire and_dcpl_274;
  wire and_dcpl_276;
  wire and_dcpl_278;
  wire and_dcpl_281;
  wire and_dcpl_284;
  wire and_dcpl_287;
  wire [64:0] z_out_1;
  wire [10:0] z_out_2;
  wire [11:0] nl_z_out_2;
  wire [8:0] z_out_4;
  wire [9:0] nl_z_out_4;
  wire and_dcpl_343;
  reg [63:0] p_sva;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [63:0] modExp_result_sva;
  reg [63:0] tmp_2_lpi_4_dfm;
  reg modExp_exp_1_7_1_sva;
  reg modExp_exp_1_6_1_sva;
  reg modExp_exp_1_5_1_sva;
  reg modExp_exp_1_4_1_sva;
  reg modExp_exp_1_3_1_sva;
  reg modExp_exp_1_2_1_sva;
  reg modExp_exp_1_1_1_sva;
  reg modExp_exp_1_0_1_sva_1;
  reg [63:0] modExp_while_if_mul_mut;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_if_mul_mut;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_1_mul_mut;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_mul_mut;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_2_mul_mut;
  reg [63:0] VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_if_mul_mut;
  reg [63:0] VEC_LOOP_2_COMP_LOOP_1_mul_mut;
  reg [63:0] VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_mul_mut;
  reg [63:0] VEC_LOOP_2_COMP_LOOP_2_mul_mut;
  reg [63:0] modExp_while_mul_itm;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_mul_itm;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_if_mul_itm;
  reg [63:0] COMP_LOOP_mux_1_itm;
  reg [63:0] VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_mul_itm;
  reg [63:0] VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_if_mul_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [63:0] modulo_result_rem_cmp_a_mx0w0;
  wire [127:0] nl_modulo_result_rem_cmp_a_mx0w0;
  wire [63:0] VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w7;
  wire [64:0] nl_VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w7;
  wire [63:0] modExp_while_mul_itm_mx0w10;
  wire [127:0] nl_modExp_while_mul_itm_mx0w10;
  wire [63:0] VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
  wire signed [128:0] nl_VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire operator_64_false_acc_mut_mx0c0;
  wire VEC_LOOP_j_1_12_0_sva_11_0_mx0c1;
  wire modExp_result_sva_mx0c0;
  wire [62:0] operator_64_false_slc_modExp_exp_63_1_3;
  wire [63:0] modulo_qr_sva_1_mx0w8;
  wire [64:0] nl_modulo_qr_sva_1_mx0w8;
  wire VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c0;
  wire VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c1;
  wire tmp_2_lpi_4_dfm_mx0c1;
  wire modExp_1_while_and_11;
  wire modExp_result_and_rgt;
  wire modExp_result_and_1_rgt;
  wire COMP_LOOP_or_2_cse;
  wire COMP_LOOP_or_4_cse;
  wire mux_150_cse;
  wire nor_140_cse;
  wire mux_tmp;
  wire mux_195_itm;
  wire COMP_LOOP_nor_3_itm;
  wire COMP_LOOP_or_23_itm;
  wire COMP_LOOP_or_24_itm;
  wire z_out_5_8;
  wire mux_372_cse;
  wire and_468_cse;

  wire[0:0] and_105_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] nor_nl;
  wire[0:0] and_106_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] and_107_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] and_299_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] and_300_nl;
  wire[0:0] nor_152_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] and_301_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] nor_153_nl;
  wire[0:0] nor_154_nl;
  wire[0:0] nor_155_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] or_188_nl;
  wire[0:0] or_187_nl;
  wire[0:0] and_111_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] or_195_nl;
  wire[0:0] and_114_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] nor_151_nl;
  wire[0:0] nor_218_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] nand_80_nl;
  wire[0:0] or_512_nl;
  wire[0:0] mux_160_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] nor_144_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] nor_145_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] and_292_nl;
  wire[0:0] nor_146_nl;
  wire[0:0] nor_208_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] nand_64_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] nand_65_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] nor_209_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] or_500_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] nand_50_nl;
  wire[0:0] or_213_nl;
  wire[0:0] or_501_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] nand_52_nl;
  wire[0:0] nor_143_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] and_291_nl;
  wire[0:0] and_128_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] and_287_nl;
  wire[0:0] nor_138_nl;
  wire[0:0] and_130_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] nor_137_nl;
  wire[0:0] nor_214_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] or_509_nl;
  wire[0:0] nand_73_nl;
  wire[0:0] and_135_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] or_228_nl;
  wire[0:0] and_138_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] or_493_nl;
  wire[0:0] nor_135_nl;
  wire[0:0] and_141_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] and_285_nl;
  wire[0:0] nor_134_nl;
  wire[0:0] and_145_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] and_284_nl;
  wire[0:0] nor_133_nl;
  wire[0:0] and_147_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] and_148_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] nor_132_nl;
  wire[0:0] nand_85_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] nor_128_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] nor_129_nl;
  wire[0:0] nor_130_nl;
  wire[0:0] nor_131_nl;
  wire[0:0] and_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] nor_248_nl;
  wire[0:0] nor_249_nl;
  wire[0:0] nor_250_nl;
  wire[0:0] nor_251_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] nor_124_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] or_296_nl;
  wire[0:0] or_294_nl;
  wire[0:0] and_176_nl;
  wire[0:0] r_or_nl;
  wire[0:0] r_or_1_nl;
  wire[0:0] and_189_nl;
  wire[0:0] and_193_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] or_533_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] or_314_nl;
  wire[0:0] or_312_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] and_195_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] nor_122_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] or_534_nl;
  wire[0:0] COMP_LOOP_and_nl;
  wire[0:0] COMP_LOOP_and_1_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] or_329_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] nor_120_nl;
  wire[0:0] and_276_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] or_325_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] or_324_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] or_323_nl;
  wire[0:0] or_322_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] or_319_nl;
  wire[0:0] COMP_LOOP_mux1h_13_nl;
  wire[0:0] COMP_LOOP_and_5_nl;
  wire[0:0] and_212_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] nor_113_nl;
  wire[0:0] nor_114_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] nor_115_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] nand_48_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] and_270_nl;
  wire[0:0] or_344_nl;
  wire[0:0] nor_116_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] or_341_nl;
  wire[0:0] or_339_nl;
  wire[0:0] mux_303_nl;
  wire[9:0] VEC_LOOP_1_COMP_LOOP_1_acc_11_nl;
  wire[10:0] nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl;
  wire[11:0] COMP_LOOP_mux_21_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] mux_317_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] nor_70_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] or_396_nl;
  wire[0:0] or_394_nl;
  wire[0:0] and_230_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] and_339_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] and_341_nl;
  wire[0:0] nor_102_nl;
  wire[0:0] nor_103_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] nor_104_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] and_268_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] nor_107_nl;
  wire[0:0] nor_108_nl;
  wire[0:0] COMP_LOOP_mux1h_23_nl;
  wire[0:0] nor_213_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] nand_42_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] and_257_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] and_258_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] and_260_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] COMP_LOOP_mux1h_40_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] or_438_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] and_247_nl;
  wire[0:0] nand_37_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] or_466_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] and_246_nl;
  wire[0:0] nand_36_nl;
  wire[0:0] or_496_nl;
  wire[0:0] nor_190_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] or_105_nl;
  wire[0:0] or_123_nl;
  wire[0:0] nor_148_nl;
  wire[0:0] nor_149_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] or_511_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] or_201_nl;
  wire[0:0] nand_78_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] or_238_nl;
  wire[0:0] or_246_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] or_267_nl;
  wire[0:0] or_36_nl;
  wire[0:0] nand_28_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] or_42_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] or_303_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] or_318_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] nor_118_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] or_336_nl;
  wire[0:0] nor_119_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] or_354_nl;
  wire[0:0] and_272_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] or_347_nl;
  wire[0:0] or_346_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] nor_99_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] nand_43_nl;
  wire[0:0] nor_100_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] nand_70_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] and_249_nl;
  wire[0:0] and_250_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] and_335_nl;
  wire[0:0] and_336_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] nand_71_nl;
  wire[0:0] nand_72_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] and_337_nl;
  wire[0:0] and_338_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] or_47_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] or_257_nl;
  wire[0:0] nand_74_nl;
  wire[0:0] nor_125_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] or_400_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] or_302_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] or_298_nl;
  wire[0:0] nor_220_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] nand_83_nl;
  wire[0:0] or_513_nl;
  wire[0:0] and_65_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] nor_185_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] and_314_nl;
  wire[0:0] nor_186_nl;
  wire[0:0] nor_187_nl;
  wire[0:0] and_67_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] nor_183_nl;
  wire[0:0] and_313_nl;
  wire[0:0] nor_184_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] nand_69_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] nor_177_nl;
  wire[0:0] nor_178_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] or_140_nl;
  wire[0:0] or_139_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] or_505_nl;
  wire[0:0] or_506_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] or_507_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] or_133_nl;
  wire[0:0] or_131_nl;
  wire[0:0] or_508_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] and_310_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] and_311_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] nor_170_nl;
  wire[0:0] nor_171_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] nor_172_nl;
  wire[0:0] nor_173_nl;
  wire[0:0] nor_174_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] nor_175_nl;
  wire[0:0] nor_176_nl;
  wire[0:0] or_147_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] nand_63_nl;
  wire[0:0] or_144_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] nand_67_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] and_340_nl;
  wire[0:0] and_308_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] nor_163_nl;
  wire[0:0] nor_164_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] or_502_nl;
  wire[0:0] or_503_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] nand_68_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] nor_167_nl;
  wire[0:0] nor_168_nl;
  wire[0:0] or_504_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] and_304_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] and_305_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] and_306_nl;
  wire[0:0] nor_156_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] nor_157_nl;
  wire[0:0] nor_158_nl;
  wire[0:0] nor_159_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] nand_12_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] nor_160_nl;
  wire[0:0] nor_161_nl;
  wire[0:0] or_173_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] or_172_nl;
  wire[0:0] or_170_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] nor_233_nl;
  wire[0:0] nor_234_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] or_nl;
  wire[0:0] or_532_nl;
  wire[0:0] nand_86_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] nor_232_nl;
  wire[0:0] and_466_nl;
  wire[0:0] nor_224_nl;
  wire[0:0] nor_225_nl;
  wire[0:0] or_537_nl;
  wire[0:0] or_536_nl;
  wire[10:0] acc_nl;
  wire[11:0] nl_acc_nl;
  wire[9:0] COMP_LOOP_mux_18_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nand_1_nl;
  wire[65:0] acc_1_nl;
  wire[66:0] nl_acc_1_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_53_nl;
  wire[0:0] COMP_LOOP_mux_19_nl;
  wire[50:0] COMP_LOOP_or_31_nl;
  wire[50:0] COMP_LOOP_and_65_nl;
  wire[50:0] COMP_LOOP_mux1h_70_nl;
  wire[1:0] COMP_LOOP_or_32_nl;
  wire[1:0] COMP_LOOP_and_66_nl;
  wire[1:0] COMP_LOOP_mux1h_71_nl;
  wire[0:0] COMP_LOOP_nor_60_nl;
  wire[9:0] COMP_LOOP_mux1h_72_nl;
  wire[8:0] COMP_LOOP_acc_18_nl;
  wire[9:0] nl_COMP_LOOP_acc_18_nl;
  wire[0:0] COMP_LOOP_or_33_nl;
  wire[0:0] COMP_LOOP_or_34_nl;
  wire[0:0] COMP_LOOP_or_35_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_54_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_55_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_56_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_57_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_58_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_59_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_60_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_61_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_62_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_63_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_64_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_65_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_66_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_67_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_68_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_69_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_70_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_71_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_72_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_73_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_74_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_75_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_76_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_77_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_78_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_79_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_80_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_81_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_82_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_83_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_84_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_85_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_86_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_87_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_88_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_89_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_90_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_91_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_92_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_93_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_94_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_95_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_96_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_97_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_98_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_99_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_100_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_101_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_102_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_103_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_104_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_105_nl;
  wire[1:0] COMP_LOOP_or_36_nl;
  wire[1:0] COMP_LOOP_and_67_nl;
  wire[1:0] COMP_LOOP_mux1h_73_nl;
  wire[0:0] COMP_LOOP_nor_62_nl;
  wire[9:0] COMP_LOOP_or_37_nl;
  wire[9:0] COMP_LOOP_mux1h_74_nl;
  wire[0:0] COMP_LOOP_or_38_nl;
  wire[0:0] COMP_LOOP_or_39_nl;
  wire[10:0] COMP_LOOP_mux_20_nl;
  wire[7:0] STAGE_LOOP_mux_2_nl;
  wire[8:0] operator_64_false_1_acc_nl;
  wire[9:0] nl_operator_64_false_1_acc_nl;
  wire[0:0] operator_64_false_1_mux_10_nl;
  wire[0:0] operator_64_false_1_mux_11_nl;
  wire[0:0] operator_64_false_1_mux_12_nl;
  wire[0:0] operator_64_false_1_mux_13_nl;
  wire[0:0] operator_64_false_1_mux_14_nl;
  wire[0:0] operator_64_false_1_mux_15_nl;
  wire[0:0] operator_64_false_1_mux_16_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[64:0] operator_64_false_acc_1_nl;
  wire[65:0] nl_operator_64_false_acc_1_nl;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_10_tr0;
  assign nl_operator_64_false_acc_1_nl = ({1'b1 , (~ operator_66_true_div_cmp_z_oreg)})
      + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_acc_1_nl = nl_operator_64_false_acc_1_nl[64:0];
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_10_tr0 = ~ (readslicef_65_1_64(operator_64_false_acc_1_nl));
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0 = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_76_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_76_tr0 = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_1[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0 = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_76_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_76_tr0 = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0 = z_out_1[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_11_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_11_tr0 = ~ (z_out_1[2]);
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_1_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_1_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_1_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_1_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd1)) modulo_result_rem_cmp (
      .a(modulo_result_rem_cmp_a),
      .b(modulo_result_rem_cmp_b),
      .z(modulo_result_rem_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_wait_dp inPlaceNTT_DIT_core_wait_dp_inst (
      .clk(clk),
      .operator_66_true_div_cmp_z(operator_66_true_div_cmp_z),
      .operator_66_true_div_cmp_z_oreg(operator_66_true_div_cmp_z_oreg)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_10_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_10_tr0[0:0]),
      .modExp_while_C_47_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_1_COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_47_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_1_COMP_LOOP_C_76_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_76_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_47_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_C_152_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_47_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_2_COMP_LOOP_C_76_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_76_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_47_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_C_152_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0[0:0]),
      .STAGE_LOOP_C_11_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_11_tr0[0:0])
    );
  assign nand_51_cse = ~((fsm_output[2:1]==2'b11));
  assign or_210_cse = (fsm_output[1]) | (fsm_output[7]);
  assign nor_140_cse = ~((fsm_output[1:0]!=2'b00));
  assign operator_66_true_div_cmp_b = {1'b0, reg_operator_66_true_div_cmp_b_reg};
  assign or_96_cse = (fsm_output[3:2]!=2'b00);
  assign and_282_cse = (fsm_output[1:0]==2'b11);
  assign and_171_m1c = and_dcpl_75 & and_dcpl_36;
  assign modExp_result_and_rgt = (~ modExp_while_and_1_itm) & and_171_m1c;
  assign modExp_result_and_1_rgt = modExp_while_and_1_itm & and_171_m1c;
  assign or_89_cse = (fsm_output[3:1]!=3'b100);
  assign and_271_cse = (fsm_output[2:1]==2'b11);
  assign or_492_cse = (fsm_output[2:1]!=2'b00);
  assign COMP_LOOP_or_2_cse = (and_dcpl_38 & and_dcpl_33 & and_dcpl_36) | ((fsm_output[3:1]==3'b011)
      & and_dcpl_33 & and_dcpl_61 & (~ (fsm_output[6])) & and_dcpl_20);
  assign or_71_cse = (fsm_output[1:0]!=2'b00);
  assign or_74_cse = (fsm_output[8:7]!=2'b00);
  assign and_259_cse = (fsm_output[5:4]==2'b11);
  assign COMP_LOOP_or_4_cse = (and_dcpl_44 & and_dcpl_24 & and_dcpl_41 & and_dcpl_20)
      | (and_dcpl_58 & and_dcpl_24 & and_dcpl_41 & and_dcpl) | (and_dcpl_37 & (~
      (fsm_output[2])) & and_dcpl_24 & and_dcpl_68 & and_dcpl_20) | (and_dcpl_75
      & and_dcpl_73);
  assign nl_modulo_result_rem_cmp_a_mx0w0 = modExp_result_sva * COMP_LOOP_mux_1_itm;
  assign modulo_result_rem_cmp_a_mx0w0 = nl_modulo_result_rem_cmp_a_mx0w0[63:0];
  assign or_52_cse = (fsm_output[3:1]!=3'b011);
  assign nl_VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w7 = tmp_2_lpi_4_dfm + COMP_LOOP_mux_1_itm_mx1;
  assign VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w7 = nl_VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w7[63:0];
  assign nl_modExp_while_mul_itm_mx0w10 = COMP_LOOP_mux_1_itm * COMP_LOOP_mux_1_itm;
  assign modExp_while_mul_itm_mx0w10 = nl_modExp_while_mul_itm_mx0w10[63:0];
  assign nl_VEC_LOOP_1_COMP_LOOP_1_mul_mut_1 = $signed(VEC_LOOP_1_COMP_LOOP_1_acc_8_itm)
      * $signed(conv_u2s_64_65(COMP_LOOP_mux_1_itm));
  assign VEC_LOOP_1_COMP_LOOP_1_mul_mut_1 = nl_VEC_LOOP_1_COMP_LOOP_1_mul_mut_1[63:0];
  assign and_334_cse = (fsm_output[3:0]==4'b1111);
  assign operator_64_false_slc_modExp_exp_63_1_3 = MUX_v_63_2_2((operator_66_true_div_cmp_z_oreg[63:1]),
      (VEC_LOOP_1_COMP_LOOP_1_acc_8_itm[63:1]), and_dcpl_157);
  assign nl_modulo_qr_sva_1_mx0w8 = (operator_64_false_acc_mut[63:0]) + p_sva;
  assign modulo_qr_sva_1_mx0w8 = nl_modulo_qr_sva_1_mx0w8[63:0];
  assign COMP_LOOP_mux_1_itm_mx1 = MUX_v_64_2_2((operator_64_false_acc_mut[63:0]),
      modulo_qr_sva_1_mx0w8, operator_64_false_acc_mut[63]);
  assign modExp_1_while_and_11 = (operator_64_false_acc_mut[63]) & modExp_exp_1_0_1_sva;
  assign or_tmp_1 = (fsm_output[8:6]!=3'b000);
  assign nor_tmp_1 = or_492_cse & (fsm_output[3]);
  assign nor_tmp_2 = (fsm_output[3:2]==2'b11);
  assign or_tmp_11 = (fsm_output[3:1]!=3'b010);
  assign or_25_cse = (fsm_output[3:1]!=3'b000);
  assign or_tmp_19 = and_271_cse | (fsm_output[3]);
  assign or_tmp_29 = (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[2]);
  assign and_dcpl = (fsm_output[7]) & (~ (fsm_output[9]));
  assign or_tmp_52 = (~ (fsm_output[7])) | (fsm_output[9]);
  assign or_100_cse = (fsm_output[3:0]!=4'b0000);
  assign and_tmp_10 = (fsm_output[4]) & or_100_cse;
  assign or_496_nl = (fsm_output[8:0]!=9'b000000000);
  assign or_105_nl = (fsm_output[8]) | and_tmp_10;
  assign mux_99_nl = MUX_s_1_2_2((fsm_output[8]), or_105_nl, fsm_output[5]);
  assign nor_190_nl = ~((fsm_output[7:6]!=2'b00) | mux_99_nl);
  assign not_tmp_63 = MUX_s_1_2_2(or_496_nl, nor_190_nl, fsm_output[9]);
  assign and_dcpl_20 = ~((fsm_output[7]) | (fsm_output[9]));
  assign and_dcpl_23 = ~((fsm_output[8]) | (fsm_output[5]) | (fsm_output[6]) | (~
      and_dcpl_20));
  assign and_dcpl_24 = ~((fsm_output[0]) | (fsm_output[4]));
  assign and_dcpl_25 = ~((fsm_output[3]) | (fsm_output[1]));
  assign and_dcpl_26 = and_dcpl_25 & (~ (fsm_output[2]));
  assign and_dcpl_30 = (~ (fsm_output[8])) & (fsm_output[5]);
  assign and_dcpl_31 = and_dcpl_30 & (~ (fsm_output[6]));
  assign and_dcpl_32 = and_dcpl_31 & (~ (fsm_output[7])) & (fsm_output[9]);
  assign and_dcpl_33 = (~ (fsm_output[0])) & (fsm_output[4]);
  assign and_dcpl_36 = and_dcpl_31 & and_dcpl_20;
  assign and_dcpl_37 = (fsm_output[3]) & (~ (fsm_output[1]));
  assign and_dcpl_38 = and_dcpl_37 & (fsm_output[2]);
  assign and_dcpl_41 = and_dcpl_30 & (fsm_output[6]);
  assign and_dcpl_43 = (fsm_output[3]) & (fsm_output[1]);
  assign and_dcpl_44 = and_dcpl_43 & (fsm_output[2]);
  assign and_dcpl_52 = (fsm_output[0]) & (fsm_output[5]);
  assign or_123_nl = (fsm_output[3:1]!=3'b001);
  assign mux_tmp_106 = MUX_s_1_2_2(or_89_cse, or_123_nl, fsm_output[8]);
  assign and_dcpl_58 = and_dcpl_43 & (~ (fsm_output[2]));
  assign and_dcpl_61 = (fsm_output[8]) & (fsm_output[5]);
  assign and_dcpl_68 = and_dcpl_61 & (fsm_output[6]);
  assign and_dcpl_73 = and_dcpl_68 & and_dcpl;
  assign and_dcpl_75 = and_dcpl_25 & (fsm_output[2]) & and_dcpl_24;
  assign and_dcpl_79 = (~ (fsm_output[0])) & (fsm_output[5]) & (~ (fsm_output[9]));
  assign not_tmp_94 = ~((COMP_LOOP_acc_1_cse_2_sva[0]) & (fsm_output[7]));
  assign and_dcpl_91 = and_dcpl_38 & and_dcpl_24 & and_dcpl_23;
  assign and_dcpl_93 = (~ (fsm_output[8])) & (~ (fsm_output[6])) & and_dcpl_20;
  assign mux_tmp_137 = MUX_s_1_2_2(or_96_cse, or_25_cse, fsm_output[0]);
  assign mux_tmp_138 = MUX_s_1_2_2(and_dcpl_44, nor_tmp_2, fsm_output[0]);
  assign or_tmp_154 = (fsm_output[4]) | mux_tmp_138;
  assign and_dcpl_98 = ~((fsm_output[9:7]!=3'b000));
  assign mux_tmp_146 = MUX_s_1_2_2(or_tmp_19, or_96_cse, fsm_output[0]);
  assign and_tmp_11 = (fsm_output[4]) & mux_tmp_146;
  assign not_tmp_111 = ~((fsm_output[5:0]==6'b111111));
  assign and_dcpl_100 = (~ (fsm_output[8])) & (fsm_output[6]);
  assign or_tmp_167 = ((fsm_output[2:0]==3'b111)) | (fsm_output[3]);
  assign nor_148_nl = ~((fsm_output[8]) | (~ (fsm_output[3])));
  assign nor_149_nl = ~((~ (fsm_output[8])) | (fsm_output[3]));
  assign mux_150_cse = MUX_s_1_2_2(nor_148_nl, nor_149_nl, fsm_output[1]);
  assign nand_17_nl = ~((fsm_output[7]) & mux_150_cse);
  assign or_201_nl = (fsm_output[7]) | (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[3]);
  assign mux_151_nl = MUX_s_1_2_2(nand_17_nl, or_201_nl, fsm_output[2]);
  assign or_511_nl = (fsm_output[6:5]!=2'b00) | mux_151_nl;
  assign nand_78_nl = ~((fsm_output[5]) & (fsm_output[6]) & (fsm_output[2]) & (fsm_output[7])
      & (fsm_output[1]) & (fsm_output[8]) & (fsm_output[3]));
  assign mux_152_nl = MUX_s_1_2_2(or_511_nl, nand_78_nl, fsm_output[4]);
  assign and_dcpl_106 = ~(mux_152_nl | (fsm_output[0]) | (fsm_output[9]));
  assign nor_tmp_38 = ((fsm_output[2:0]!=3'b000)) & (fsm_output[3]);
  assign mux_tmp_157 = MUX_s_1_2_2(nor_tmp_2, nor_tmp_1, fsm_output[0]);
  assign and_dcpl_108 = and_259_cse & (~ (fsm_output[6]));
  assign and_dcpl_109 = and_dcpl_108 & and_dcpl;
  assign or_tmp_189 = (fsm_output[2]) | (~ and_dcpl_43);
  assign mux_tmp_171 = MUX_s_1_2_2(or_tmp_189, or_tmp_11, fsm_output[8]);
  assign and_dcpl_110 = ~(mux_tmp_171 | (fsm_output[0]));
  assign and_dcpl_111 = and_dcpl_110 & and_dcpl_109;
  assign and_dcpl_113 = (fsm_output[9:7]==3'b001);
  assign and_dcpl_119 = (fsm_output[9:7]==3'b010);
  assign not_tmp_141 = ~((fsm_output[5:4]==2'b11) & nor_tmp_38);
  assign and_dcpl_121 = (fsm_output[8]) & (fsm_output[6]);
  assign or_tmp_201 = (fsm_output[4]) | mux_tmp_157;
  assign and_dcpl_127 = (fsm_output[9:7]==3'b011);
  assign or_tmp_204 = (fsm_output[4:1]!=4'b0000);
  assign and_dcpl_136 = ~((~(or_492_cse ^ (fsm_output[3]))) | (fsm_output[4]) | (fsm_output[8])
      | (fsm_output[5]) | (fsm_output[6]) | (~ and_dcpl_20));
  assign or_238_nl = (fsm_output[8]) | (fsm_output[4]);
  assign mux_181_nl = MUX_s_1_2_2((fsm_output[8]), or_238_nl, fsm_output[5]);
  assign or_tmp_207 = (fsm_output[7:6]!=2'b00) | mux_181_nl;
  assign and_dcpl_137 = (fsm_output[0]) & (~ (fsm_output[4]));
  assign and_dcpl_144 = and_dcpl_58 & (~((fsm_output[4]) ^ (fsm_output[5]))) & (fsm_output[0])
      & (~ (fsm_output[8])) & (~ (fsm_output[6])) & and_dcpl_20;
  assign or_246_nl = (~ (fsm_output[8])) | (~ (fsm_output[7])) | (fsm_output[2])
      | (fsm_output[9]) | (fsm_output[6]);
  assign or_267_nl = (~ (fsm_output[7])) | (~ (fsm_output[2])) | (fsm_output[9])
      | (fsm_output[6]);
  assign or_36_nl = (fsm_output[7]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[2]);
  assign mux_184_nl = MUX_s_1_2_2(or_267_nl, or_36_nl, fsm_output[8]);
  assign mux_tmp_185 = MUX_s_1_2_2(or_246_nl, mux_184_nl, fsm_output[1]);
  assign or_42_nl = (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[2]));
  assign mux_32_nl = MUX_s_1_2_2(or_42_nl, or_tmp_29, fsm_output[7]);
  assign nand_28_nl = ~((fsm_output[8]) & (fsm_output[1]) & (~ mux_32_nl));
  assign mux_tmp_187 = MUX_s_1_2_2(nand_28_nl, mux_tmp_185, fsm_output[4]);
  assign mux_188_nl = MUX_s_1_2_2((fsm_output[6]), (~ (fsm_output[6])), fsm_output[9]);
  assign nand_23_nl = ~((fsm_output[2]) & mux_188_nl);
  assign mux_189_nl = MUX_s_1_2_2(nand_23_nl, or_tmp_29, fsm_output[7]);
  assign or_252_cse = (fsm_output[1]) | (fsm_output[8]) | mux_189_nl;
  assign and_dcpl_151 = (fsm_output[6:4]==3'b110);
  assign and_dcpl_152 = and_dcpl_151 & and_dcpl;
  assign and_dcpl_153 = and_dcpl_110 & and_dcpl_152;
  assign and_dcpl_155 = (fsm_output[0]) & (fsm_output[4]);
  assign and_dcpl_157 = and_dcpl_58 & and_dcpl_155 & and_dcpl_36;
  assign or_tmp_263 = (fsm_output[4:1]!=4'b0110);
  assign and_dcpl_164 = and_dcpl_155 & (fsm_output[5]) & (~ (fsm_output[6])) & (~
      (fsm_output[9]));
  assign or_tmp_267 = (fsm_output[1]) | (~ (fsm_output[3]));
  assign or_303_nl = (~ (fsm_output[1])) | (fsm_output[3]);
  assign mux_tmp_236 = MUX_s_1_2_2(or_tmp_267, or_303_nl, fsm_output[8]);
  assign and_dcpl_165 = ~(mux_tmp_236 | (~((fsm_output[2]) ^ (fsm_output[7]))));
  assign and_dcpl_166 = and_dcpl_165 & and_dcpl_164;
  assign and_dcpl_167 = (fsm_output[6]) & (~ (fsm_output[9]));
  assign mux_237_nl = MUX_s_1_2_2((~ and_dcpl_44), or_89_cse, fsm_output[8]);
  assign mux_238_nl = MUX_s_1_2_2(mux_237_nl, mux_tmp_171, fsm_output[7]);
  assign and_dcpl_171 = (~ mux_238_nl) & (fsm_output[0]);
  assign and_tmp_17 = (fsm_output[4]) & or_96_cse;
  assign or_tmp_271 = (fsm_output[4:0]!=5'b10100);
  assign or_tmp_273 = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[2]) | (~
      and_dcpl_43);
  assign or_tmp_279 = (fsm_output[4:0]!=5'b01100);
  assign and_dcpl_179 = (fsm_output[7:5]==3'b110);
  assign or_318_nl = (fsm_output[4:1]!=4'b1001);
  assign mux_255_nl = MUX_s_1_2_2(or_318_nl, or_tmp_263, fsm_output[8]);
  assign and_dcpl_181 = ~(mux_255_nl | (fsm_output[0]));
  assign or_tmp_283 = (fsm_output[6]) | (fsm_output[4]);
  assign mux_tmp_256 = MUX_s_1_2_2((fsm_output[6]), or_tmp_283, fsm_output[5]);
  assign or_tmp_284 = (fsm_output[7]) | mux_tmp_256;
  assign nor_tmp_56 = (fsm_output[6:5]==2'b11);
  assign nor_tmp_57 = (fsm_output[6:4]==3'b111);
  assign mux_tmp_263 = MUX_s_1_2_2((~ or_tmp_283), (fsm_output[4]), fsm_output[5]);
  assign nor_tmp_59 = (fsm_output[6]) & (fsm_output[4]);
  assign mux_tmp_269 = MUX_s_1_2_2((~ or_tmp_283), nor_tmp_59, fsm_output[5]);
  assign mux_271_nl = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[6]);
  assign mux_tmp_272 = MUX_s_1_2_2(mux_271_nl, nor_tmp_59, fsm_output[5]);
  assign and_tmp_19 = (fsm_output[5]) & or_tmp_283;
  assign or_tmp_295 = (~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[3]);
  assign or_336_nl = (fsm_output[8]) | (~ (fsm_output[2])) | (fsm_output[3]);
  assign mux_291_nl = MUX_s_1_2_2(or_tmp_295, or_336_nl, fsm_output[1]);
  assign nor_118_nl = ~((~ (fsm_output[4])) | (fsm_output[5]) | (fsm_output[7]) |
      mux_291_nl);
  assign or_354_nl = (fsm_output[8]) | (fsm_output[2]) | (~ (fsm_output[3]));
  assign mux_290_nl = MUX_s_1_2_2(or_354_nl, or_tmp_295, fsm_output[1]);
  assign nor_119_nl = ~((fsm_output[4]) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | mux_290_nl);
  assign mux_292_nl = MUX_s_1_2_2(nor_118_nl, nor_119_nl, fsm_output[0]);
  assign and_dcpl_186 = mux_292_nl & and_dcpl_167;
  assign and_dcpl_187 = and_dcpl_108 & and_dcpl_20;
  assign and_dcpl_189 = (~ mux_tmp_236) & (fsm_output[2]) & (fsm_output[0]);
  assign and_dcpl_190 = and_dcpl_189 & and_dcpl_187;
  assign and_273_cse = (fsm_output[2]) & (fsm_output[7]);
  assign and_272_nl = (fsm_output[2]) & (fsm_output[7]) & (fsm_output[8]);
  assign or_347_nl = and_273_cse | (fsm_output[8]);
  assign or_346_nl = (fsm_output[2]) | (fsm_output[7]) | (fsm_output[8]);
  assign mux_295_nl = MUX_s_1_2_2(or_347_nl, or_346_nl, fsm_output[1]);
  assign mux_tmp_296 = MUX_s_1_2_2(and_272_nl, mux_295_nl, fsm_output[3]);
  assign and_dcpl_193 = (~ mux_tmp_236) & (~ (fsm_output[2])) & (fsm_output[0]);
  assign and_dcpl_194 = and_dcpl_193 & and_dcpl_109;
  assign mux_304_nl = MUX_s_1_2_2(nand_51_cse, or_492_cse, fsm_output[8]);
  assign and_dcpl_197 = (~ mux_304_nl) & (fsm_output[3]) & (~ (fsm_output[0]));
  assign and_dcpl_198 = and_dcpl_197 & and_dcpl_187;
  assign or_dcpl_39 = (fsm_output[7]) | (fsm_output[9]);
  assign or_dcpl_44 = or_tmp_267 | (~ (fsm_output[2]));
  assign and_dcpl_202 = and_dcpl_151 & and_dcpl_20;
  assign or_tmp_335 = (fsm_output[9]) | (~((fsm_output[7:6]!=2'b00)));
  assign mux_tmp_314 = MUX_s_1_2_2(or_tmp_335, (fsm_output[9]), fsm_output[5]);
  assign or_tmp_337 = (fsm_output[9]) | (~ or_tmp_1);
  assign mux_319_nl = MUX_s_1_2_2((~ or_tmp_1), or_tmp_1, fsm_output[9]);
  assign mux_tmp_320 = MUX_s_1_2_2(mux_319_nl, or_tmp_335, fsm_output[5]);
  assign or_tmp_341 = ~((fsm_output[8]) & (fsm_output[2]) & (fsm_output[1]) & (~
      (fsm_output[3])));
  assign mux_tmp_326 = MUX_s_1_2_2(or_dcpl_44, or_52_cse, fsm_output[8]);
  assign or_dcpl_58 = ~((fsm_output[0]) & (fsm_output[4]));
  assign nand_43_nl = ~((fsm_output[3:1]==3'b111));
  assign mux_342_nl = MUX_s_1_2_2(nand_43_nl, or_89_cse, fsm_output[8]);
  assign nor_99_nl = ~((~ (fsm_output[4])) | (fsm_output[6]) | (fsm_output[7]) |
      mux_342_nl);
  assign nor_100_nl = ~((fsm_output[4]) | (~ (fsm_output[6])) | (~ (fsm_output[7]))
      | mux_tmp_106);
  assign mux_343_nl = MUX_s_1_2_2(nor_99_nl, nor_100_nl, fsm_output[0]);
  assign and_dcpl_211 = mux_343_nl & (fsm_output[5]) & (~ (fsm_output[9]));
  assign nor_tmp_77 = ((fsm_output[2]) | (fsm_output[7]) | (fsm_output[4])) & (fsm_output[5]);
  assign nor_tmp_79 = (and_273_cse | (fsm_output[4])) & (fsm_output[5]);
  assign nor_tmp_81 = (fsm_output[2]) & (fsm_output[7]) & (fsm_output[4]) & (fsm_output[5]);
  assign and_249_nl = ((fsm_output[0]) | (fsm_output[7])) & (fsm_output[8]) & (fsm_output[4])
      & (fsm_output[5]);
  assign and_250_nl = or_74_cse & (fsm_output[5:4]==2'b11);
  assign mux_358_nl = MUX_s_1_2_2(and_249_nl, and_250_nl, fsm_output[1]);
  assign nand_70_nl = ~((fsm_output[3]) & mux_358_nl);
  assign and_335_nl = (((fsm_output[1]) & (fsm_output[0]) & (fsm_output[7]) & (fsm_output[8]))
      | (fsm_output[4])) & (fsm_output[5]);
  assign and_336_nl = ((or_71_cse & (fsm_output[7])) | (fsm_output[8]) | (fsm_output[4]))
      & (fsm_output[5]);
  assign mux_357_nl = MUX_s_1_2_2(and_335_nl, and_336_nl, fsm_output[3]);
  assign mux_359_nl = MUX_s_1_2_2(nand_70_nl, mux_357_nl, fsm_output[6]);
  assign nand_71_nl = ~((fsm_output[7]) & (fsm_output[8]) & (fsm_output[4]) & (fsm_output[5]));
  assign nand_72_nl = ~((and_282_cse | (fsm_output[8:7]!=2'b00)) & (fsm_output[5:4]==2'b11));
  assign mux_355_nl = MUX_s_1_2_2(nand_71_nl, nand_72_nl, fsm_output[3]);
  assign and_337_nl = (((fsm_output[8:7]==2'b11)) | (fsm_output[4])) & (fsm_output[5]);
  assign and_338_nl = ((fsm_output[1]) | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[4]))
      & (fsm_output[5]);
  assign mux_354_nl = MUX_s_1_2_2(and_337_nl, and_338_nl, fsm_output[3]);
  assign mux_356_nl = MUX_s_1_2_2(mux_355_nl, mux_354_nl, fsm_output[6]);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, mux_356_nl, fsm_output[2]);
  assign and_dcpl_214 = ~(mux_360_nl | (fsm_output[9]));
  assign or_dcpl_62 = (fsm_output[8]) | (~ (fsm_output[5]));
  assign or_dcpl_63 = or_dcpl_62 | (fsm_output[6]);
  assign or_dcpl_68 = (fsm_output[0]) | (fsm_output[4]);
  assign or_dcpl_72 = or_dcpl_62 | (~ (fsm_output[6]));
  assign or_dcpl_82 = ~((fsm_output[8]) & (fsm_output[5]));
  assign or_dcpl_83 = or_dcpl_82 | (fsm_output[6]);
  assign or_dcpl_84 = or_dcpl_83 | or_dcpl_39;
  assign or_dcpl_89 = or_dcpl_82 | (~ (fsm_output[6]));
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_26 & and_dcpl_33 & and_dcpl_32;
  assign operator_64_false_acc_mut_mx0c0 = and_dcpl_26 & and_dcpl_137 & and_dcpl_23;
  assign or_47_nl = (fsm_output[8]) | (~ (fsm_output[1])) | (fsm_output[7]) | (fsm_output[6])
      | (fsm_output[9]) | (fsm_output[2]);
  assign mux_210_nl = MUX_s_1_2_2(or_252_cse, or_47_nl, fsm_output[4]);
  assign mux_194_nl = MUX_s_1_2_2(mux_tmp_187, mux_210_nl, fsm_output[3]);
  assign nand_24_nl = ~((fsm_output[5]) & (~ mux_194_nl));
  assign mux_190_nl = MUX_s_1_2_2(mux_tmp_185, or_252_cse, fsm_output[4]);
  assign mux_191_nl = MUX_s_1_2_2(mux_190_nl, mux_tmp_187, fsm_output[3]);
  assign or_257_nl = (fsm_output[4]) | (fsm_output[8]) | (~ (fsm_output[1])) | (fsm_output[7])
      | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[6]);
  assign nand_74_nl = ~((fsm_output[4]) & (fsm_output[8]) & (~ (fsm_output[1])) &
      (fsm_output[7]) & (fsm_output[6]) & (~ (fsm_output[9])) & (fsm_output[2]));
  assign mux_183_nl = MUX_s_1_2_2(or_257_nl, nand_74_nl, fsm_output[3]);
  assign mux_192_nl = MUX_s_1_2_2(mux_191_nl, mux_183_nl, fsm_output[5]);
  assign mux_195_itm = MUX_s_1_2_2(nand_24_nl, mux_192_nl, fsm_output[0]);
  assign VEC_LOOP_j_1_12_0_sva_11_0_mx0c1 = and_dcpl_44 & and_dcpl_137 & and_dcpl_32;
  assign nor_125_nl = ~((fsm_output[8:4]!=5'b00000) | nor_tmp_2);
  assign modExp_result_sva_mx0c0 = MUX_s_1_2_2(nor_125_nl, or_tmp_207, fsm_output[9]);
  assign VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c0
      = (~ mux_tmp_236) & (fsm_output[2]) & (~ (fsm_output[0])) & and_dcpl_187;
  assign VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c1
      = and_dcpl_197 & and_dcpl_202;
  assign or_400_nl = (~ (VEC_LOOP_j_1_12_0_sva_11_0[0])) | (fsm_output[8]) | (~ (fsm_output[2]))
      | (fsm_output[1]) | (~ (fsm_output[3]));
  assign mux_330_nl = MUX_s_1_2_2(or_tmp_341, mux_tmp_326, VEC_LOOP_j_1_12_0_sva_11_0[0]);
  assign mux_331_nl = MUX_s_1_2_2(or_400_nl, mux_330_nl, reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]);
  assign nand_32_nl = ~((COMP_LOOP_acc_1_cse_2_sva[0]) & (~ mux_tmp_106));
  assign mux_332_nl = MUX_s_1_2_2(mux_331_nl, nand_32_nl, fsm_output[7]);
  assign tmp_2_lpi_4_dfm_mx0c1 = (~ mux_332_nl) & and_dcpl_164;
  assign or_302_nl = (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[2]) | (~
      and_dcpl_43);
  assign or_298_nl = (fsm_output[4:1]!=4'b0011);
  assign mux_234_nl = MUX_s_1_2_2(or_tmp_263, or_298_nl, fsm_output[8]);
  assign mux_235_nl = MUX_s_1_2_2(or_302_nl, mux_234_nl, fsm_output[6]);
  assign and_178_m1c = (~ mux_235_nl) & and_dcpl_52 & and_dcpl_20;
  assign nand_83_nl = ~((fsm_output[8]) & (fsm_output[4]) & (fsm_output[1]) & (fsm_output[3]));
  assign or_513_nl = (fsm_output[8]) | (fsm_output[4]) | (fsm_output[1]) | (fsm_output[3]);
  assign mux_102_nl = MUX_s_1_2_2(nand_83_nl, or_513_nl, fsm_output[5]);
  assign nor_220_nl = ~(mux_102_nl | (fsm_output[2]) | (fsm_output[0]) | (fsm_output[6])
      | (~ and_dcpl));
  assign nor_185_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[4])) | (fsm_output[2])
      | (~ (fsm_output[1])) | (fsm_output[3]));
  assign and_314_nl = (fsm_output[4:1]==4'b1011);
  assign nor_186_nl = ~((fsm_output[4:1]!=4'b1000));
  assign mux_103_nl = MUX_s_1_2_2(and_314_nl, nor_186_nl, fsm_output[8]);
  assign mux_104_nl = MUX_s_1_2_2(nor_185_nl, mux_103_nl, fsm_output[7]);
  assign nor_187_nl = ~((fsm_output[7]) | (fsm_output[8]) | (fsm_output[4]) | (~
      (fsm_output[2])) | (fsm_output[1]) | (~ (fsm_output[3])));
  assign mux_105_nl = MUX_s_1_2_2(mux_104_nl, nor_187_nl, fsm_output[9]);
  assign and_65_nl = mux_105_nl & and_dcpl_52 & (~ (fsm_output[6]));
  assign nor_183_nl = ~((fsm_output[5]) | (~ (fsm_output[8])) | (~ (fsm_output[2]))
      | (fsm_output[1]) | (~ (fsm_output[3])));
  assign and_313_nl = (fsm_output[5]) & (~ mux_tmp_106);
  assign mux_107_nl = MUX_s_1_2_2(nor_183_nl, and_313_nl, fsm_output[7]);
  assign nor_184_nl = ~((fsm_output[7]) | (fsm_output[5]) | (fsm_output[8]) | (~
      (fsm_output[2])) | (~ (fsm_output[1])) | (fsm_output[3]));
  assign mux_108_nl = MUX_s_1_2_2(mux_107_nl, nor_184_nl, fsm_output[9]);
  assign and_67_nl = mux_108_nl & and_dcpl_33 & (~ (fsm_output[6]));
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_11_5_2(z_out_2, (z_out_1[12:2]), COMP_LOOP_acc_psp_1_sva,
      (COMP_LOOP_acc_10_cse_12_1_1_sva[11:1]), (COMP_LOOP_acc_1_cse_2_sva[11:1]),
      {COMP_LOOP_or_2_cse , COMP_LOOP_or_4_cse , nor_220_nl , and_65_nl , and_67_nl});
  assign vec_rsc_0_0_i_da_d_pff = COMP_LOOP_mux_1_itm_mx1;
  assign nor_177_nl = ~((fsm_output[0]) | (~ (fsm_output[3])) | (~ (fsm_output[1]))
      | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) | (fsm_output[9:7]!=3'b011));
  assign or_140_nl = (~ (fsm_output[1])) | (fsm_output[8]) | (~ (fsm_output[9]))
      | (fsm_output[7]);
  assign or_139_nl = (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[9]) | (fsm_output[7]);
  assign mux_113_nl = MUX_s_1_2_2(or_140_nl, or_139_nl, fsm_output[3]);
  assign nor_178_nl = ~((fsm_output[0]) | (COMP_LOOP_acc_1_cse_2_sva[0]) | mux_113_nl);
  assign mux_114_nl = MUX_s_1_2_2(nor_177_nl, nor_178_nl, fsm_output[2]);
  assign nand_69_nl = ~((fsm_output[4]) & mux_114_nl);
  assign or_505_nl = (fsm_output[0]) | (fsm_output[3]) | (fsm_output[1]) | (VEC_LOOP_j_1_12_0_sva_11_0[0])
      | (fsm_output[9:7]!=3'b001);
  assign or_506_nl = (~ (fsm_output[0])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[0])
      | (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_111_nl = MUX_s_1_2_2(or_505_nl, or_506_nl, fsm_output[2]);
  assign or_133_nl = (fsm_output[9:7]!=3'b011);
  assign or_131_nl = (fsm_output[9:7]!=3'b010);
  assign mux_109_nl = MUX_s_1_2_2(or_133_nl, or_131_nl, fsm_output[1]);
  assign or_507_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[0])
      | mux_109_nl;
  assign or_508_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[0])
      | (~ (fsm_output[1])) | (fsm_output[8]) | (fsm_output[9]) | (~ (fsm_output[7]));
  assign mux_110_nl = MUX_s_1_2_2(or_507_nl, or_508_nl, fsm_output[2]);
  assign mux_112_nl = MUX_s_1_2_2(mux_111_nl, mux_110_nl, fsm_output[4]);
  assign mux_115_nl = MUX_s_1_2_2(nand_69_nl, mux_112_nl, fsm_output[5]);
  assign vec_rsc_0_0_i_wea_d_pff = ~(mux_115_nl | (fsm_output[6]));
  assign nor_170_nl = ~((~ (fsm_output[1])) | (z_out_1[1]) | (~ (fsm_output[7])));
  assign nor_171_nl = ~((~ (fsm_output[1])) | (z_out_1[1]) | (fsm_output[7]));
  assign mux_120_nl = MUX_s_1_2_2(nor_170_nl, nor_171_nl, fsm_output[2]);
  assign and_311_nl = (fsm_output[3]) & mux_120_nl;
  assign nor_172_nl = ~((fsm_output[2:1]!=2'b10) | (z_out_1[1]) | (~ (fsm_output[7])));
  assign nor_173_nl = ~((fsm_output[2:1]!=2'b00) | (z_out_1[1]) | (fsm_output[7]));
  assign mux_119_nl = MUX_s_1_2_2(nor_172_nl, nor_173_nl, fsm_output[3]);
  assign mux_121_nl = MUX_s_1_2_2(and_311_nl, mux_119_nl, fsm_output[8]);
  assign and_310_nl = (fsm_output[6]) & mux_121_nl;
  assign nor_175_nl = ~((fsm_output[1]) | (~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[0]) | (~ (fsm_output[7])));
  assign nor_176_nl = ~((fsm_output[1]) | (VEC_LOOP_j_1_12_0_sva_11_0[0]) | (fsm_output[7]));
  assign mux_117_nl = MUX_s_1_2_2(nor_175_nl, nor_176_nl, fsm_output[2]);
  assign nand_6_nl = ~((fsm_output[3]) & mux_117_nl);
  assign nand_63_nl = ~((fsm_output[1]) & VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm
      & (~ (COMP_LOOP_acc_1_cse_2_sva[0])) & (fsm_output[7]));
  assign or_144_nl = (~ (fsm_output[1])) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) |
      (fsm_output[7]);
  assign mux_116_nl = MUX_s_1_2_2(nand_63_nl, or_144_nl, fsm_output[2]);
  assign or_147_nl = (fsm_output[3]) | mux_116_nl;
  assign mux_118_nl = MUX_s_1_2_2(nand_6_nl, or_147_nl, fsm_output[8]);
  assign nor_174_nl = ~((fsm_output[6]) | mux_118_nl);
  assign mux_122_nl = MUX_s_1_2_2(and_310_nl, nor_174_nl, fsm_output[4]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = mux_122_nl & and_dcpl_79;
  assign and_340_nl = (~ (fsm_output[0])) & (fsm_output[3]) & (fsm_output[1]) & (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      & (fsm_output[9:7]==3'b011);
  assign nor_163_nl = ~((~ (fsm_output[1])) | (fsm_output[8]) | (~ (fsm_output[9]))
      | (fsm_output[7]));
  assign nor_164_nl = ~((fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[9]) |
      (fsm_output[7]));
  assign mux_127_nl = MUX_s_1_2_2(nor_163_nl, nor_164_nl, fsm_output[3]);
  assign and_308_nl = (~((fsm_output[0]) | (~ (COMP_LOOP_acc_1_cse_2_sva[0])))) &
      mux_127_nl;
  assign mux_128_nl = MUX_s_1_2_2(and_340_nl, and_308_nl, fsm_output[2]);
  assign nand_67_nl = ~((fsm_output[4]) & mux_128_nl);
  assign or_502_nl = (fsm_output[0]) | (fsm_output[3]) | (fsm_output[1]) | (~ (VEC_LOOP_j_1_12_0_sva_11_0[0]))
      | (fsm_output[9:7]!=3'b001);
  assign or_503_nl = (~ (fsm_output[0])) | (~ (fsm_output[3])) | (~ (COMP_LOOP_acc_10_cse_12_1_1_sva[0]))
      | (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_125_nl = MUX_s_1_2_2(or_502_nl, or_503_nl, fsm_output[2]);
  assign nor_167_nl = ~((fsm_output[9:7]!=3'b011));
  assign nor_168_nl = ~((fsm_output[9:7]!=3'b010));
  assign mux_123_nl = MUX_s_1_2_2(nor_167_nl, nor_168_nl, fsm_output[1]);
  assign nand_68_nl = ~((~((~ (fsm_output[0])) | (fsm_output[3]) | (~ (COMP_LOOP_acc_10_cse_12_1_1_sva[0]))))
      & mux_123_nl);
  assign or_504_nl = (~ (fsm_output[0])) | (fsm_output[3]) | (~ (COMP_LOOP_acc_10_cse_12_1_1_sva[0]))
      | (~ (fsm_output[1])) | (fsm_output[8]) | (fsm_output[9]) | (~ (fsm_output[7]));
  assign mux_124_nl = MUX_s_1_2_2(nand_68_nl, or_504_nl, fsm_output[2]);
  assign mux_126_nl = MUX_s_1_2_2(mux_125_nl, mux_124_nl, fsm_output[4]);
  assign mux_129_nl = MUX_s_1_2_2(nand_67_nl, mux_126_nl, fsm_output[5]);
  assign vec_rsc_0_1_i_wea_d_pff = ~(mux_129_nl | (fsm_output[6]));
  assign and_306_nl = (fsm_output[1]) & (z_out_1[1]) & (fsm_output[7]);
  assign nor_156_nl = ~((~ (fsm_output[1])) | (~ (z_out_1[1])) | (fsm_output[7]));
  assign mux_134_nl = MUX_s_1_2_2(and_306_nl, nor_156_nl, fsm_output[2]);
  assign and_305_nl = (fsm_output[3]) & mux_134_nl;
  assign nor_157_nl = ~((fsm_output[2:1]!=2'b10) | (~((z_out_1[1]) & (fsm_output[7]))));
  assign nor_158_nl = ~((fsm_output[2:1]!=2'b00) | (~ (z_out_1[1])) | (fsm_output[7]));
  assign mux_133_nl = MUX_s_1_2_2(nor_157_nl, nor_158_nl, fsm_output[3]);
  assign mux_135_nl = MUX_s_1_2_2(and_305_nl, mux_133_nl, fsm_output[8]);
  assign and_304_nl = (fsm_output[6]) & mux_135_nl;
  assign nor_160_nl = ~((fsm_output[1]) | (~ VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm)
      | not_tmp_94);
  assign nor_161_nl = ~((fsm_output[1]) | (~ (VEC_LOOP_j_1_12_0_sva_11_0[0])) | (fsm_output[7]));
  assign mux_131_nl = MUX_s_1_2_2(nor_160_nl, nor_161_nl, fsm_output[2]);
  assign nand_12_nl = ~((fsm_output[3]) & mux_131_nl);
  assign or_172_nl = (~((fsm_output[1]) & VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm))
      | not_tmp_94;
  assign or_170_nl = (~ (fsm_output[1])) | (~ (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]))
      | (fsm_output[7]);
  assign mux_130_nl = MUX_s_1_2_2(or_172_nl, or_170_nl, fsm_output[2]);
  assign or_173_nl = (fsm_output[3]) | mux_130_nl;
  assign mux_132_nl = MUX_s_1_2_2(nand_12_nl, or_173_nl, fsm_output[8]);
  assign nor_159_nl = ~((fsm_output[6]) | mux_132_nl);
  assign mux_136_nl = MUX_s_1_2_2(and_304_nl, nor_159_nl, fsm_output[4]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = mux_136_nl & and_dcpl_79;
  assign nor_233_nl = ~((~ (fsm_output[8])) | (fsm_output[3]) | (~ (fsm_output[2])));
  assign nor_234_nl = ~((fsm_output[8]) | (~ (fsm_output[3])) | (fsm_output[2]));
  assign mux_365_nl = MUX_s_1_2_2(nor_233_nl, nor_234_nl, fsm_output[1]);
  assign and_dcpl_232 = mux_365_nl & (fsm_output[5]) & (fsm_output[6]) & (~ (fsm_output[4]))
      & (~ (fsm_output[9])) & (fsm_output[7]) & (~ (fsm_output[0]));
  assign or_nl = (fsm_output[7:2]!=6'b100010);
  assign or_532_nl = (fsm_output[7:2]!=6'b000001);
  assign mux_367_nl = MUX_s_1_2_2(or_nl, or_532_nl, fsm_output[8]);
  assign nor_232_nl = ~((fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[5]) |
      (fsm_output[4]) | (fsm_output[6]));
  assign and_466_nl = (fsm_output[2]) & (fsm_output[7]) & (fsm_output[5]) & (fsm_output[4])
      & (fsm_output[6]);
  assign mux_366_nl = MUX_s_1_2_2(nor_232_nl, and_466_nl, fsm_output[3]);
  assign nand_86_nl = ~((fsm_output[8]) & mux_366_nl);
  assign mux_368_nl = MUX_s_1_2_2(mux_367_nl, nand_86_nl, fsm_output[1]);
  assign and_dcpl_234 = ~(mux_368_nl | (fsm_output[9]) | (fsm_output[0]));
  assign and_dcpl_239 = (~ (fsm_output[6])) & (fsm_output[4]);
  assign and_dcpl_241 = mux_150_cse & and_dcpl_239 & (fsm_output[5]) & (~ (fsm_output[9]))
      & (~ (fsm_output[7])) & (fsm_output[2]) & (~ (fsm_output[0]));
  assign and_dcpl_242 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_244 = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]));
  assign and_dcpl_247 = ~((fsm_output[6]) | (fsm_output[4]));
  assign and_dcpl_249 = and_dcpl_247 & (~ (fsm_output[5])) & and_dcpl_20;
  assign and_dcpl_250 = and_dcpl_249 & and_dcpl_244 & and_dcpl_242;
  assign and_dcpl_253 = (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[8]));
  assign and_dcpl_255 = and_dcpl_249 & and_dcpl_253 & nor_140_cse;
  assign and_dcpl_256 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_261 = and_dcpl_202 & and_dcpl_253 & and_dcpl_256;
  assign and_dcpl_262 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_266 = and_dcpl_151 & (~ (fsm_output[9])) & (fsm_output[7]);
  assign and_dcpl_267 = and_dcpl_266 & and_dcpl_262 & (~ (fsm_output[8])) & and_dcpl_256;
  assign and_dcpl_270 = and_dcpl_202 & and_dcpl_262 & (fsm_output[8]) & nor_140_cse;
  assign and_dcpl_272 = (fsm_output[2]) & (~ (fsm_output[3])) & (fsm_output[8]);
  assign and_dcpl_274 = and_dcpl_266 & and_dcpl_272 & nor_140_cse;
  assign and_dcpl_276 = and_dcpl_239 & (fsm_output[5]);
  assign and_dcpl_278 = and_dcpl_276 & and_dcpl_20 & and_dcpl_272 & and_dcpl_242;
  assign and_dcpl_281 = (fsm_output[9]) & (~ (fsm_output[7]));
  assign and_dcpl_284 = and_dcpl_247 & (fsm_output[5]) & and_dcpl_281 & and_dcpl_253
      & (fsm_output[1:0]==2'b11);
  assign and_dcpl_287 = and_dcpl_276 & and_dcpl_281 & and_dcpl_244 & nor_140_cse;
  assign nor_224_nl = ~((~ (fsm_output[8])) | (fsm_output[2]));
  assign nor_225_nl = ~((fsm_output[8]) | (~ (fsm_output[2])));
  assign mux_372_cse = MUX_s_1_2_2(nor_224_nl, nor_225_nl, fsm_output[1]);
  assign and_dcpl_343 = mux_372_cse & (~ (fsm_output[6])) & (fsm_output[4]) & (fsm_output[5])
      & (~ (fsm_output[9])) & (~ (fsm_output[7])) & (fsm_output[3]) & (~ (fsm_output[0]));
  assign or_537_nl = (fsm_output[0]) | (~((fsm_output[7:6]==2'b11)));
  assign or_536_nl = (~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[7]);
  assign mux_tmp = MUX_s_1_2_2(or_537_nl, or_536_nl, fsm_output[4]);
  assign COMP_LOOP_nor_3_itm = ~(and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287);
  assign COMP_LOOP_or_23_itm = and_dcpl_261 | and_dcpl_267;
  assign COMP_LOOP_or_24_itm = and_dcpl_270 | and_dcpl_274;
  always @(posedge clk) begin
    if ( ~ not_tmp_63 ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_26 & and_dcpl_24 & and_dcpl_23) | STAGE_LOOP_i_3_0_sva_mx0c1 )
        begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, (z_out_4[3:0]), STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ not_tmp_63 ) begin
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_1_obj_ld_cse <= 1'b0;
      modExp_exp_1_0_1_sva <= 1'b0;
      modExp_while_and_itm <= 1'b0;
      modExp_while_and_1_itm <= 1'b0;
      modExp_exp_1_1_1_sva <= 1'b0;
      modExp_exp_1_7_1_sva <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_1_obj_ld_cse <= and_dcpl_26 & and_dcpl_33 & (fsm_output[9:5]==5'b10001)
          & (~ (z_out_1[2]));
      modExp_exp_1_0_1_sva <= (COMP_LOOP_mux1h_13_nl & (~ and_dcpl_190)) | and_dcpl_194;
      modExp_while_and_itm <= (~ (modulo_result_rem_cmp_z[63])) & modExp_exp_1_0_1_sva;
      modExp_while_and_1_itm <= (modulo_result_rem_cmp_z[63]) & modExp_exp_1_0_1_sva;
      modExp_exp_1_1_1_sva <= COMP_LOOP_mux1h_23_nl & (~(and_dcpl_189 & and_dcpl_202));
      modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_40_nl & (~(and_dcpl_193 & and_dcpl_152));
    end
  end
  always @(posedge clk) begin
    modulo_result_rem_cmp_a <= MUX1HOT_v_64_20_2(modulo_result_rem_cmp_a_mx0w0, modExp_while_if_mul_mut,
        modExp_while_mul_itm, VEC_LOOP_1_COMP_LOOP_1_mul_mut_1, VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_if_mul_mut,
        VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_mul_itm, VEC_LOOP_1_COMP_LOOP_1_mul_mut,
        VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w7, COMP_LOOP_mux_1_itm, VEC_LOOP_1_COMP_LOOP_1_acc_8_itm,
        modExp_while_mul_itm_mx0w10, VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_mul_mut,
        VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_if_mul_itm, VEC_LOOP_1_COMP_LOOP_2_mul_mut,
        VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_if_mul_mut, VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_mul_itm,
        VEC_LOOP_2_COMP_LOOP_1_mul_mut, VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_mul_mut,
        VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_if_mul_itm, VEC_LOOP_2_COMP_LOOP_2_mul_mut,
        {and_dcpl_91 , and_105_nl , and_106_nl , and_107_nl , and_111_nl , and_114_nl
        , nor_218_nl , and_dcpl_106 , mux_160_nl , nor_208_nl , and_dcpl_111 , and_128_nl
        , and_130_nl , nor_214_nl , and_135_nl , and_138_nl , and_141_nl , and_145_nl
        , and_147_nl , and_148_nl});
    modulo_result_rem_cmp_b <= p_sva;
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_1, operator_64_false_acc_mut,
        and_dcpl_136);
    reg_operator_66_true_div_cmp_b_reg <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_136);
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_132_nl, or_tmp_207, fsm_output[9]) ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_acc_mut <= 65'b00000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( operator_64_false_acc_mut_mx0c0 | and_dcpl_144 | (~ mux_195_itm) )
        begin
      operator_64_false_acc_mut <= MUX1HOT_v_65_3_2(z_out_1, ({2'b00 , operator_64_false_slc_modExp_exp_63_1_3}),
          ({1'b0 , modulo_result_rem_cmp_z}), {operator_64_false_acc_mut_mx0c0 ,
          and_dcpl_144 , (~ mux_195_itm)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_1_12_0_sva_11_0 <= 12'b000000000000;
    end
    else if ( and_dcpl_144 | VEC_LOOP_j_1_12_0_sva_11_0_mx0c1 ) begin
      VEC_LOOP_j_1_12_0_sva_11_0 <= MUX_v_12_2_2(12'b000000000000, (z_out_1[11:0]),
          VEC_LOOP_j_1_12_0_sva_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_k_9_1_1_sva_7_0 <= 8'b00000000;
    end
    else if ( MUX_s_1_2_2(and_nl, nor_251_nl, fsm_output[8]) ) begin
      COMP_LOOP_k_9_1_1_sva_7_0 <= MUX_v_8_2_2(8'b00000000, (z_out_4[7:0]), nand_85_nl);
    end
  end
  always @(posedge clk) begin
    if ( (modExp_exp_1_0_1_sva | modExp_while_and_itm | modExp_while_and_1_itm |
        modExp_result_sva_mx0c0 | (~ mux_233_nl)) & (modExp_result_sva_mx0c0 | modExp_result_and_rgt
        | modExp_result_and_1_rgt) ) begin
      modExp_result_sva <= MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          (operator_64_false_acc_mut[63:0]), modulo_qr_sva_1_mx0w8, {modExp_result_sva_mx0c0
          , modExp_result_and_rgt , modExp_result_and_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_253_nl, or_534_nl, fsm_output[9]) ) begin
      COMP_LOOP_mux_1_itm <= MUX1HOT_v_64_7_2(r_sva, (operator_64_false_acc_mut[63:0]),
          modulo_qr_sva_1_mx0w8, modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
          VEC_LOOP_1_COMP_LOOP_1_acc_5_mut_mx0w7, {and_176_nl , r_or_nl , r_or_1_nl
          , and_dcpl_166 , and_189_nl , and_193_nl , and_dcpl_106});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_1_COMP_LOOP_1_acc_8_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( (modExp_exp_1_0_1_sva | and_dcpl_144 | and_dcpl_166 | and_dcpl_106)
        & mux_289_nl ) begin
      VEC_LOOP_1_COMP_LOOP_1_acc_8_itm <= MUX1HOT_v_64_5_2(({1'b0 , operator_64_false_slc_modExp_exp_63_1_3}),
          64'b0000000000000000000000000000000000000000000000000000000000000001, (operator_64_false_acc_mut[63:0]),
          modulo_qr_sva_1_mx0w8, (z_out_1[63:0]), {and_dcpl_144 , and_dcpl_166 ,
          COMP_LOOP_and_nl , COMP_LOOP_and_1_nl , and_dcpl_106});
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_303_nl & and_dcpl_93) ) begin
      modExp_while_if_mul_mut <= modulo_result_rem_cmp_a_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva <= 1'b0;
    end
    else if ( and_dcpl_91 | and_dcpl_198 | and_dcpl_153 ) begin
      exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva <= MUX1HOT_s_1_3_2((~ (z_out_1[63])),
          (~ z_out_5_8), (~ (readslicef_10_1_9(VEC_LOOP_1_COMP_LOOP_1_acc_11_nl))),
          {and_dcpl_91 , and_dcpl_198 , and_dcpl_153});
    end
  end
  always @(posedge clk) begin
    if ( ~(or_dcpl_44 | (~ (fsm_output[0])) | (fsm_output[4]) | (fsm_output[8]) |
        (fsm_output[5]) | (fsm_output[6]) | or_dcpl_39) ) begin
      modExp_while_mul_itm <= modExp_while_mul_itm_mx0w10;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_or_2_cse ) begin
      COMP_LOOP_acc_psp_1_sva <= z_out_2;
    end
  end
  always @(posedge clk) begin
    if ( VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c0
        | VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c1
        | and_dcpl_111 ) begin
      VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm
          <= MUX1HOT_s_1_3_2((z_out_1[9]), (z_out[9]), z_out_5_8, {VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c0
          , VEC_LOOP_1_COMP_LOOP_1_operator_64_false_1_slc_operator_64_false_1_acc_9_1_itm_mx0c1
          , and_dcpl_111});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_320, mux_324_nl, fsm_output[4]) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= nl_COMP_LOOP_acc_1_cse_2_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( ((~ mux_329_nl) & and_dcpl_164) | tmp_2_lpi_4_dfm_mx0c1 ) begin
      tmp_2_lpi_4_dfm <= MUX_v_64_2_2(vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, tmp_2_lpi_4_dfm_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_0_1_sva_1 <= 1'b0;
    end
    else if ( ~(mux_340_nl & (~ (fsm_output[9]))) ) begin
      modExp_exp_1_0_1_sva_1 <= MUX_s_1_2_2((COMP_LOOP_k_9_1_1_sva_7_0[0]), modExp_exp_1_1_1_sva,
          and_230_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_2_1_sva <= 1'b0;
    end
    else if ( ~ and_dcpl_214 ) begin
      modExp_exp_1_2_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[1]), modExp_exp_1_3_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[2]), {and_dcpl_190 , and_dcpl_211 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_3_1_sva <= 1'b0;
    end
    else if ( ~ and_dcpl_214 ) begin
      modExp_exp_1_3_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[2]), modExp_exp_1_4_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[3]), {and_dcpl_190 , and_dcpl_211 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_4_1_sva <= 1'b0;
    end
    else if ( ~ and_dcpl_214 ) begin
      modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[3]), modExp_exp_1_5_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[4]), {and_dcpl_190 , and_dcpl_211 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_5_1_sva <= 1'b0;
    end
    else if ( ~ and_dcpl_214 ) begin
      modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[4]), modExp_exp_1_6_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[5]), {and_dcpl_190 , and_dcpl_211 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_6_1_sva <= 1'b0;
    end
    else if ( ~ and_dcpl_214 ) begin
      modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_1_1_sva_7_0[5]), modExp_exp_1_7_1_sva,
          (COMP_LOOP_k_9_1_1_sva_7_0[6]), {and_dcpl_190 , and_dcpl_211 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( ~((~ mux_361_nl) & and_dcpl_98) ) begin
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_if_mul_mut <= VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~((~ and_dcpl_44) | or_dcpl_58 | or_dcpl_63 | or_dcpl_39) ) begin
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_mul_itm <= modExp_while_mul_itm_mx0w10;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= 12'b000000000000;
    end
    else if ( COMP_LOOP_or_4_cse ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_1[12:1];
    end
  end
  always @(posedge clk) begin
    if ( ~(or_25_cse | (fsm_output[0]) | (~ (fsm_output[4])) | or_dcpl_72 | or_dcpl_39)
        ) begin
      VEC_LOOP_1_COMP_LOOP_1_mul_mut <= VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_273 | or_dcpl_63 | or_tmp_52) ) begin
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_mul_mut <= modExp_while_mul_itm_mx0w10;
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_362_nl & and_dcpl_113) ) begin
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_if_mul_itm <= VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_279 | or_dcpl_72 | or_tmp_52) ) begin
      VEC_LOOP_1_COMP_LOOP_2_mul_mut <= VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~((~ mux_363_nl) & and_dcpl_119) ) begin
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_if_mul_mut <= VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_89_cse | or_dcpl_58 | or_dcpl_84) ) begin
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_mul_itm <= modExp_while_mul_itm_mx0w10;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_189 | or_dcpl_68 | or_dcpl_89 | or_dcpl_39) ) begin
      VEC_LOOP_2_COMP_LOOP_1_mul_mut <= VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_tmp_271 | or_dcpl_83 | or_tmp_52) ) begin
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_mul_mut <= modExp_while_mul_itm_mx0w10;
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_364_nl & and_dcpl_127) ) begin
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_if_mul_itm <= VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_52_cse | or_dcpl_68 | or_dcpl_89 | or_tmp_52) ) begin
      VEC_LOOP_2_COMP_LOOP_2_mul_mut <= VEC_LOOP_1_COMP_LOOP_1_mul_mut_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_VEC_LOOP_1_acc_1_psp_ftd_1 <= 12'b000000000000;
    end
    else if ( ~(or_tmp_11 | or_dcpl_58 | or_dcpl_84) ) begin
      reg_VEC_LOOP_1_acc_1_psp_ftd_1 <= z_out_1[11:0];
    end
  end
  assign nor_nl = ~((fsm_output[4]) | mux_tmp_137);
  assign mux_139_nl = MUX_s_1_2_2(or_tmp_154, nor_nl, fsm_output[5]);
  assign and_105_nl = mux_139_nl & and_dcpl_93;
  assign mux_140_nl = MUX_s_1_2_2(mux_tmp_137, (~ nor_tmp_1), fsm_output[4]);
  assign and_106_nl = mux_140_nl & and_dcpl_36;
  assign and_300_nl = (fsm_output[8]) & (fsm_output[1]) & (fsm_output[7]) & (fsm_output[2]);
  assign nor_152_nl = ~((fsm_output[8]) | (fsm_output[1]) | (fsm_output[7]) | (fsm_output[2]));
  assign mux_144_nl = MUX_s_1_2_2(and_300_nl, nor_152_nl, fsm_output[4]);
  assign and_299_nl = (fsm_output[6]) & mux_144_nl;
  assign nor_153_nl = ~((~ (fsm_output[1])) | (fsm_output[7]) | (~ (fsm_output[2])));
  assign nor_154_nl = ~((fsm_output[1]) | (fsm_output[7]) | (fsm_output[2]));
  assign mux_142_nl = MUX_s_1_2_2(nor_153_nl, nor_154_nl, fsm_output[8]);
  assign and_301_nl = (fsm_output[4]) & mux_142_nl;
  assign or_188_nl = (fsm_output[1]) | (~((fsm_output[7]) & (fsm_output[2])));
  assign or_187_nl = (~ (fsm_output[1])) | (fsm_output[7]) | (fsm_output[2]);
  assign mux_141_nl = MUX_s_1_2_2(or_188_nl, or_187_nl, fsm_output[8]);
  assign nor_155_nl = ~((fsm_output[4]) | mux_141_nl);
  assign mux_143_nl = MUX_s_1_2_2(and_301_nl, nor_155_nl, fsm_output[6]);
  assign mux_145_nl = MUX_s_1_2_2(and_299_nl, mux_143_nl, fsm_output[3]);
  assign and_107_nl = mux_145_nl & and_dcpl_79;
  assign or_195_nl = (fsm_output[5]) | and_tmp_11;
  assign mux_147_nl = MUX_s_1_2_2(not_tmp_111, or_195_nl, fsm_output[6]);
  assign and_111_nl = (~ mux_147_nl) & and_dcpl_98;
  assign nor_151_nl = ~((fsm_output[4]) | nor_tmp_2);
  assign mux_148_nl = MUX_s_1_2_2(and_tmp_11, nor_151_nl, fsm_output[5]);
  assign and_114_nl = mux_148_nl & and_dcpl_100 & and_dcpl_20;
  assign nand_80_nl = ~((fsm_output[6:4]==3'b111) & or_100_cse);
  assign or_512_nl = (fsm_output[6:4]!=3'b000) | or_tmp_167;
  assign mux_149_nl = MUX_s_1_2_2(nand_80_nl, or_512_nl, fsm_output[7]);
  assign nor_218_nl = ~(mux_149_nl | (fsm_output[9:8]!=2'b00));
  assign mux_158_nl = MUX_s_1_2_2((~ mux_tmp_146), mux_tmp_157, fsm_output[4]);
  assign nor_144_nl = ~((fsm_output[6]) | (fsm_output[5]) | (~ (fsm_output[8])) |
      mux_158_nl);
  assign mux_154_nl = MUX_s_1_2_2((~ nor_tmp_38), and_334_cse, fsm_output[4]);
  assign mux_153_nl = MUX_s_1_2_2((~ mux_tmp_137), nor_tmp_38, fsm_output[4]);
  assign mux_155_nl = MUX_s_1_2_2(mux_154_nl, mux_153_nl, fsm_output[8]);
  assign nor_145_nl = ~((fsm_output[5]) | mux_155_nl);
  assign and_292_nl = (fsm_output[5]) & (fsm_output[8]) & (fsm_output[4]) & (fsm_output[0])
      & (fsm_output[2]) & (fsm_output[1]) & (fsm_output[3]);
  assign mux_156_nl = MUX_s_1_2_2(nor_145_nl, and_292_nl, fsm_output[6]);
  assign mux_159_nl = MUX_s_1_2_2(nor_144_nl, mux_156_nl, fsm_output[7]);
  assign nor_146_nl = ~((fsm_output[8:5]!=4'b0000) | and_tmp_11);
  assign mux_160_nl = MUX_s_1_2_2(mux_159_nl, nor_146_nl, fsm_output[9]);
  assign mux_168_nl = MUX_s_1_2_2(or_74_cse, (~ or_74_cse), fsm_output[9]);
  assign nand_64_nl = ~((fsm_output[5]) & mux_168_nl);
  assign nor_209_nl = ~((fsm_output[8]) | (fsm_output[2]) | (fsm_output[7]));
  assign mux_167_nl = MUX_s_1_2_2(or_74_cse, nor_209_nl, fsm_output[9]);
  assign nand_65_nl = ~((fsm_output[5]) & mux_167_nl);
  assign mux_169_nl = MUX_s_1_2_2(nand_64_nl, nand_65_nl, fsm_output[3]);
  assign nand_66_nl = ~((~((~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[2]))))
      & (~(nor_140_cse | (fsm_output[7]))));
  assign nand_50_nl = ~(nand_51_cse & (fsm_output[7]));
  assign or_213_nl = (fsm_output[2]) | (fsm_output[1]) | (fsm_output[7]);
  assign mux_164_nl = MUX_s_1_2_2(nand_50_nl, or_213_nl, fsm_output[8]);
  assign or_500_nl = (fsm_output[9]) | mux_164_nl;
  assign mux_165_nl = MUX_s_1_2_2(nand_66_nl, or_500_nl, fsm_output[5]);
  assign nand_52_nl = ~((fsm_output[2]) & (fsm_output[0]) & (fsm_output[1]) & (fsm_output[7]));
  assign and_291_nl = (fsm_output[1]) & (fsm_output[7]);
  assign mux_161_nl = MUX_s_1_2_2(and_291_nl, or_210_cse, fsm_output[0]);
  assign nor_143_nl = ~((fsm_output[2]) | mux_161_nl);
  assign mux_162_nl = MUX_s_1_2_2(nand_52_nl, nor_143_nl, fsm_output[8]);
  assign mux_163_nl = MUX_s_1_2_2(mux_162_nl, or_74_cse, fsm_output[9]);
  assign or_501_nl = (fsm_output[5]) | mux_163_nl;
  assign mux_166_nl = MUX_s_1_2_2(mux_165_nl, or_501_nl, fsm_output[3]);
  assign mux_170_nl = MUX_s_1_2_2(mux_169_nl, mux_166_nl, fsm_output[4]);
  assign nor_208_nl = ~(mux_170_nl | (fsm_output[6]));
  assign and_287_nl = (fsm_output[5:4]==2'b11) & mux_tmp_157;
  assign nor_138_nl = ~((fsm_output[5]) | and_tmp_10);
  assign mux_172_nl = MUX_s_1_2_2(and_287_nl, nor_138_nl, fsm_output[6]);
  assign and_128_nl = mux_172_nl & and_dcpl_113;
  assign nor_137_nl = ~((fsm_output[4:3]!=2'b00));
  assign mux_173_nl = MUX_s_1_2_2(and_tmp_10, nor_137_nl, fsm_output[5]);
  assign and_130_nl = mux_173_nl & and_dcpl_100 & and_dcpl;
  assign or_509_nl = (fsm_output[6]) | (fsm_output[5]) | (~ (fsm_output[8])) | (fsm_output[4])
      | mux_tmp_137;
  assign nand_73_nl = ~((fsm_output[6]) & (fsm_output[5]) & (~ (fsm_output[8])) &
      or_tmp_154);
  assign mux_174_nl = MUX_s_1_2_2(or_509_nl, nand_73_nl, fsm_output[7]);
  assign nor_214_nl = ~(mux_174_nl | (fsm_output[9]));
  assign or_228_nl = (fsm_output[5:4]!=2'b00) | and_334_cse;
  assign mux_175_nl = MUX_s_1_2_2(not_tmp_141, or_228_nl, fsm_output[6]);
  assign and_135_nl = (~ mux_175_nl) & and_dcpl_119;
  assign or_493_nl = (fsm_output[4]) | and_334_cse;
  assign nor_135_nl = ~((fsm_output[4]) | or_tmp_19);
  assign mux_176_nl = MUX_s_1_2_2(or_493_nl, nor_135_nl, fsm_output[5]);
  assign and_138_nl = mux_176_nl & and_dcpl_121 & and_dcpl_20;
  assign and_285_nl = (fsm_output[6:5]==2'b11) & or_tmp_201;
  assign nor_134_nl = ~((fsm_output[6:0]!=7'b0000000));
  assign mux_177_nl = MUX_s_1_2_2(and_285_nl, nor_134_nl, fsm_output[7]);
  assign and_141_nl = mux_177_nl & (fsm_output[9:8]==2'b01);
  assign and_284_nl = (fsm_output[5:4]==2'b11) & mux_tmp_146;
  assign nor_133_nl = ~((fsm_output[5:4]!=2'b00) | mux_tmp_157);
  assign mux_178_nl = MUX_s_1_2_2(and_284_nl, nor_133_nl, fsm_output[6]);
  assign and_145_nl = mux_178_nl & and_dcpl_127;
  assign mux_179_nl = MUX_s_1_2_2(or_tmp_201, (~ or_tmp_204), fsm_output[5]);
  assign and_147_nl = mux_179_nl & and_dcpl_121 & and_dcpl;
  assign mux_180_nl = MUX_s_1_2_2(or_tmp_167, (~ mux_tmp_138), fsm_output[4]);
  assign and_148_nl = mux_180_nl & and_dcpl_73;
  assign COMP_LOOP_and_5_nl = (~ and_dcpl_157) & and_dcpl_144;
  assign nor_113_nl = ~((~ (fsm_output[3])) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[8]));
  assign nor_114_nl = ~((fsm_output[3]) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[8]));
  assign mux_300_nl = MUX_s_1_2_2(nor_113_nl, nor_114_nl, fsm_output[5]);
  assign nor_115_nl = ~((fsm_output[8:7]!=2'b00));
  assign mux_299_nl = MUX_s_1_2_2(nor_115_nl, mux_tmp_296, fsm_output[5]);
  assign mux_301_nl = MUX_s_1_2_2(mux_300_nl, mux_299_nl, fsm_output[4]);
  assign and_270_nl = or_492_cse & (fsm_output[8:7]==2'b11);
  assign or_344_nl = and_271_cse | (fsm_output[8:7]!=2'b00);
  assign mux_294_nl = MUX_s_1_2_2(and_270_nl, or_344_nl, fsm_output[3]);
  assign mux_297_nl = MUX_s_1_2_2(mux_tmp_296, mux_294_nl, fsm_output[0]);
  assign nand_48_nl = ~((fsm_output[5]) & mux_297_nl);
  assign or_341_nl = (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[8]));
  assign or_339_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[8]);
  assign mux_293_nl = MUX_s_1_2_2(or_341_nl, or_339_nl, fsm_output[1]);
  assign nor_116_nl = ~((fsm_output[5]) | (~((fsm_output[0]) | (fsm_output[3]) |
      mux_293_nl)));
  assign mux_298_nl = MUX_s_1_2_2(nand_48_nl, nor_116_nl, fsm_output[4]);
  assign mux_302_nl = MUX_s_1_2_2(mux_301_nl, mux_298_nl, fsm_output[6]);
  assign and_212_nl = mux_302_nl & (~ (fsm_output[9]));
  assign COMP_LOOP_mux1h_13_nl = MUX1HOT_s_1_4_2((operator_66_true_div_cmp_z_oreg[0]),
      (VEC_LOOP_1_COMP_LOOP_1_acc_8_itm[0]), modExp_exp_1_0_1_sva_1, modExp_exp_1_0_1_sva,
      {COMP_LOOP_and_5_nl , and_dcpl_157 , and_dcpl_186 , and_212_nl});
  assign and_257_nl = or_492_cse & (fsm_output[7]) & (fsm_output[4]) & (fsm_output[5]);
  assign and_258_nl = ((fsm_output[2]) | (fsm_output[7])) & (fsm_output[5:4]==2'b11);
  assign mux_350_nl = MUX_s_1_2_2(nor_tmp_81, and_258_nl, fsm_output[1]);
  assign mux_351_nl = MUX_s_1_2_2(and_257_nl, mux_350_nl, fsm_output[0]);
  assign nand_42_nl = ~((fsm_output[3]) & mux_351_nl);
  assign mux_348_nl = MUX_s_1_2_2(nor_tmp_79, nor_tmp_77, or_71_cse);
  assign mux_349_nl = MUX_s_1_2_2(and_259_cse, mux_348_nl, fsm_output[3]);
  assign mux_352_nl = MUX_s_1_2_2(nand_42_nl, mux_349_nl, fsm_output[6]);
  assign and_260_nl = ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[7]))
      & (fsm_output[5:4]==2'b11);
  assign mux_346_nl = MUX_s_1_2_2(nor_tmp_81, and_260_nl, fsm_output[3]);
  assign mux_344_nl = MUX_s_1_2_2(nor_tmp_79, nor_tmp_77, and_282_cse);
  assign mux_345_nl = MUX_s_1_2_2(mux_344_nl, (fsm_output[5]), fsm_output[3]);
  assign mux_347_nl = MUX_s_1_2_2((~ mux_346_nl), mux_345_nl, fsm_output[6]);
  assign mux_353_nl = MUX_s_1_2_2(mux_352_nl, mux_347_nl, fsm_output[8]);
  assign nor_213_nl = ~(mux_353_nl | (fsm_output[9]));
  assign COMP_LOOP_mux1h_23_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_1_1_sva_7_0[7]),
      modExp_exp_1_2_1_sva, modExp_exp_1_1_1_sva, (COMP_LOOP_k_9_1_1_sva_7_0[1]),
      {and_dcpl_190 , and_dcpl_211 , nor_213_nl , and_dcpl_194});
  assign COMP_LOOP_mux1h_40_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_1_1_sva_7_0[6]),
      modExp_exp_1_1_1_sva, modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_1_1_sva_7_0[7]),
      {and_dcpl_190 , and_dcpl_198 , and_dcpl_214 , and_dcpl_194});
  assign nor_132_nl = ~((fsm_output[8:1]!=8'b00000000));
  assign nor_128_nl = ~((fsm_output[8]) | (fsm_output[4]) | (fsm_output[2]) | (~
      and_dcpl_43));
  assign nor_129_nl = ~((~ (fsm_output[4])) | (fsm_output[2]) | (~ and_dcpl_43));
  assign nor_130_nl = ~((fsm_output[4:1]!=4'b1010));
  assign mux_216_nl = MUX_s_1_2_2(nor_129_nl, nor_130_nl, fsm_output[8]);
  assign mux_217_nl = MUX_s_1_2_2(nor_128_nl, mux_216_nl, fsm_output[5]);
  assign nor_131_nl = ~((~ (fsm_output[5])) | (fsm_output[8]) | (fsm_output[4]) |
      (~ and_dcpl_44));
  assign mux_218_nl = MUX_s_1_2_2(mux_217_nl, nor_131_nl, fsm_output[9]);
  assign nand_85_nl = ~(mux_218_nl & (fsm_output[0]) & (~ (fsm_output[6])) & (~ (fsm_output[7])));
  assign nor_248_nl = ~((fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[0])) |
      (fsm_output[6]) | (fsm_output[7]));
  assign nor_249_nl = ~((fsm_output[9]) | mux_tmp);
  assign mux_374_nl = MUX_s_1_2_2(nor_248_nl, nor_249_nl, fsm_output[5]);
  assign nor_250_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[9])) | (fsm_output[4])
      | (~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[7]));
  assign mux_375_nl = MUX_s_1_2_2(mux_374_nl, nor_250_nl, fsm_output[2]);
  assign and_nl = (fsm_output[3]) & (fsm_output[1]) & mux_375_nl;
  assign nor_251_nl = ~((fsm_output[3]) | (fsm_output[1]) | (~ (fsm_output[2])) |
      (~ (fsm_output[5])) | (fsm_output[9]) | mux_tmp);
  assign or_296_nl = (fsm_output[8]) | (fsm_output[4]) | nor_tmp_2;
  assign or_294_nl = (fsm_output[8]) | (fsm_output[4]) | (fsm_output[0]) | (~ (fsm_output[2]))
      | (fsm_output[1]) | (fsm_output[3]);
  assign mux_232_nl = MUX_s_1_2_2(or_296_nl, or_294_nl, fsm_output[5]);
  assign nor_124_nl = ~((fsm_output[7:6]!=2'b00) | mux_232_nl);
  assign mux_233_nl = MUX_s_1_2_2(nor_124_nl, or_tmp_207, fsm_output[9]);
  assign and_176_nl = and_dcpl_58 & and_dcpl_137 & and_dcpl_23;
  assign r_or_nl = ((~ (operator_64_false_acc_mut[63])) & and_178_m1c) | (and_dcpl_181
      & and_dcpl_179 & (~ (fsm_output[9])) & (~ (operator_64_false_acc_mut[63])));
  assign r_or_1_nl = ((operator_64_false_acc_mut[63]) & and_178_m1c) | (and_dcpl_181
      & and_dcpl_179 & (~ (fsm_output[9])) & (operator_64_false_acc_mut[63]));
  assign and_189_nl = and_dcpl_171 & (~ (fsm_output[4])) & (~ (COMP_LOOP_acc_10_cse_12_1_1_sva[0]))
      & (fsm_output[5]) & and_dcpl_167;
  assign and_193_nl = and_dcpl_171 & (~ (fsm_output[4])) & (COMP_LOOP_acc_10_cse_12_1_1_sva[0])
      & (fsm_output[5]) & and_dcpl_167;
  assign mux_250_nl = MUX_s_1_2_2((~ mux_tmp_146), nor_tmp_1, fsm_output[4]);
  assign mux_251_nl = MUX_s_1_2_2(or_tmp_279, mux_250_nl, fsm_output[8]);
  assign or_314_nl = (~ (fsm_output[4])) | (fsm_output[0]) | (~ and_dcpl_44);
  assign or_312_nl = (fsm_output[4:0]!=5'b11000);
  assign mux_249_nl = MUX_s_1_2_2(or_314_nl, or_312_nl, fsm_output[8]);
  assign mux_252_nl = MUX_s_1_2_2(mux_251_nl, mux_249_nl, fsm_output[5]);
  assign or_533_nl = (fsm_output[6]) | mux_252_nl;
  assign mux_245_nl = MUX_s_1_2_2((~ nor_tmp_38), and_dcpl_44, fsm_output[4]);
  assign mux_244_nl = MUX_s_1_2_2((~ mux_tmp_137), (fsm_output[3]), fsm_output[4]);
  assign mux_246_nl = MUX_s_1_2_2(mux_245_nl, mux_244_nl, fsm_output[8]);
  assign mux_243_nl = MUX_s_1_2_2(or_tmp_273, or_tmp_271, fsm_output[8]);
  assign mux_247_nl = MUX_s_1_2_2(mux_246_nl, mux_243_nl, fsm_output[5]);
  assign and_195_nl = (fsm_output[4]) & mux_tmp_137;
  assign mux_241_nl = MUX_s_1_2_2(and_195_nl, or_tmp_154, fsm_output[8]);
  assign nor_122_nl = ~((fsm_output[4]) | nor_tmp_1);
  assign mux_239_nl = MUX_s_1_2_2((~ or_96_cse), and_334_cse, fsm_output[4]);
  assign mux_240_nl = MUX_s_1_2_2(nor_122_nl, mux_239_nl, fsm_output[8]);
  assign mux_242_nl = MUX_s_1_2_2(mux_241_nl, mux_240_nl, fsm_output[5]);
  assign mux_248_nl = MUX_s_1_2_2(mux_247_nl, (~ mux_242_nl), fsm_output[6]);
  assign mux_253_nl = MUX_s_1_2_2(or_533_nl, mux_248_nl, fsm_output[7]);
  assign or_534_nl = (fsm_output[8:5]!=4'b0000) | and_tmp_17;
  assign COMP_LOOP_and_nl = (~ modExp_1_while_and_11) & and_dcpl_186;
  assign COMP_LOOP_and_1_nl = modExp_1_while_and_11 & and_dcpl_186;
  assign mux_284_nl = MUX_s_1_2_2(mux_tmp_269, mux_tmp_263, and_282_cse);
  assign mux_282_nl = MUX_s_1_2_2(mux_tmp_263, and_tmp_19, fsm_output[0]);
  assign mux_283_nl = MUX_s_1_2_2(mux_282_nl, nor_tmp_57, fsm_output[1]);
  assign mux_285_nl = MUX_s_1_2_2(mux_284_nl, mux_283_nl, fsm_output[7]);
  assign mux_286_nl = MUX_s_1_2_2(mux_tmp_269, mux_285_nl, fsm_output[3]);
  assign mux_279_nl = MUX_s_1_2_2(mux_tmp_272, mux_tmp_263, or_71_cse);
  assign mux_278_nl = MUX_s_1_2_2(mux_tmp_263, and_tmp_19, and_282_cse);
  assign mux_280_nl = MUX_s_1_2_2(mux_279_nl, mux_278_nl, fsm_output[7]);
  assign mux_277_nl = MUX_s_1_2_2(nor_tmp_57, nor_tmp_56, or_210_cse);
  assign mux_281_nl = MUX_s_1_2_2(mux_280_nl, mux_277_nl, fsm_output[3]);
  assign mux_287_nl = MUX_s_1_2_2(mux_286_nl, mux_281_nl, fsm_output[8]);
  assign or_329_nl = (fsm_output[1:0]!=2'b10);
  assign mux_273_nl = MUX_s_1_2_2(mux_tmp_272, mux_tmp_269, or_329_nl);
  assign mux_270_nl = MUX_s_1_2_2(mux_tmp_269, mux_tmp_263, or_71_cse);
  assign mux_274_nl = MUX_s_1_2_2(mux_273_nl, mux_270_nl, fsm_output[7]);
  assign mux_267_nl = MUX_s_1_2_2(and_259_cse, nor_tmp_57, fsm_output[1]);
  assign mux_268_nl = MUX_s_1_2_2(mux_267_nl, nor_tmp_56, fsm_output[7]);
  assign mux_275_nl = MUX_s_1_2_2(mux_274_nl, mux_268_nl, fsm_output[3]);
  assign mux_264_nl = MUX_s_1_2_2(mux_tmp_263, and_259_cse, or_71_cse);
  assign mux_262_nl = MUX_s_1_2_2(nor_tmp_57, nor_tmp_56, fsm_output[1]);
  assign mux_265_nl = MUX_s_1_2_2(mux_264_nl, mux_262_nl, fsm_output[7]);
  assign nor_120_nl = ~((fsm_output[5:4]!=2'b10));
  assign and_276_nl = (fsm_output[7]) & (fsm_output[1]) & (fsm_output[0]);
  assign mux_261_nl = MUX_s_1_2_2(nor_tmp_56, nor_120_nl, and_276_nl);
  assign mux_266_nl = MUX_s_1_2_2(mux_265_nl, mux_261_nl, fsm_output[3]);
  assign mux_276_nl = MUX_s_1_2_2(mux_275_nl, mux_266_nl, fsm_output[8]);
  assign mux_288_nl = MUX_s_1_2_2(mux_287_nl, mux_276_nl, fsm_output[2]);
  assign or_323_nl = (fsm_output[6:5]!=2'b00);
  assign mux_258_nl = MUX_s_1_2_2(mux_tmp_256, or_323_nl, and_282_cse);
  assign or_324_nl = (fsm_output[7]) | mux_258_nl;
  assign mux_259_nl = MUX_s_1_2_2(or_tmp_284, or_324_nl, fsm_output[3]);
  assign or_325_nl = (fsm_output[8]) | mux_259_nl;
  assign or_319_nl = (fsm_output[7:5]!=3'b000);
  assign mux_257_nl = MUX_s_1_2_2(or_tmp_284, or_319_nl, fsm_output[3]);
  assign or_322_nl = (fsm_output[8]) | mux_257_nl;
  assign mux_260_nl = MUX_s_1_2_2(or_325_nl, or_322_nl, fsm_output[2]);
  assign mux_289_nl = MUX_s_1_2_2(mux_288_nl, mux_260_nl, fsm_output[9]);
  assign mux_303_nl = MUX_s_1_2_2(or_tmp_154, (~ or_tmp_204), fsm_output[5]);
  assign nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl = ({z_out_4 , 1'b0}) + ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))})
      + 10'b0000000001;
  assign VEC_LOOP_1_COMP_LOOP_1_acc_11_nl = nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl[9:0];
  assign COMP_LOOP_mux_21_nl = MUX_v_12_2_2(VEC_LOOP_j_1_12_0_sva_11_0, reg_VEC_LOOP_1_acc_1_psp_ftd_1,
      and_468_cse);
  assign nl_COMP_LOOP_acc_1_cse_2_sva  = COMP_LOOP_mux_21_nl + conv_u2u_9_12({COMP_LOOP_k_9_1_1_sva_7_0
      , 1'b1});
  assign mux_323_nl = MUX_s_1_2_2(mux_tmp_320, or_tmp_337, fsm_output[3]);
  assign mux_317_nl = MUX_s_1_2_2(or_tmp_335, or_tmp_337, fsm_output[5]);
  assign mux_318_nl = MUX_s_1_2_2(mux_317_nl, mux_tmp_314, fsm_output[0]);
  assign mux_321_nl = MUX_s_1_2_2(mux_tmp_320, mux_318_nl, fsm_output[3]);
  assign nor_70_nl = ~((fsm_output[0]) | (~ (fsm_output[5])));
  assign mux_315_nl = MUX_s_1_2_2(or_tmp_337, or_tmp_335, nor_70_nl);
  assign mux_316_nl = MUX_s_1_2_2(mux_315_nl, mux_tmp_314, fsm_output[3]);
  assign mux_322_nl = MUX_s_1_2_2(mux_321_nl, mux_316_nl, fsm_output[1]);
  assign mux_324_nl = MUX_s_1_2_2(mux_323_nl, mux_322_nl, fsm_output[2]);
  assign mux_327_nl = MUX_s_1_2_2(mux_tmp_326, or_tmp_341, VEC_LOOP_j_1_12_0_sva_11_0[0]);
  assign or_396_nl = (VEC_LOOP_j_1_12_0_sva_11_0[0]) | (fsm_output[8]) | (~ (fsm_output[2]))
      | (fsm_output[1]) | (~ (fsm_output[3]));
  assign mux_328_nl = MUX_s_1_2_2(mux_327_nl, or_396_nl, reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]);
  assign or_394_nl = (COMP_LOOP_acc_1_cse_2_sva[0]) | mux_tmp_106;
  assign mux_329_nl = MUX_s_1_2_2(mux_328_nl, or_394_nl, fsm_output[7]);
  assign and_230_nl = and_dcpl_165 & and_dcpl_137 & (fsm_output[5]) & and_dcpl_167;
  assign and_341_nl = (~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[8]))) &
      (fsm_output[6]);
  assign nor_102_nl = ~((fsm_output[8]) | (~ (fsm_output[6])));
  assign mux_337_nl = MUX_s_1_2_2(and_341_nl, nor_102_nl, fsm_output[2]);
  assign nor_103_nl = ~((fsm_output[2]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[8])
      | (~ (fsm_output[6])));
  assign mux_338_nl = MUX_s_1_2_2(mux_337_nl, nor_103_nl, fsm_output[3]);
  assign and_339_nl = (fsm_output[7]) & mux_338_nl;
  assign mux_339_nl = MUX_s_1_2_2((fsm_output[6]), and_339_nl, fsm_output[5]);
  assign nor_104_nl = ~((fsm_output[3]) | and_271_cse | (fsm_output[8]) | (~ (fsm_output[6])));
  assign mux_335_nl = MUX_s_1_2_2(nor_104_nl, (fsm_output[6]), fsm_output[7]);
  assign and_268_nl = (fsm_output[3]) & (~((~(and_271_cse | (fsm_output[8]))) | (fsm_output[6])));
  assign nor_107_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[6]));
  assign nor_108_nl = ~((~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[8])))
      | (fsm_output[6]));
  assign mux_333_nl = MUX_s_1_2_2(nor_107_nl, nor_108_nl, fsm_output[3]);
  assign mux_334_nl = MUX_s_1_2_2(and_268_nl, mux_333_nl, fsm_output[7]);
  assign mux_336_nl = MUX_s_1_2_2(mux_335_nl, mux_334_nl, fsm_output[5]);
  assign mux_340_nl = MUX_s_1_2_2(mux_339_nl, mux_336_nl, fsm_output[4]);
  assign or_438_nl = (fsm_output[5]) | and_tmp_17;
  assign mux_361_nl = MUX_s_1_2_2(not_tmp_111, or_438_nl, fsm_output[6]);
  assign and_247_nl = (fsm_output[5:2]==4'b1111);
  assign nand_37_nl = ~((fsm_output[5]) & ((fsm_output[4]) | or_tmp_167));
  assign mux_362_nl = MUX_s_1_2_2(and_247_nl, nand_37_nl, fsm_output[6]);
  assign or_466_nl = (fsm_output[5:4]!=2'b00) | and_dcpl_44;
  assign mux_363_nl = MUX_s_1_2_2(not_tmp_141, or_466_nl, fsm_output[6]);
  assign and_246_nl = (fsm_output[5:4]==2'b11) & or_tmp_19;
  assign nand_36_nl = ~((fsm_output[5]) & ((fsm_output[4:0]!=5'b00000)));
  assign mux_364_nl = MUX_s_1_2_2(and_246_nl, nand_36_nl, fsm_output[6]);
  assign COMP_LOOP_mux_18_nl = MUX_v_10_2_2(({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))}),
      STAGE_LOOP_lshift_psp_sva, and_dcpl_232);
  assign COMP_LOOP_COMP_LOOP_nand_1_nl = ~(and_dcpl_232 & (~(mux_372_cse & (fsm_output[5])
      & (fsm_output[6]) & (~((fsm_output[4]) | (fsm_output[9]) | (fsm_output[7])))
      & (fsm_output[3]) & (~ (fsm_output[0])))));
  assign nl_acc_nl = ({COMP_LOOP_mux_18_nl , COMP_LOOP_COMP_LOOP_nand_1_nl}) + conv_u2u_10_11({COMP_LOOP_k_9_1_1_sva_7_0
      , 2'b11});
  assign acc_nl = nl_acc_nl[10:0];
  assign z_out = readslicef_11_10_1(acc_nl);
  assign COMP_LOOP_mux_19_nl = MUX_s_1_2_2((tmp_2_lpi_4_dfm[63]), (p_sva[63]), and_dcpl_250);
  assign COMP_LOOP_COMP_LOOP_or_53_nl = (COMP_LOOP_mux_19_nl & COMP_LOOP_nor_3_itm)
      | and_dcpl_241 | and_dcpl_255;
  assign COMP_LOOP_mux1h_70_nl = MUX1HOT_v_51_3_2((tmp_2_lpi_4_dfm[62:12]), (p_sva[62:12]),
      (~ (operator_64_false_acc_mut[62:12])), {and_dcpl_234 , and_dcpl_250 , and_dcpl_255});
  assign COMP_LOOP_and_65_nl = MUX_v_51_2_2(51'b000000000000000000000000000000000000000000000000000,
      COMP_LOOP_mux1h_70_nl, COMP_LOOP_nor_3_itm);
  assign COMP_LOOP_or_31_nl = MUX_v_51_2_2(COMP_LOOP_and_65_nl, 51'b111111111111111111111111111111111111111111111111111,
      and_dcpl_241);
  assign COMP_LOOP_mux1h_71_nl = MUX1HOT_v_2_5_2((tmp_2_lpi_4_dfm[11:10]), (p_sva[11:10]),
      (~ (operator_64_false_acc_mut[11:10])), (VEC_LOOP_j_1_12_0_sva_11_0[11:10]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:10]), {and_dcpl_234 , and_dcpl_250 , and_dcpl_255
      , and_dcpl_278 , and_dcpl_284});
  assign COMP_LOOP_nor_60_nl = ~(and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_287);
  assign COMP_LOOP_and_66_nl = MUX_v_2_2_2(2'b00, COMP_LOOP_mux1h_71_nl, COMP_LOOP_nor_60_nl);
  assign COMP_LOOP_or_32_nl = MUX_v_2_2_2(COMP_LOOP_and_66_nl, 2'b11, and_dcpl_241);
  assign nl_COMP_LOOP_acc_18_nl = (STAGE_LOOP_lshift_psp_sva[9:1]) + conv_u2u_8_9(COMP_LOOP_k_9_1_1_sva_7_0);
  assign COMP_LOOP_acc_18_nl = nl_COMP_LOOP_acc_18_nl[8:0];
  assign COMP_LOOP_or_33_nl = and_dcpl_261 | and_dcpl_270;
  assign COMP_LOOP_or_34_nl = and_dcpl_267 | and_dcpl_274;
  assign COMP_LOOP_mux1h_72_nl = MUX1HOT_v_10_9_2((tmp_2_lpi_4_dfm[9:0]), ({1'b1
      , (~ COMP_LOOP_k_9_1_1_sva_7_0) , 1'b1}), (p_sva[9:0]), (~ (operator_64_false_acc_mut[9:0])),
      ({COMP_LOOP_acc_18_nl , (STAGE_LOOP_lshift_psp_sva[0])}), z_out, (VEC_LOOP_j_1_12_0_sva_11_0[9:0]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[9:0]), ({7'b0000000 , (z_out_4[3:1])}), {and_dcpl_234
      , and_dcpl_241 , and_dcpl_250 , and_dcpl_255 , COMP_LOOP_or_33_nl , COMP_LOOP_or_34_nl
      , and_dcpl_278 , and_dcpl_284 , and_dcpl_287});
  assign COMP_LOOP_or_35_nl = (~(and_dcpl_241 | and_dcpl_250 | and_dcpl_255 | and_dcpl_261
      | and_dcpl_267 | and_dcpl_270 | and_dcpl_274 | and_dcpl_278 | and_dcpl_284
      | and_dcpl_287)) | and_dcpl_234;
  assign COMP_LOOP_COMP_LOOP_or_54_nl = (~((COMP_LOOP_mux_1_itm_mx1[63]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_55_nl = (~((COMP_LOOP_mux_1_itm_mx1[62]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_56_nl = (~((COMP_LOOP_mux_1_itm_mx1[61]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_57_nl = (~((COMP_LOOP_mux_1_itm_mx1[60]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_58_nl = (~((COMP_LOOP_mux_1_itm_mx1[59]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_59_nl = (~((COMP_LOOP_mux_1_itm_mx1[58]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_60_nl = (~((COMP_LOOP_mux_1_itm_mx1[57]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_61_nl = (~((COMP_LOOP_mux_1_itm_mx1[56]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_62_nl = (~((COMP_LOOP_mux_1_itm_mx1[55]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_63_nl = (~((COMP_LOOP_mux_1_itm_mx1[54]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_64_nl = (~((COMP_LOOP_mux_1_itm_mx1[53]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_65_nl = (~((COMP_LOOP_mux_1_itm_mx1[52]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_66_nl = (~((COMP_LOOP_mux_1_itm_mx1[51]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_67_nl = (~((COMP_LOOP_mux_1_itm_mx1[50]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_68_nl = (~((COMP_LOOP_mux_1_itm_mx1[49]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_69_nl = (~((COMP_LOOP_mux_1_itm_mx1[48]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_70_nl = (~((COMP_LOOP_mux_1_itm_mx1[47]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_71_nl = (~((COMP_LOOP_mux_1_itm_mx1[46]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_72_nl = (~((COMP_LOOP_mux_1_itm_mx1[45]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_73_nl = (~((COMP_LOOP_mux_1_itm_mx1[44]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_74_nl = (~((COMP_LOOP_mux_1_itm_mx1[43]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_75_nl = (~((COMP_LOOP_mux_1_itm_mx1[42]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_76_nl = (~((COMP_LOOP_mux_1_itm_mx1[41]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_77_nl = (~((COMP_LOOP_mux_1_itm_mx1[40]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_78_nl = (~((COMP_LOOP_mux_1_itm_mx1[39]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_79_nl = (~((COMP_LOOP_mux_1_itm_mx1[38]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_80_nl = (~((COMP_LOOP_mux_1_itm_mx1[37]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_81_nl = (~((COMP_LOOP_mux_1_itm_mx1[36]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_82_nl = (~((COMP_LOOP_mux_1_itm_mx1[35]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_83_nl = (~((COMP_LOOP_mux_1_itm_mx1[34]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_84_nl = (~((COMP_LOOP_mux_1_itm_mx1[33]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_85_nl = (~((COMP_LOOP_mux_1_itm_mx1[32]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_86_nl = (~((COMP_LOOP_mux_1_itm_mx1[31]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_87_nl = (~((COMP_LOOP_mux_1_itm_mx1[30]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_88_nl = (~((COMP_LOOP_mux_1_itm_mx1[29]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_89_nl = (~((COMP_LOOP_mux_1_itm_mx1[28]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_90_nl = (~((COMP_LOOP_mux_1_itm_mx1[27]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_91_nl = (~((COMP_LOOP_mux_1_itm_mx1[26]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_92_nl = (~((COMP_LOOP_mux_1_itm_mx1[25]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_93_nl = (~((COMP_LOOP_mux_1_itm_mx1[24]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_94_nl = (~((COMP_LOOP_mux_1_itm_mx1[23]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_95_nl = (~((COMP_LOOP_mux_1_itm_mx1[22]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_96_nl = (~((COMP_LOOP_mux_1_itm_mx1[21]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_97_nl = (~((COMP_LOOP_mux_1_itm_mx1[20]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_98_nl = (~((COMP_LOOP_mux_1_itm_mx1[19]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_99_nl = (~((COMP_LOOP_mux_1_itm_mx1[18]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_100_nl = (~((COMP_LOOP_mux_1_itm_mx1[17]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_101_nl = (~((COMP_LOOP_mux_1_itm_mx1[16]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_102_nl = (~((COMP_LOOP_mux_1_itm_mx1[15]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_103_nl = (~((COMP_LOOP_mux_1_itm_mx1[14]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_104_nl = (~((COMP_LOOP_mux_1_itm_mx1[13]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_COMP_LOOP_or_105_nl = (~((COMP_LOOP_mux_1_itm_mx1[12]) | and_dcpl_241
      | and_dcpl_255 | and_dcpl_261 | and_dcpl_267 | and_dcpl_270 | and_dcpl_274
      | and_dcpl_278 | and_dcpl_284 | and_dcpl_287)) | and_dcpl_250;
  assign COMP_LOOP_mux1h_73_nl = MUX1HOT_v_2_3_2((~ (COMP_LOOP_mux_1_itm_mx1[11:10])),
      (VEC_LOOP_j_1_12_0_sva_11_0[11:10]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:10]),
      {and_dcpl_234 , COMP_LOOP_or_23_itm , COMP_LOOP_or_24_itm});
  assign COMP_LOOP_nor_62_nl = ~(and_dcpl_241 | and_dcpl_255 | and_dcpl_278 | and_dcpl_284
      | and_dcpl_287);
  assign COMP_LOOP_and_67_nl = MUX_v_2_2_2(2'b00, COMP_LOOP_mux1h_73_nl, COMP_LOOP_nor_62_nl);
  assign COMP_LOOP_or_36_nl = MUX_v_2_2_2(COMP_LOOP_and_67_nl, 2'b11, and_dcpl_250);
  assign COMP_LOOP_or_38_nl = and_dcpl_241 | and_dcpl_255;
  assign COMP_LOOP_or_39_nl = and_dcpl_278 | and_dcpl_284;
  assign COMP_LOOP_mux1h_74_nl = MUX1HOT_v_10_6_2((~ (COMP_LOOP_mux_1_itm_mx1[9:0])),
      10'b0000000001, (VEC_LOOP_j_1_12_0_sva_11_0[9:0]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[9:0]),
      STAGE_LOOP_lshift_psp_sva, 10'b0000000011, {and_dcpl_234 , COMP_LOOP_or_38_nl
      , COMP_LOOP_or_23_itm , COMP_LOOP_or_24_itm , COMP_LOOP_or_39_nl , and_dcpl_287});
  assign COMP_LOOP_or_37_nl = MUX_v_10_2_2(COMP_LOOP_mux1h_74_nl, 10'b1111111111,
      and_dcpl_250);
  assign nl_acc_1_nl = conv_u2u_65_66({COMP_LOOP_COMP_LOOP_or_53_nl , COMP_LOOP_or_31_nl
      , COMP_LOOP_or_32_nl , COMP_LOOP_mux1h_72_nl , COMP_LOOP_or_35_nl}) + conv_s2u_65_66({COMP_LOOP_COMP_LOOP_or_54_nl
      , COMP_LOOP_COMP_LOOP_or_55_nl , COMP_LOOP_COMP_LOOP_or_56_nl , COMP_LOOP_COMP_LOOP_or_57_nl
      , COMP_LOOP_COMP_LOOP_or_58_nl , COMP_LOOP_COMP_LOOP_or_59_nl , COMP_LOOP_COMP_LOOP_or_60_nl
      , COMP_LOOP_COMP_LOOP_or_61_nl , COMP_LOOP_COMP_LOOP_or_62_nl , COMP_LOOP_COMP_LOOP_or_63_nl
      , COMP_LOOP_COMP_LOOP_or_64_nl , COMP_LOOP_COMP_LOOP_or_65_nl , COMP_LOOP_COMP_LOOP_or_66_nl
      , COMP_LOOP_COMP_LOOP_or_67_nl , COMP_LOOP_COMP_LOOP_or_68_nl , COMP_LOOP_COMP_LOOP_or_69_nl
      , COMP_LOOP_COMP_LOOP_or_70_nl , COMP_LOOP_COMP_LOOP_or_71_nl , COMP_LOOP_COMP_LOOP_or_72_nl
      , COMP_LOOP_COMP_LOOP_or_73_nl , COMP_LOOP_COMP_LOOP_or_74_nl , COMP_LOOP_COMP_LOOP_or_75_nl
      , COMP_LOOP_COMP_LOOP_or_76_nl , COMP_LOOP_COMP_LOOP_or_77_nl , COMP_LOOP_COMP_LOOP_or_78_nl
      , COMP_LOOP_COMP_LOOP_or_79_nl , COMP_LOOP_COMP_LOOP_or_80_nl , COMP_LOOP_COMP_LOOP_or_81_nl
      , COMP_LOOP_COMP_LOOP_or_82_nl , COMP_LOOP_COMP_LOOP_or_83_nl , COMP_LOOP_COMP_LOOP_or_84_nl
      , COMP_LOOP_COMP_LOOP_or_85_nl , COMP_LOOP_COMP_LOOP_or_86_nl , COMP_LOOP_COMP_LOOP_or_87_nl
      , COMP_LOOP_COMP_LOOP_or_88_nl , COMP_LOOP_COMP_LOOP_or_89_nl , COMP_LOOP_COMP_LOOP_or_90_nl
      , COMP_LOOP_COMP_LOOP_or_91_nl , COMP_LOOP_COMP_LOOP_or_92_nl , COMP_LOOP_COMP_LOOP_or_93_nl
      , COMP_LOOP_COMP_LOOP_or_94_nl , COMP_LOOP_COMP_LOOP_or_95_nl , COMP_LOOP_COMP_LOOP_or_96_nl
      , COMP_LOOP_COMP_LOOP_or_97_nl , COMP_LOOP_COMP_LOOP_or_98_nl , COMP_LOOP_COMP_LOOP_or_99_nl
      , COMP_LOOP_COMP_LOOP_or_100_nl , COMP_LOOP_COMP_LOOP_or_101_nl , COMP_LOOP_COMP_LOOP_or_102_nl
      , COMP_LOOP_COMP_LOOP_or_103_nl , COMP_LOOP_COMP_LOOP_or_104_nl , COMP_LOOP_COMP_LOOP_or_105_nl
      , COMP_LOOP_or_36_nl , COMP_LOOP_or_37_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[65:0];
  assign z_out_1 = readslicef_66_65_1(acc_1_nl);
  assign and_468_cse = (fsm_output[6:4]==3'b011) & and_dcpl_20 & (fsm_output[2])
      & (~ (fsm_output[3])) & (fsm_output[8]) & (fsm_output[1]) & (~ (fsm_output[0]));
  assign COMP_LOOP_mux_20_nl = MUX_v_11_2_2((VEC_LOOP_j_1_12_0_sva_11_0[11:1]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:1]),
      and_468_cse);
  assign nl_z_out_2 = COMP_LOOP_mux_20_nl + conv_u2u_8_11(COMP_LOOP_k_9_1_1_sva_7_0);
  assign z_out_2 = nl_z_out_2[10:0];
  assign STAGE_LOOP_mux_2_nl = MUX_v_8_2_2(({4'b0000 , STAGE_LOOP_i_3_0_sva}), COMP_LOOP_k_9_1_1_sva_7_0,
      and_dcpl_232);
  assign nl_z_out_4 = conv_u2u_8_9(STAGE_LOOP_mux_2_nl) + 9'b000000001;
  assign z_out_4 = nl_z_out_4[8:0];
  assign operator_64_false_1_mux_10_nl = MUX_s_1_2_2((~ modExp_exp_1_7_1_sva), (~
      modExp_exp_1_1_1_sva), and_dcpl_343);
  assign operator_64_false_1_mux_11_nl = MUX_s_1_2_2((~ modExp_exp_1_6_1_sva), (~
      modExp_exp_1_7_1_sva), and_dcpl_343);
  assign operator_64_false_1_mux_12_nl = MUX_s_1_2_2((~ modExp_exp_1_5_1_sva), (~
      modExp_exp_1_6_1_sva), and_dcpl_343);
  assign operator_64_false_1_mux_13_nl = MUX_s_1_2_2((~ modExp_exp_1_4_1_sva), (~
      modExp_exp_1_5_1_sva), and_dcpl_343);
  assign operator_64_false_1_mux_14_nl = MUX_s_1_2_2((~ modExp_exp_1_3_1_sva), (~
      modExp_exp_1_4_1_sva), and_dcpl_343);
  assign operator_64_false_1_mux_15_nl = MUX_s_1_2_2((~ modExp_exp_1_2_1_sva), (~
      modExp_exp_1_3_1_sva), and_dcpl_343);
  assign operator_64_false_1_mux_16_nl = MUX_s_1_2_2((~ modExp_exp_1_1_1_sva), (~
      modExp_exp_1_2_1_sva), and_dcpl_343);
  assign nl_operator_64_false_1_acc_nl = ({1'b1 , operator_64_false_1_mux_10_nl ,
      operator_64_false_1_mux_11_nl , operator_64_false_1_mux_12_nl , operator_64_false_1_mux_13_nl
      , operator_64_false_1_mux_14_nl , operator_64_false_1_mux_15_nl , operator_64_false_1_mux_16_nl
      , (~ modExp_exp_1_0_1_sva_1)}) + 9'b000000001;
  assign operator_64_false_1_acc_nl = nl_operator_64_false_1_acc_nl[8:0];
  assign z_out_5_8 = readslicef_9_1_8(operator_64_false_1_acc_nl);

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_6_2;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [5:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    MUX1HOT_v_10_6_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_9_2;
    input [9:0] input_8;
    input [9:0] input_7;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [8:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    result = result | ( input_6 & {10{sel[6]}});
    result = result | ( input_7 & {10{sel[7]}});
    result = result | ( input_8 & {10{sel[8]}});
    MUX1HOT_v_10_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_5_2;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [4:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    result = result | ( input_3 & {11{sel[3]}});
    result = result | ( input_4 & {11{sel[4]}});
    MUX1HOT_v_11_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_5_2;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [4:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    result = result | ( input_4 & {2{sel[4]}});
    MUX1HOT_v_2_5_2 = result;
  end
  endfunction


  function automatic [50:0] MUX1HOT_v_51_3_2;
    input [50:0] input_2;
    input [50:0] input_1;
    input [50:0] input_0;
    input [2:0] sel;
    reg [50:0] result;
  begin
    result = input_0 & {51{sel[0]}};
    result = result | ( input_1 & {51{sel[1]}});
    result = result | ( input_2 & {51{sel[2]}});
    MUX1HOT_v_51_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_20_2;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [19:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    MUX1HOT_v_64_20_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_5_2;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [4:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    MUX1HOT_v_64_5_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_7_2;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [6:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    MUX1HOT_v_64_7_2 = result;
  end
  endfunction


  function automatic [64:0] MUX1HOT_v_65_3_2;
    input [64:0] input_2;
    input [64:0] input_1;
    input [64:0] input_0;
    input [2:0] sel;
    reg [64:0] result;
  begin
    result = input_0 & {65{sel[0]}};
    result = result | ( input_1 & {65{sel[1]}});
    result = result | ( input_2 & {65{sel[2]}});
    MUX1HOT_v_65_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [50:0] MUX_v_51_2_2;
    input [50:0] input_0;
    input [50:0] input_1;
    input [0:0] sel;
    reg [50:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_51_2_2 = result;
  end
  endfunction


  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [0:0] readslicef_65_1_64;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 64;
    readslicef_65_1_64 = tmp[0:0];
  end
  endfunction


  function automatic [64:0] readslicef_66_65_1;
    input [65:0] vector;
    reg [65:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_66_65_1 = tmp[64:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [65:0] conv_s2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_s2u_65_66 = {vector[64], vector};
  end
  endfunction


  function automatic [64:0] conv_u2s_64_65 ;
    input [63:0]  vector ;
  begin
    conv_u2s_64_65 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_11 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [65:0] conv_u2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_u2u_65_66 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [10:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [10:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [64:0] operator_66_true_div_cmp_a;
  wire [10:0] operator_66_true_div_cmp_b;
  wire [64:0] operator_66_true_div_cmp_z;
  wire [10:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(operator_66_true_div_cmp_b),
      .z(operator_66_true_div_cmp_z)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_11_64_2048_2048_64_1_gen
      vec_rsc_0_0_i (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_11_64_2048_2048_64_1_gen
      vec_rsc_0_1_i (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .operator_66_true_div_cmp_a(operator_66_true_div_cmp_a),
      .operator_66_true_div_cmp_b(operator_66_true_div_cmp_b),
      .operator_66_true_div_cmp_z(operator_66_true_div_cmp_z),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff)
    );
endmodule



