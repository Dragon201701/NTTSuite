
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Wed Jun 30 21:47:46 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [8:0] adra;
  input [8:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_8_tr0, modExp_while_C_40_tr0, COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_1_while_C_40_tr0, COMP_LOOP_C_65_tr0, COMP_LOOP_2_modExp_1_while_C_40_tr0,
      COMP_LOOP_C_130_tr0, COMP_LOOP_3_modExp_1_while_C_40_tr0, COMP_LOOP_C_195_tr0,
      COMP_LOOP_4_modExp_1_while_C_40_tr0, COMP_LOOP_C_260_tr0, COMP_LOOP_5_modExp_1_while_C_40_tr0,
      COMP_LOOP_C_325_tr0, COMP_LOOP_6_modExp_1_while_C_40_tr0, COMP_LOOP_C_390_tr0,
      COMP_LOOP_7_modExp_1_while_C_40_tr0, COMP_LOOP_C_455_tr0, COMP_LOOP_8_modExp_1_while_C_40_tr0,
      COMP_LOOP_C_520_tr0, VEC_LOOP_C_0_tr0, STAGE_LOOP_C_9_tr0
);
  input clk;
  input rst;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;
  input STAGE_LOOP_C_8_tr0;
  input modExp_while_C_40_tr0;
  input COMP_LOOP_C_1_tr0;
  input COMP_LOOP_1_modExp_1_while_C_40_tr0;
  input COMP_LOOP_C_65_tr0;
  input COMP_LOOP_2_modExp_1_while_C_40_tr0;
  input COMP_LOOP_C_130_tr0;
  input COMP_LOOP_3_modExp_1_while_C_40_tr0;
  input COMP_LOOP_C_195_tr0;
  input COMP_LOOP_4_modExp_1_while_C_40_tr0;
  input COMP_LOOP_C_260_tr0;
  input COMP_LOOP_5_modExp_1_while_C_40_tr0;
  input COMP_LOOP_C_325_tr0;
  input COMP_LOOP_6_modExp_1_while_C_40_tr0;
  input COMP_LOOP_C_390_tr0;
  input COMP_LOOP_7_modExp_1_while_C_40_tr0;
  input COMP_LOOP_C_455_tr0;
  input COMP_LOOP_8_modExp_1_while_C_40_tr0;
  input COMP_LOOP_C_520_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_9_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 10'd0,
    STAGE_LOOP_C_0 = 10'd1,
    STAGE_LOOP_C_1 = 10'd2,
    STAGE_LOOP_C_2 = 10'd3,
    STAGE_LOOP_C_3 = 10'd4,
    STAGE_LOOP_C_4 = 10'd5,
    STAGE_LOOP_C_5 = 10'd6,
    STAGE_LOOP_C_6 = 10'd7,
    STAGE_LOOP_C_7 = 10'd8,
    STAGE_LOOP_C_8 = 10'd9,
    modExp_while_C_0 = 10'd10,
    modExp_while_C_1 = 10'd11,
    modExp_while_C_2 = 10'd12,
    modExp_while_C_3 = 10'd13,
    modExp_while_C_4 = 10'd14,
    modExp_while_C_5 = 10'd15,
    modExp_while_C_6 = 10'd16,
    modExp_while_C_7 = 10'd17,
    modExp_while_C_8 = 10'd18,
    modExp_while_C_9 = 10'd19,
    modExp_while_C_10 = 10'd20,
    modExp_while_C_11 = 10'd21,
    modExp_while_C_12 = 10'd22,
    modExp_while_C_13 = 10'd23,
    modExp_while_C_14 = 10'd24,
    modExp_while_C_15 = 10'd25,
    modExp_while_C_16 = 10'd26,
    modExp_while_C_17 = 10'd27,
    modExp_while_C_18 = 10'd28,
    modExp_while_C_19 = 10'd29,
    modExp_while_C_20 = 10'd30,
    modExp_while_C_21 = 10'd31,
    modExp_while_C_22 = 10'd32,
    modExp_while_C_23 = 10'd33,
    modExp_while_C_24 = 10'd34,
    modExp_while_C_25 = 10'd35,
    modExp_while_C_26 = 10'd36,
    modExp_while_C_27 = 10'd37,
    modExp_while_C_28 = 10'd38,
    modExp_while_C_29 = 10'd39,
    modExp_while_C_30 = 10'd40,
    modExp_while_C_31 = 10'd41,
    modExp_while_C_32 = 10'd42,
    modExp_while_C_33 = 10'd43,
    modExp_while_C_34 = 10'd44,
    modExp_while_C_35 = 10'd45,
    modExp_while_C_36 = 10'd46,
    modExp_while_C_37 = 10'd47,
    modExp_while_C_38 = 10'd48,
    modExp_while_C_39 = 10'd49,
    modExp_while_C_40 = 10'd50,
    COMP_LOOP_C_0 = 10'd51,
    COMP_LOOP_C_1 = 10'd52,
    COMP_LOOP_1_modExp_1_while_C_0 = 10'd53,
    COMP_LOOP_1_modExp_1_while_C_1 = 10'd54,
    COMP_LOOP_1_modExp_1_while_C_2 = 10'd55,
    COMP_LOOP_1_modExp_1_while_C_3 = 10'd56,
    COMP_LOOP_1_modExp_1_while_C_4 = 10'd57,
    COMP_LOOP_1_modExp_1_while_C_5 = 10'd58,
    COMP_LOOP_1_modExp_1_while_C_6 = 10'd59,
    COMP_LOOP_1_modExp_1_while_C_7 = 10'd60,
    COMP_LOOP_1_modExp_1_while_C_8 = 10'd61,
    COMP_LOOP_1_modExp_1_while_C_9 = 10'd62,
    COMP_LOOP_1_modExp_1_while_C_10 = 10'd63,
    COMP_LOOP_1_modExp_1_while_C_11 = 10'd64,
    COMP_LOOP_1_modExp_1_while_C_12 = 10'd65,
    COMP_LOOP_1_modExp_1_while_C_13 = 10'd66,
    COMP_LOOP_1_modExp_1_while_C_14 = 10'd67,
    COMP_LOOP_1_modExp_1_while_C_15 = 10'd68,
    COMP_LOOP_1_modExp_1_while_C_16 = 10'd69,
    COMP_LOOP_1_modExp_1_while_C_17 = 10'd70,
    COMP_LOOP_1_modExp_1_while_C_18 = 10'd71,
    COMP_LOOP_1_modExp_1_while_C_19 = 10'd72,
    COMP_LOOP_1_modExp_1_while_C_20 = 10'd73,
    COMP_LOOP_1_modExp_1_while_C_21 = 10'd74,
    COMP_LOOP_1_modExp_1_while_C_22 = 10'd75,
    COMP_LOOP_1_modExp_1_while_C_23 = 10'd76,
    COMP_LOOP_1_modExp_1_while_C_24 = 10'd77,
    COMP_LOOP_1_modExp_1_while_C_25 = 10'd78,
    COMP_LOOP_1_modExp_1_while_C_26 = 10'd79,
    COMP_LOOP_1_modExp_1_while_C_27 = 10'd80,
    COMP_LOOP_1_modExp_1_while_C_28 = 10'd81,
    COMP_LOOP_1_modExp_1_while_C_29 = 10'd82,
    COMP_LOOP_1_modExp_1_while_C_30 = 10'd83,
    COMP_LOOP_1_modExp_1_while_C_31 = 10'd84,
    COMP_LOOP_1_modExp_1_while_C_32 = 10'd85,
    COMP_LOOP_1_modExp_1_while_C_33 = 10'd86,
    COMP_LOOP_1_modExp_1_while_C_34 = 10'd87,
    COMP_LOOP_1_modExp_1_while_C_35 = 10'd88,
    COMP_LOOP_1_modExp_1_while_C_36 = 10'd89,
    COMP_LOOP_1_modExp_1_while_C_37 = 10'd90,
    COMP_LOOP_1_modExp_1_while_C_38 = 10'd91,
    COMP_LOOP_1_modExp_1_while_C_39 = 10'd92,
    COMP_LOOP_1_modExp_1_while_C_40 = 10'd93,
    COMP_LOOP_C_2 = 10'd94,
    COMP_LOOP_C_3 = 10'd95,
    COMP_LOOP_C_4 = 10'd96,
    COMP_LOOP_C_5 = 10'd97,
    COMP_LOOP_C_6 = 10'd98,
    COMP_LOOP_C_7 = 10'd99,
    COMP_LOOP_C_8 = 10'd100,
    COMP_LOOP_C_9 = 10'd101,
    COMP_LOOP_C_10 = 10'd102,
    COMP_LOOP_C_11 = 10'd103,
    COMP_LOOP_C_12 = 10'd104,
    COMP_LOOP_C_13 = 10'd105,
    COMP_LOOP_C_14 = 10'd106,
    COMP_LOOP_C_15 = 10'd107,
    COMP_LOOP_C_16 = 10'd108,
    COMP_LOOP_C_17 = 10'd109,
    COMP_LOOP_C_18 = 10'd110,
    COMP_LOOP_C_19 = 10'd111,
    COMP_LOOP_C_20 = 10'd112,
    COMP_LOOP_C_21 = 10'd113,
    COMP_LOOP_C_22 = 10'd114,
    COMP_LOOP_C_23 = 10'd115,
    COMP_LOOP_C_24 = 10'd116,
    COMP_LOOP_C_25 = 10'd117,
    COMP_LOOP_C_26 = 10'd118,
    COMP_LOOP_C_27 = 10'd119,
    COMP_LOOP_C_28 = 10'd120,
    COMP_LOOP_C_29 = 10'd121,
    COMP_LOOP_C_30 = 10'd122,
    COMP_LOOP_C_31 = 10'd123,
    COMP_LOOP_C_32 = 10'd124,
    COMP_LOOP_C_33 = 10'd125,
    COMP_LOOP_C_34 = 10'd126,
    COMP_LOOP_C_35 = 10'd127,
    COMP_LOOP_C_36 = 10'd128,
    COMP_LOOP_C_37 = 10'd129,
    COMP_LOOP_C_38 = 10'd130,
    COMP_LOOP_C_39 = 10'd131,
    COMP_LOOP_C_40 = 10'd132,
    COMP_LOOP_C_41 = 10'd133,
    COMP_LOOP_C_42 = 10'd134,
    COMP_LOOP_C_43 = 10'd135,
    COMP_LOOP_C_44 = 10'd136,
    COMP_LOOP_C_45 = 10'd137,
    COMP_LOOP_C_46 = 10'd138,
    COMP_LOOP_C_47 = 10'd139,
    COMP_LOOP_C_48 = 10'd140,
    COMP_LOOP_C_49 = 10'd141,
    COMP_LOOP_C_50 = 10'd142,
    COMP_LOOP_C_51 = 10'd143,
    COMP_LOOP_C_52 = 10'd144,
    COMP_LOOP_C_53 = 10'd145,
    COMP_LOOP_C_54 = 10'd146,
    COMP_LOOP_C_55 = 10'd147,
    COMP_LOOP_C_56 = 10'd148,
    COMP_LOOP_C_57 = 10'd149,
    COMP_LOOP_C_58 = 10'd150,
    COMP_LOOP_C_59 = 10'd151,
    COMP_LOOP_C_60 = 10'd152,
    COMP_LOOP_C_61 = 10'd153,
    COMP_LOOP_C_62 = 10'd154,
    COMP_LOOP_C_63 = 10'd155,
    COMP_LOOP_C_64 = 10'd156,
    COMP_LOOP_C_65 = 10'd157,
    COMP_LOOP_C_66 = 10'd158,
    COMP_LOOP_2_modExp_1_while_C_0 = 10'd159,
    COMP_LOOP_2_modExp_1_while_C_1 = 10'd160,
    COMP_LOOP_2_modExp_1_while_C_2 = 10'd161,
    COMP_LOOP_2_modExp_1_while_C_3 = 10'd162,
    COMP_LOOP_2_modExp_1_while_C_4 = 10'd163,
    COMP_LOOP_2_modExp_1_while_C_5 = 10'd164,
    COMP_LOOP_2_modExp_1_while_C_6 = 10'd165,
    COMP_LOOP_2_modExp_1_while_C_7 = 10'd166,
    COMP_LOOP_2_modExp_1_while_C_8 = 10'd167,
    COMP_LOOP_2_modExp_1_while_C_9 = 10'd168,
    COMP_LOOP_2_modExp_1_while_C_10 = 10'd169,
    COMP_LOOP_2_modExp_1_while_C_11 = 10'd170,
    COMP_LOOP_2_modExp_1_while_C_12 = 10'd171,
    COMP_LOOP_2_modExp_1_while_C_13 = 10'd172,
    COMP_LOOP_2_modExp_1_while_C_14 = 10'd173,
    COMP_LOOP_2_modExp_1_while_C_15 = 10'd174,
    COMP_LOOP_2_modExp_1_while_C_16 = 10'd175,
    COMP_LOOP_2_modExp_1_while_C_17 = 10'd176,
    COMP_LOOP_2_modExp_1_while_C_18 = 10'd177,
    COMP_LOOP_2_modExp_1_while_C_19 = 10'd178,
    COMP_LOOP_2_modExp_1_while_C_20 = 10'd179,
    COMP_LOOP_2_modExp_1_while_C_21 = 10'd180,
    COMP_LOOP_2_modExp_1_while_C_22 = 10'd181,
    COMP_LOOP_2_modExp_1_while_C_23 = 10'd182,
    COMP_LOOP_2_modExp_1_while_C_24 = 10'd183,
    COMP_LOOP_2_modExp_1_while_C_25 = 10'd184,
    COMP_LOOP_2_modExp_1_while_C_26 = 10'd185,
    COMP_LOOP_2_modExp_1_while_C_27 = 10'd186,
    COMP_LOOP_2_modExp_1_while_C_28 = 10'd187,
    COMP_LOOP_2_modExp_1_while_C_29 = 10'd188,
    COMP_LOOP_2_modExp_1_while_C_30 = 10'd189,
    COMP_LOOP_2_modExp_1_while_C_31 = 10'd190,
    COMP_LOOP_2_modExp_1_while_C_32 = 10'd191,
    COMP_LOOP_2_modExp_1_while_C_33 = 10'd192,
    COMP_LOOP_2_modExp_1_while_C_34 = 10'd193,
    COMP_LOOP_2_modExp_1_while_C_35 = 10'd194,
    COMP_LOOP_2_modExp_1_while_C_36 = 10'd195,
    COMP_LOOP_2_modExp_1_while_C_37 = 10'd196,
    COMP_LOOP_2_modExp_1_while_C_38 = 10'd197,
    COMP_LOOP_2_modExp_1_while_C_39 = 10'd198,
    COMP_LOOP_2_modExp_1_while_C_40 = 10'd199,
    COMP_LOOP_C_67 = 10'd200,
    COMP_LOOP_C_68 = 10'd201,
    COMP_LOOP_C_69 = 10'd202,
    COMP_LOOP_C_70 = 10'd203,
    COMP_LOOP_C_71 = 10'd204,
    COMP_LOOP_C_72 = 10'd205,
    COMP_LOOP_C_73 = 10'd206,
    COMP_LOOP_C_74 = 10'd207,
    COMP_LOOP_C_75 = 10'd208,
    COMP_LOOP_C_76 = 10'd209,
    COMP_LOOP_C_77 = 10'd210,
    COMP_LOOP_C_78 = 10'd211,
    COMP_LOOP_C_79 = 10'd212,
    COMP_LOOP_C_80 = 10'd213,
    COMP_LOOP_C_81 = 10'd214,
    COMP_LOOP_C_82 = 10'd215,
    COMP_LOOP_C_83 = 10'd216,
    COMP_LOOP_C_84 = 10'd217,
    COMP_LOOP_C_85 = 10'd218,
    COMP_LOOP_C_86 = 10'd219,
    COMP_LOOP_C_87 = 10'd220,
    COMP_LOOP_C_88 = 10'd221,
    COMP_LOOP_C_89 = 10'd222,
    COMP_LOOP_C_90 = 10'd223,
    COMP_LOOP_C_91 = 10'd224,
    COMP_LOOP_C_92 = 10'd225,
    COMP_LOOP_C_93 = 10'd226,
    COMP_LOOP_C_94 = 10'd227,
    COMP_LOOP_C_95 = 10'd228,
    COMP_LOOP_C_96 = 10'd229,
    COMP_LOOP_C_97 = 10'd230,
    COMP_LOOP_C_98 = 10'd231,
    COMP_LOOP_C_99 = 10'd232,
    COMP_LOOP_C_100 = 10'd233,
    COMP_LOOP_C_101 = 10'd234,
    COMP_LOOP_C_102 = 10'd235,
    COMP_LOOP_C_103 = 10'd236,
    COMP_LOOP_C_104 = 10'd237,
    COMP_LOOP_C_105 = 10'd238,
    COMP_LOOP_C_106 = 10'd239,
    COMP_LOOP_C_107 = 10'd240,
    COMP_LOOP_C_108 = 10'd241,
    COMP_LOOP_C_109 = 10'd242,
    COMP_LOOP_C_110 = 10'd243,
    COMP_LOOP_C_111 = 10'd244,
    COMP_LOOP_C_112 = 10'd245,
    COMP_LOOP_C_113 = 10'd246,
    COMP_LOOP_C_114 = 10'd247,
    COMP_LOOP_C_115 = 10'd248,
    COMP_LOOP_C_116 = 10'd249,
    COMP_LOOP_C_117 = 10'd250,
    COMP_LOOP_C_118 = 10'd251,
    COMP_LOOP_C_119 = 10'd252,
    COMP_LOOP_C_120 = 10'd253,
    COMP_LOOP_C_121 = 10'd254,
    COMP_LOOP_C_122 = 10'd255,
    COMP_LOOP_C_123 = 10'd256,
    COMP_LOOP_C_124 = 10'd257,
    COMP_LOOP_C_125 = 10'd258,
    COMP_LOOP_C_126 = 10'd259,
    COMP_LOOP_C_127 = 10'd260,
    COMP_LOOP_C_128 = 10'd261,
    COMP_LOOP_C_129 = 10'd262,
    COMP_LOOP_C_130 = 10'd263,
    COMP_LOOP_C_131 = 10'd264,
    COMP_LOOP_3_modExp_1_while_C_0 = 10'd265,
    COMP_LOOP_3_modExp_1_while_C_1 = 10'd266,
    COMP_LOOP_3_modExp_1_while_C_2 = 10'd267,
    COMP_LOOP_3_modExp_1_while_C_3 = 10'd268,
    COMP_LOOP_3_modExp_1_while_C_4 = 10'd269,
    COMP_LOOP_3_modExp_1_while_C_5 = 10'd270,
    COMP_LOOP_3_modExp_1_while_C_6 = 10'd271,
    COMP_LOOP_3_modExp_1_while_C_7 = 10'd272,
    COMP_LOOP_3_modExp_1_while_C_8 = 10'd273,
    COMP_LOOP_3_modExp_1_while_C_9 = 10'd274,
    COMP_LOOP_3_modExp_1_while_C_10 = 10'd275,
    COMP_LOOP_3_modExp_1_while_C_11 = 10'd276,
    COMP_LOOP_3_modExp_1_while_C_12 = 10'd277,
    COMP_LOOP_3_modExp_1_while_C_13 = 10'd278,
    COMP_LOOP_3_modExp_1_while_C_14 = 10'd279,
    COMP_LOOP_3_modExp_1_while_C_15 = 10'd280,
    COMP_LOOP_3_modExp_1_while_C_16 = 10'd281,
    COMP_LOOP_3_modExp_1_while_C_17 = 10'd282,
    COMP_LOOP_3_modExp_1_while_C_18 = 10'd283,
    COMP_LOOP_3_modExp_1_while_C_19 = 10'd284,
    COMP_LOOP_3_modExp_1_while_C_20 = 10'd285,
    COMP_LOOP_3_modExp_1_while_C_21 = 10'd286,
    COMP_LOOP_3_modExp_1_while_C_22 = 10'd287,
    COMP_LOOP_3_modExp_1_while_C_23 = 10'd288,
    COMP_LOOP_3_modExp_1_while_C_24 = 10'd289,
    COMP_LOOP_3_modExp_1_while_C_25 = 10'd290,
    COMP_LOOP_3_modExp_1_while_C_26 = 10'd291,
    COMP_LOOP_3_modExp_1_while_C_27 = 10'd292,
    COMP_LOOP_3_modExp_1_while_C_28 = 10'd293,
    COMP_LOOP_3_modExp_1_while_C_29 = 10'd294,
    COMP_LOOP_3_modExp_1_while_C_30 = 10'd295,
    COMP_LOOP_3_modExp_1_while_C_31 = 10'd296,
    COMP_LOOP_3_modExp_1_while_C_32 = 10'd297,
    COMP_LOOP_3_modExp_1_while_C_33 = 10'd298,
    COMP_LOOP_3_modExp_1_while_C_34 = 10'd299,
    COMP_LOOP_3_modExp_1_while_C_35 = 10'd300,
    COMP_LOOP_3_modExp_1_while_C_36 = 10'd301,
    COMP_LOOP_3_modExp_1_while_C_37 = 10'd302,
    COMP_LOOP_3_modExp_1_while_C_38 = 10'd303,
    COMP_LOOP_3_modExp_1_while_C_39 = 10'd304,
    COMP_LOOP_3_modExp_1_while_C_40 = 10'd305,
    COMP_LOOP_C_132 = 10'd306,
    COMP_LOOP_C_133 = 10'd307,
    COMP_LOOP_C_134 = 10'd308,
    COMP_LOOP_C_135 = 10'd309,
    COMP_LOOP_C_136 = 10'd310,
    COMP_LOOP_C_137 = 10'd311,
    COMP_LOOP_C_138 = 10'd312,
    COMP_LOOP_C_139 = 10'd313,
    COMP_LOOP_C_140 = 10'd314,
    COMP_LOOP_C_141 = 10'd315,
    COMP_LOOP_C_142 = 10'd316,
    COMP_LOOP_C_143 = 10'd317,
    COMP_LOOP_C_144 = 10'd318,
    COMP_LOOP_C_145 = 10'd319,
    COMP_LOOP_C_146 = 10'd320,
    COMP_LOOP_C_147 = 10'd321,
    COMP_LOOP_C_148 = 10'd322,
    COMP_LOOP_C_149 = 10'd323,
    COMP_LOOP_C_150 = 10'd324,
    COMP_LOOP_C_151 = 10'd325,
    COMP_LOOP_C_152 = 10'd326,
    COMP_LOOP_C_153 = 10'd327,
    COMP_LOOP_C_154 = 10'd328,
    COMP_LOOP_C_155 = 10'd329,
    COMP_LOOP_C_156 = 10'd330,
    COMP_LOOP_C_157 = 10'd331,
    COMP_LOOP_C_158 = 10'd332,
    COMP_LOOP_C_159 = 10'd333,
    COMP_LOOP_C_160 = 10'd334,
    COMP_LOOP_C_161 = 10'd335,
    COMP_LOOP_C_162 = 10'd336,
    COMP_LOOP_C_163 = 10'd337,
    COMP_LOOP_C_164 = 10'd338,
    COMP_LOOP_C_165 = 10'd339,
    COMP_LOOP_C_166 = 10'd340,
    COMP_LOOP_C_167 = 10'd341,
    COMP_LOOP_C_168 = 10'd342,
    COMP_LOOP_C_169 = 10'd343,
    COMP_LOOP_C_170 = 10'd344,
    COMP_LOOP_C_171 = 10'd345,
    COMP_LOOP_C_172 = 10'd346,
    COMP_LOOP_C_173 = 10'd347,
    COMP_LOOP_C_174 = 10'd348,
    COMP_LOOP_C_175 = 10'd349,
    COMP_LOOP_C_176 = 10'd350,
    COMP_LOOP_C_177 = 10'd351,
    COMP_LOOP_C_178 = 10'd352,
    COMP_LOOP_C_179 = 10'd353,
    COMP_LOOP_C_180 = 10'd354,
    COMP_LOOP_C_181 = 10'd355,
    COMP_LOOP_C_182 = 10'd356,
    COMP_LOOP_C_183 = 10'd357,
    COMP_LOOP_C_184 = 10'd358,
    COMP_LOOP_C_185 = 10'd359,
    COMP_LOOP_C_186 = 10'd360,
    COMP_LOOP_C_187 = 10'd361,
    COMP_LOOP_C_188 = 10'd362,
    COMP_LOOP_C_189 = 10'd363,
    COMP_LOOP_C_190 = 10'd364,
    COMP_LOOP_C_191 = 10'd365,
    COMP_LOOP_C_192 = 10'd366,
    COMP_LOOP_C_193 = 10'd367,
    COMP_LOOP_C_194 = 10'd368,
    COMP_LOOP_C_195 = 10'd369,
    COMP_LOOP_C_196 = 10'd370,
    COMP_LOOP_4_modExp_1_while_C_0 = 10'd371,
    COMP_LOOP_4_modExp_1_while_C_1 = 10'd372,
    COMP_LOOP_4_modExp_1_while_C_2 = 10'd373,
    COMP_LOOP_4_modExp_1_while_C_3 = 10'd374,
    COMP_LOOP_4_modExp_1_while_C_4 = 10'd375,
    COMP_LOOP_4_modExp_1_while_C_5 = 10'd376,
    COMP_LOOP_4_modExp_1_while_C_6 = 10'd377,
    COMP_LOOP_4_modExp_1_while_C_7 = 10'd378,
    COMP_LOOP_4_modExp_1_while_C_8 = 10'd379,
    COMP_LOOP_4_modExp_1_while_C_9 = 10'd380,
    COMP_LOOP_4_modExp_1_while_C_10 = 10'd381,
    COMP_LOOP_4_modExp_1_while_C_11 = 10'd382,
    COMP_LOOP_4_modExp_1_while_C_12 = 10'd383,
    COMP_LOOP_4_modExp_1_while_C_13 = 10'd384,
    COMP_LOOP_4_modExp_1_while_C_14 = 10'd385,
    COMP_LOOP_4_modExp_1_while_C_15 = 10'd386,
    COMP_LOOP_4_modExp_1_while_C_16 = 10'd387,
    COMP_LOOP_4_modExp_1_while_C_17 = 10'd388,
    COMP_LOOP_4_modExp_1_while_C_18 = 10'd389,
    COMP_LOOP_4_modExp_1_while_C_19 = 10'd390,
    COMP_LOOP_4_modExp_1_while_C_20 = 10'd391,
    COMP_LOOP_4_modExp_1_while_C_21 = 10'd392,
    COMP_LOOP_4_modExp_1_while_C_22 = 10'd393,
    COMP_LOOP_4_modExp_1_while_C_23 = 10'd394,
    COMP_LOOP_4_modExp_1_while_C_24 = 10'd395,
    COMP_LOOP_4_modExp_1_while_C_25 = 10'd396,
    COMP_LOOP_4_modExp_1_while_C_26 = 10'd397,
    COMP_LOOP_4_modExp_1_while_C_27 = 10'd398,
    COMP_LOOP_4_modExp_1_while_C_28 = 10'd399,
    COMP_LOOP_4_modExp_1_while_C_29 = 10'd400,
    COMP_LOOP_4_modExp_1_while_C_30 = 10'd401,
    COMP_LOOP_4_modExp_1_while_C_31 = 10'd402,
    COMP_LOOP_4_modExp_1_while_C_32 = 10'd403,
    COMP_LOOP_4_modExp_1_while_C_33 = 10'd404,
    COMP_LOOP_4_modExp_1_while_C_34 = 10'd405,
    COMP_LOOP_4_modExp_1_while_C_35 = 10'd406,
    COMP_LOOP_4_modExp_1_while_C_36 = 10'd407,
    COMP_LOOP_4_modExp_1_while_C_37 = 10'd408,
    COMP_LOOP_4_modExp_1_while_C_38 = 10'd409,
    COMP_LOOP_4_modExp_1_while_C_39 = 10'd410,
    COMP_LOOP_4_modExp_1_while_C_40 = 10'd411,
    COMP_LOOP_C_197 = 10'd412,
    COMP_LOOP_C_198 = 10'd413,
    COMP_LOOP_C_199 = 10'd414,
    COMP_LOOP_C_200 = 10'd415,
    COMP_LOOP_C_201 = 10'd416,
    COMP_LOOP_C_202 = 10'd417,
    COMP_LOOP_C_203 = 10'd418,
    COMP_LOOP_C_204 = 10'd419,
    COMP_LOOP_C_205 = 10'd420,
    COMP_LOOP_C_206 = 10'd421,
    COMP_LOOP_C_207 = 10'd422,
    COMP_LOOP_C_208 = 10'd423,
    COMP_LOOP_C_209 = 10'd424,
    COMP_LOOP_C_210 = 10'd425,
    COMP_LOOP_C_211 = 10'd426,
    COMP_LOOP_C_212 = 10'd427,
    COMP_LOOP_C_213 = 10'd428,
    COMP_LOOP_C_214 = 10'd429,
    COMP_LOOP_C_215 = 10'd430,
    COMP_LOOP_C_216 = 10'd431,
    COMP_LOOP_C_217 = 10'd432,
    COMP_LOOP_C_218 = 10'd433,
    COMP_LOOP_C_219 = 10'd434,
    COMP_LOOP_C_220 = 10'd435,
    COMP_LOOP_C_221 = 10'd436,
    COMP_LOOP_C_222 = 10'd437,
    COMP_LOOP_C_223 = 10'd438,
    COMP_LOOP_C_224 = 10'd439,
    COMP_LOOP_C_225 = 10'd440,
    COMP_LOOP_C_226 = 10'd441,
    COMP_LOOP_C_227 = 10'd442,
    COMP_LOOP_C_228 = 10'd443,
    COMP_LOOP_C_229 = 10'd444,
    COMP_LOOP_C_230 = 10'd445,
    COMP_LOOP_C_231 = 10'd446,
    COMP_LOOP_C_232 = 10'd447,
    COMP_LOOP_C_233 = 10'd448,
    COMP_LOOP_C_234 = 10'd449,
    COMP_LOOP_C_235 = 10'd450,
    COMP_LOOP_C_236 = 10'd451,
    COMP_LOOP_C_237 = 10'd452,
    COMP_LOOP_C_238 = 10'd453,
    COMP_LOOP_C_239 = 10'd454,
    COMP_LOOP_C_240 = 10'd455,
    COMP_LOOP_C_241 = 10'd456,
    COMP_LOOP_C_242 = 10'd457,
    COMP_LOOP_C_243 = 10'd458,
    COMP_LOOP_C_244 = 10'd459,
    COMP_LOOP_C_245 = 10'd460,
    COMP_LOOP_C_246 = 10'd461,
    COMP_LOOP_C_247 = 10'd462,
    COMP_LOOP_C_248 = 10'd463,
    COMP_LOOP_C_249 = 10'd464,
    COMP_LOOP_C_250 = 10'd465,
    COMP_LOOP_C_251 = 10'd466,
    COMP_LOOP_C_252 = 10'd467,
    COMP_LOOP_C_253 = 10'd468,
    COMP_LOOP_C_254 = 10'd469,
    COMP_LOOP_C_255 = 10'd470,
    COMP_LOOP_C_256 = 10'd471,
    COMP_LOOP_C_257 = 10'd472,
    COMP_LOOP_C_258 = 10'd473,
    COMP_LOOP_C_259 = 10'd474,
    COMP_LOOP_C_260 = 10'd475,
    COMP_LOOP_C_261 = 10'd476,
    COMP_LOOP_5_modExp_1_while_C_0 = 10'd477,
    COMP_LOOP_5_modExp_1_while_C_1 = 10'd478,
    COMP_LOOP_5_modExp_1_while_C_2 = 10'd479,
    COMP_LOOP_5_modExp_1_while_C_3 = 10'd480,
    COMP_LOOP_5_modExp_1_while_C_4 = 10'd481,
    COMP_LOOP_5_modExp_1_while_C_5 = 10'd482,
    COMP_LOOP_5_modExp_1_while_C_6 = 10'd483,
    COMP_LOOP_5_modExp_1_while_C_7 = 10'd484,
    COMP_LOOP_5_modExp_1_while_C_8 = 10'd485,
    COMP_LOOP_5_modExp_1_while_C_9 = 10'd486,
    COMP_LOOP_5_modExp_1_while_C_10 = 10'd487,
    COMP_LOOP_5_modExp_1_while_C_11 = 10'd488,
    COMP_LOOP_5_modExp_1_while_C_12 = 10'd489,
    COMP_LOOP_5_modExp_1_while_C_13 = 10'd490,
    COMP_LOOP_5_modExp_1_while_C_14 = 10'd491,
    COMP_LOOP_5_modExp_1_while_C_15 = 10'd492,
    COMP_LOOP_5_modExp_1_while_C_16 = 10'd493,
    COMP_LOOP_5_modExp_1_while_C_17 = 10'd494,
    COMP_LOOP_5_modExp_1_while_C_18 = 10'd495,
    COMP_LOOP_5_modExp_1_while_C_19 = 10'd496,
    COMP_LOOP_5_modExp_1_while_C_20 = 10'd497,
    COMP_LOOP_5_modExp_1_while_C_21 = 10'd498,
    COMP_LOOP_5_modExp_1_while_C_22 = 10'd499,
    COMP_LOOP_5_modExp_1_while_C_23 = 10'd500,
    COMP_LOOP_5_modExp_1_while_C_24 = 10'd501,
    COMP_LOOP_5_modExp_1_while_C_25 = 10'd502,
    COMP_LOOP_5_modExp_1_while_C_26 = 10'd503,
    COMP_LOOP_5_modExp_1_while_C_27 = 10'd504,
    COMP_LOOP_5_modExp_1_while_C_28 = 10'd505,
    COMP_LOOP_5_modExp_1_while_C_29 = 10'd506,
    COMP_LOOP_5_modExp_1_while_C_30 = 10'd507,
    COMP_LOOP_5_modExp_1_while_C_31 = 10'd508,
    COMP_LOOP_5_modExp_1_while_C_32 = 10'd509,
    COMP_LOOP_5_modExp_1_while_C_33 = 10'd510,
    COMP_LOOP_5_modExp_1_while_C_34 = 10'd511,
    COMP_LOOP_5_modExp_1_while_C_35 = 10'd512,
    COMP_LOOP_5_modExp_1_while_C_36 = 10'd513,
    COMP_LOOP_5_modExp_1_while_C_37 = 10'd514,
    COMP_LOOP_5_modExp_1_while_C_38 = 10'd515,
    COMP_LOOP_5_modExp_1_while_C_39 = 10'd516,
    COMP_LOOP_5_modExp_1_while_C_40 = 10'd517,
    COMP_LOOP_C_262 = 10'd518,
    COMP_LOOP_C_263 = 10'd519,
    COMP_LOOP_C_264 = 10'd520,
    COMP_LOOP_C_265 = 10'd521,
    COMP_LOOP_C_266 = 10'd522,
    COMP_LOOP_C_267 = 10'd523,
    COMP_LOOP_C_268 = 10'd524,
    COMP_LOOP_C_269 = 10'd525,
    COMP_LOOP_C_270 = 10'd526,
    COMP_LOOP_C_271 = 10'd527,
    COMP_LOOP_C_272 = 10'd528,
    COMP_LOOP_C_273 = 10'd529,
    COMP_LOOP_C_274 = 10'd530,
    COMP_LOOP_C_275 = 10'd531,
    COMP_LOOP_C_276 = 10'd532,
    COMP_LOOP_C_277 = 10'd533,
    COMP_LOOP_C_278 = 10'd534,
    COMP_LOOP_C_279 = 10'd535,
    COMP_LOOP_C_280 = 10'd536,
    COMP_LOOP_C_281 = 10'd537,
    COMP_LOOP_C_282 = 10'd538,
    COMP_LOOP_C_283 = 10'd539,
    COMP_LOOP_C_284 = 10'd540,
    COMP_LOOP_C_285 = 10'd541,
    COMP_LOOP_C_286 = 10'd542,
    COMP_LOOP_C_287 = 10'd543,
    COMP_LOOP_C_288 = 10'd544,
    COMP_LOOP_C_289 = 10'd545,
    COMP_LOOP_C_290 = 10'd546,
    COMP_LOOP_C_291 = 10'd547,
    COMP_LOOP_C_292 = 10'd548,
    COMP_LOOP_C_293 = 10'd549,
    COMP_LOOP_C_294 = 10'd550,
    COMP_LOOP_C_295 = 10'd551,
    COMP_LOOP_C_296 = 10'd552,
    COMP_LOOP_C_297 = 10'd553,
    COMP_LOOP_C_298 = 10'd554,
    COMP_LOOP_C_299 = 10'd555,
    COMP_LOOP_C_300 = 10'd556,
    COMP_LOOP_C_301 = 10'd557,
    COMP_LOOP_C_302 = 10'd558,
    COMP_LOOP_C_303 = 10'd559,
    COMP_LOOP_C_304 = 10'd560,
    COMP_LOOP_C_305 = 10'd561,
    COMP_LOOP_C_306 = 10'd562,
    COMP_LOOP_C_307 = 10'd563,
    COMP_LOOP_C_308 = 10'd564,
    COMP_LOOP_C_309 = 10'd565,
    COMP_LOOP_C_310 = 10'd566,
    COMP_LOOP_C_311 = 10'd567,
    COMP_LOOP_C_312 = 10'd568,
    COMP_LOOP_C_313 = 10'd569,
    COMP_LOOP_C_314 = 10'd570,
    COMP_LOOP_C_315 = 10'd571,
    COMP_LOOP_C_316 = 10'd572,
    COMP_LOOP_C_317 = 10'd573,
    COMP_LOOP_C_318 = 10'd574,
    COMP_LOOP_C_319 = 10'd575,
    COMP_LOOP_C_320 = 10'd576,
    COMP_LOOP_C_321 = 10'd577,
    COMP_LOOP_C_322 = 10'd578,
    COMP_LOOP_C_323 = 10'd579,
    COMP_LOOP_C_324 = 10'd580,
    COMP_LOOP_C_325 = 10'd581,
    COMP_LOOP_C_326 = 10'd582,
    COMP_LOOP_6_modExp_1_while_C_0 = 10'd583,
    COMP_LOOP_6_modExp_1_while_C_1 = 10'd584,
    COMP_LOOP_6_modExp_1_while_C_2 = 10'd585,
    COMP_LOOP_6_modExp_1_while_C_3 = 10'd586,
    COMP_LOOP_6_modExp_1_while_C_4 = 10'd587,
    COMP_LOOP_6_modExp_1_while_C_5 = 10'd588,
    COMP_LOOP_6_modExp_1_while_C_6 = 10'd589,
    COMP_LOOP_6_modExp_1_while_C_7 = 10'd590,
    COMP_LOOP_6_modExp_1_while_C_8 = 10'd591,
    COMP_LOOP_6_modExp_1_while_C_9 = 10'd592,
    COMP_LOOP_6_modExp_1_while_C_10 = 10'd593,
    COMP_LOOP_6_modExp_1_while_C_11 = 10'd594,
    COMP_LOOP_6_modExp_1_while_C_12 = 10'd595,
    COMP_LOOP_6_modExp_1_while_C_13 = 10'd596,
    COMP_LOOP_6_modExp_1_while_C_14 = 10'd597,
    COMP_LOOP_6_modExp_1_while_C_15 = 10'd598,
    COMP_LOOP_6_modExp_1_while_C_16 = 10'd599,
    COMP_LOOP_6_modExp_1_while_C_17 = 10'd600,
    COMP_LOOP_6_modExp_1_while_C_18 = 10'd601,
    COMP_LOOP_6_modExp_1_while_C_19 = 10'd602,
    COMP_LOOP_6_modExp_1_while_C_20 = 10'd603,
    COMP_LOOP_6_modExp_1_while_C_21 = 10'd604,
    COMP_LOOP_6_modExp_1_while_C_22 = 10'd605,
    COMP_LOOP_6_modExp_1_while_C_23 = 10'd606,
    COMP_LOOP_6_modExp_1_while_C_24 = 10'd607,
    COMP_LOOP_6_modExp_1_while_C_25 = 10'd608,
    COMP_LOOP_6_modExp_1_while_C_26 = 10'd609,
    COMP_LOOP_6_modExp_1_while_C_27 = 10'd610,
    COMP_LOOP_6_modExp_1_while_C_28 = 10'd611,
    COMP_LOOP_6_modExp_1_while_C_29 = 10'd612,
    COMP_LOOP_6_modExp_1_while_C_30 = 10'd613,
    COMP_LOOP_6_modExp_1_while_C_31 = 10'd614,
    COMP_LOOP_6_modExp_1_while_C_32 = 10'd615,
    COMP_LOOP_6_modExp_1_while_C_33 = 10'd616,
    COMP_LOOP_6_modExp_1_while_C_34 = 10'd617,
    COMP_LOOP_6_modExp_1_while_C_35 = 10'd618,
    COMP_LOOP_6_modExp_1_while_C_36 = 10'd619,
    COMP_LOOP_6_modExp_1_while_C_37 = 10'd620,
    COMP_LOOP_6_modExp_1_while_C_38 = 10'd621,
    COMP_LOOP_6_modExp_1_while_C_39 = 10'd622,
    COMP_LOOP_6_modExp_1_while_C_40 = 10'd623,
    COMP_LOOP_C_327 = 10'd624,
    COMP_LOOP_C_328 = 10'd625,
    COMP_LOOP_C_329 = 10'd626,
    COMP_LOOP_C_330 = 10'd627,
    COMP_LOOP_C_331 = 10'd628,
    COMP_LOOP_C_332 = 10'd629,
    COMP_LOOP_C_333 = 10'd630,
    COMP_LOOP_C_334 = 10'd631,
    COMP_LOOP_C_335 = 10'd632,
    COMP_LOOP_C_336 = 10'd633,
    COMP_LOOP_C_337 = 10'd634,
    COMP_LOOP_C_338 = 10'd635,
    COMP_LOOP_C_339 = 10'd636,
    COMP_LOOP_C_340 = 10'd637,
    COMP_LOOP_C_341 = 10'd638,
    COMP_LOOP_C_342 = 10'd639,
    COMP_LOOP_C_343 = 10'd640,
    COMP_LOOP_C_344 = 10'd641,
    COMP_LOOP_C_345 = 10'd642,
    COMP_LOOP_C_346 = 10'd643,
    COMP_LOOP_C_347 = 10'd644,
    COMP_LOOP_C_348 = 10'd645,
    COMP_LOOP_C_349 = 10'd646,
    COMP_LOOP_C_350 = 10'd647,
    COMP_LOOP_C_351 = 10'd648,
    COMP_LOOP_C_352 = 10'd649,
    COMP_LOOP_C_353 = 10'd650,
    COMP_LOOP_C_354 = 10'd651,
    COMP_LOOP_C_355 = 10'd652,
    COMP_LOOP_C_356 = 10'd653,
    COMP_LOOP_C_357 = 10'd654,
    COMP_LOOP_C_358 = 10'd655,
    COMP_LOOP_C_359 = 10'd656,
    COMP_LOOP_C_360 = 10'd657,
    COMP_LOOP_C_361 = 10'd658,
    COMP_LOOP_C_362 = 10'd659,
    COMP_LOOP_C_363 = 10'd660,
    COMP_LOOP_C_364 = 10'd661,
    COMP_LOOP_C_365 = 10'd662,
    COMP_LOOP_C_366 = 10'd663,
    COMP_LOOP_C_367 = 10'd664,
    COMP_LOOP_C_368 = 10'd665,
    COMP_LOOP_C_369 = 10'd666,
    COMP_LOOP_C_370 = 10'd667,
    COMP_LOOP_C_371 = 10'd668,
    COMP_LOOP_C_372 = 10'd669,
    COMP_LOOP_C_373 = 10'd670,
    COMP_LOOP_C_374 = 10'd671,
    COMP_LOOP_C_375 = 10'd672,
    COMP_LOOP_C_376 = 10'd673,
    COMP_LOOP_C_377 = 10'd674,
    COMP_LOOP_C_378 = 10'd675,
    COMP_LOOP_C_379 = 10'd676,
    COMP_LOOP_C_380 = 10'd677,
    COMP_LOOP_C_381 = 10'd678,
    COMP_LOOP_C_382 = 10'd679,
    COMP_LOOP_C_383 = 10'd680,
    COMP_LOOP_C_384 = 10'd681,
    COMP_LOOP_C_385 = 10'd682,
    COMP_LOOP_C_386 = 10'd683,
    COMP_LOOP_C_387 = 10'd684,
    COMP_LOOP_C_388 = 10'd685,
    COMP_LOOP_C_389 = 10'd686,
    COMP_LOOP_C_390 = 10'd687,
    COMP_LOOP_C_391 = 10'd688,
    COMP_LOOP_7_modExp_1_while_C_0 = 10'd689,
    COMP_LOOP_7_modExp_1_while_C_1 = 10'd690,
    COMP_LOOP_7_modExp_1_while_C_2 = 10'd691,
    COMP_LOOP_7_modExp_1_while_C_3 = 10'd692,
    COMP_LOOP_7_modExp_1_while_C_4 = 10'd693,
    COMP_LOOP_7_modExp_1_while_C_5 = 10'd694,
    COMP_LOOP_7_modExp_1_while_C_6 = 10'd695,
    COMP_LOOP_7_modExp_1_while_C_7 = 10'd696,
    COMP_LOOP_7_modExp_1_while_C_8 = 10'd697,
    COMP_LOOP_7_modExp_1_while_C_9 = 10'd698,
    COMP_LOOP_7_modExp_1_while_C_10 = 10'd699,
    COMP_LOOP_7_modExp_1_while_C_11 = 10'd700,
    COMP_LOOP_7_modExp_1_while_C_12 = 10'd701,
    COMP_LOOP_7_modExp_1_while_C_13 = 10'd702,
    COMP_LOOP_7_modExp_1_while_C_14 = 10'd703,
    COMP_LOOP_7_modExp_1_while_C_15 = 10'd704,
    COMP_LOOP_7_modExp_1_while_C_16 = 10'd705,
    COMP_LOOP_7_modExp_1_while_C_17 = 10'd706,
    COMP_LOOP_7_modExp_1_while_C_18 = 10'd707,
    COMP_LOOP_7_modExp_1_while_C_19 = 10'd708,
    COMP_LOOP_7_modExp_1_while_C_20 = 10'd709,
    COMP_LOOP_7_modExp_1_while_C_21 = 10'd710,
    COMP_LOOP_7_modExp_1_while_C_22 = 10'd711,
    COMP_LOOP_7_modExp_1_while_C_23 = 10'd712,
    COMP_LOOP_7_modExp_1_while_C_24 = 10'd713,
    COMP_LOOP_7_modExp_1_while_C_25 = 10'd714,
    COMP_LOOP_7_modExp_1_while_C_26 = 10'd715,
    COMP_LOOP_7_modExp_1_while_C_27 = 10'd716,
    COMP_LOOP_7_modExp_1_while_C_28 = 10'd717,
    COMP_LOOP_7_modExp_1_while_C_29 = 10'd718,
    COMP_LOOP_7_modExp_1_while_C_30 = 10'd719,
    COMP_LOOP_7_modExp_1_while_C_31 = 10'd720,
    COMP_LOOP_7_modExp_1_while_C_32 = 10'd721,
    COMP_LOOP_7_modExp_1_while_C_33 = 10'd722,
    COMP_LOOP_7_modExp_1_while_C_34 = 10'd723,
    COMP_LOOP_7_modExp_1_while_C_35 = 10'd724,
    COMP_LOOP_7_modExp_1_while_C_36 = 10'd725,
    COMP_LOOP_7_modExp_1_while_C_37 = 10'd726,
    COMP_LOOP_7_modExp_1_while_C_38 = 10'd727,
    COMP_LOOP_7_modExp_1_while_C_39 = 10'd728,
    COMP_LOOP_7_modExp_1_while_C_40 = 10'd729,
    COMP_LOOP_C_392 = 10'd730,
    COMP_LOOP_C_393 = 10'd731,
    COMP_LOOP_C_394 = 10'd732,
    COMP_LOOP_C_395 = 10'd733,
    COMP_LOOP_C_396 = 10'd734,
    COMP_LOOP_C_397 = 10'd735,
    COMP_LOOP_C_398 = 10'd736,
    COMP_LOOP_C_399 = 10'd737,
    COMP_LOOP_C_400 = 10'd738,
    COMP_LOOP_C_401 = 10'd739,
    COMP_LOOP_C_402 = 10'd740,
    COMP_LOOP_C_403 = 10'd741,
    COMP_LOOP_C_404 = 10'd742,
    COMP_LOOP_C_405 = 10'd743,
    COMP_LOOP_C_406 = 10'd744,
    COMP_LOOP_C_407 = 10'd745,
    COMP_LOOP_C_408 = 10'd746,
    COMP_LOOP_C_409 = 10'd747,
    COMP_LOOP_C_410 = 10'd748,
    COMP_LOOP_C_411 = 10'd749,
    COMP_LOOP_C_412 = 10'd750,
    COMP_LOOP_C_413 = 10'd751,
    COMP_LOOP_C_414 = 10'd752,
    COMP_LOOP_C_415 = 10'd753,
    COMP_LOOP_C_416 = 10'd754,
    COMP_LOOP_C_417 = 10'd755,
    COMP_LOOP_C_418 = 10'd756,
    COMP_LOOP_C_419 = 10'd757,
    COMP_LOOP_C_420 = 10'd758,
    COMP_LOOP_C_421 = 10'd759,
    COMP_LOOP_C_422 = 10'd760,
    COMP_LOOP_C_423 = 10'd761,
    COMP_LOOP_C_424 = 10'd762,
    COMP_LOOP_C_425 = 10'd763,
    COMP_LOOP_C_426 = 10'd764,
    COMP_LOOP_C_427 = 10'd765,
    COMP_LOOP_C_428 = 10'd766,
    COMP_LOOP_C_429 = 10'd767,
    COMP_LOOP_C_430 = 10'd768,
    COMP_LOOP_C_431 = 10'd769,
    COMP_LOOP_C_432 = 10'd770,
    COMP_LOOP_C_433 = 10'd771,
    COMP_LOOP_C_434 = 10'd772,
    COMP_LOOP_C_435 = 10'd773,
    COMP_LOOP_C_436 = 10'd774,
    COMP_LOOP_C_437 = 10'd775,
    COMP_LOOP_C_438 = 10'd776,
    COMP_LOOP_C_439 = 10'd777,
    COMP_LOOP_C_440 = 10'd778,
    COMP_LOOP_C_441 = 10'd779,
    COMP_LOOP_C_442 = 10'd780,
    COMP_LOOP_C_443 = 10'd781,
    COMP_LOOP_C_444 = 10'd782,
    COMP_LOOP_C_445 = 10'd783,
    COMP_LOOP_C_446 = 10'd784,
    COMP_LOOP_C_447 = 10'd785,
    COMP_LOOP_C_448 = 10'd786,
    COMP_LOOP_C_449 = 10'd787,
    COMP_LOOP_C_450 = 10'd788,
    COMP_LOOP_C_451 = 10'd789,
    COMP_LOOP_C_452 = 10'd790,
    COMP_LOOP_C_453 = 10'd791,
    COMP_LOOP_C_454 = 10'd792,
    COMP_LOOP_C_455 = 10'd793,
    COMP_LOOP_C_456 = 10'd794,
    COMP_LOOP_8_modExp_1_while_C_0 = 10'd795,
    COMP_LOOP_8_modExp_1_while_C_1 = 10'd796,
    COMP_LOOP_8_modExp_1_while_C_2 = 10'd797,
    COMP_LOOP_8_modExp_1_while_C_3 = 10'd798,
    COMP_LOOP_8_modExp_1_while_C_4 = 10'd799,
    COMP_LOOP_8_modExp_1_while_C_5 = 10'd800,
    COMP_LOOP_8_modExp_1_while_C_6 = 10'd801,
    COMP_LOOP_8_modExp_1_while_C_7 = 10'd802,
    COMP_LOOP_8_modExp_1_while_C_8 = 10'd803,
    COMP_LOOP_8_modExp_1_while_C_9 = 10'd804,
    COMP_LOOP_8_modExp_1_while_C_10 = 10'd805,
    COMP_LOOP_8_modExp_1_while_C_11 = 10'd806,
    COMP_LOOP_8_modExp_1_while_C_12 = 10'd807,
    COMP_LOOP_8_modExp_1_while_C_13 = 10'd808,
    COMP_LOOP_8_modExp_1_while_C_14 = 10'd809,
    COMP_LOOP_8_modExp_1_while_C_15 = 10'd810,
    COMP_LOOP_8_modExp_1_while_C_16 = 10'd811,
    COMP_LOOP_8_modExp_1_while_C_17 = 10'd812,
    COMP_LOOP_8_modExp_1_while_C_18 = 10'd813,
    COMP_LOOP_8_modExp_1_while_C_19 = 10'd814,
    COMP_LOOP_8_modExp_1_while_C_20 = 10'd815,
    COMP_LOOP_8_modExp_1_while_C_21 = 10'd816,
    COMP_LOOP_8_modExp_1_while_C_22 = 10'd817,
    COMP_LOOP_8_modExp_1_while_C_23 = 10'd818,
    COMP_LOOP_8_modExp_1_while_C_24 = 10'd819,
    COMP_LOOP_8_modExp_1_while_C_25 = 10'd820,
    COMP_LOOP_8_modExp_1_while_C_26 = 10'd821,
    COMP_LOOP_8_modExp_1_while_C_27 = 10'd822,
    COMP_LOOP_8_modExp_1_while_C_28 = 10'd823,
    COMP_LOOP_8_modExp_1_while_C_29 = 10'd824,
    COMP_LOOP_8_modExp_1_while_C_30 = 10'd825,
    COMP_LOOP_8_modExp_1_while_C_31 = 10'd826,
    COMP_LOOP_8_modExp_1_while_C_32 = 10'd827,
    COMP_LOOP_8_modExp_1_while_C_33 = 10'd828,
    COMP_LOOP_8_modExp_1_while_C_34 = 10'd829,
    COMP_LOOP_8_modExp_1_while_C_35 = 10'd830,
    COMP_LOOP_8_modExp_1_while_C_36 = 10'd831,
    COMP_LOOP_8_modExp_1_while_C_37 = 10'd832,
    COMP_LOOP_8_modExp_1_while_C_38 = 10'd833,
    COMP_LOOP_8_modExp_1_while_C_39 = 10'd834,
    COMP_LOOP_8_modExp_1_while_C_40 = 10'd835,
    COMP_LOOP_C_457 = 10'd836,
    COMP_LOOP_C_458 = 10'd837,
    COMP_LOOP_C_459 = 10'd838,
    COMP_LOOP_C_460 = 10'd839,
    COMP_LOOP_C_461 = 10'd840,
    COMP_LOOP_C_462 = 10'd841,
    COMP_LOOP_C_463 = 10'd842,
    COMP_LOOP_C_464 = 10'd843,
    COMP_LOOP_C_465 = 10'd844,
    COMP_LOOP_C_466 = 10'd845,
    COMP_LOOP_C_467 = 10'd846,
    COMP_LOOP_C_468 = 10'd847,
    COMP_LOOP_C_469 = 10'd848,
    COMP_LOOP_C_470 = 10'd849,
    COMP_LOOP_C_471 = 10'd850,
    COMP_LOOP_C_472 = 10'd851,
    COMP_LOOP_C_473 = 10'd852,
    COMP_LOOP_C_474 = 10'd853,
    COMP_LOOP_C_475 = 10'd854,
    COMP_LOOP_C_476 = 10'd855,
    COMP_LOOP_C_477 = 10'd856,
    COMP_LOOP_C_478 = 10'd857,
    COMP_LOOP_C_479 = 10'd858,
    COMP_LOOP_C_480 = 10'd859,
    COMP_LOOP_C_481 = 10'd860,
    COMP_LOOP_C_482 = 10'd861,
    COMP_LOOP_C_483 = 10'd862,
    COMP_LOOP_C_484 = 10'd863,
    COMP_LOOP_C_485 = 10'd864,
    COMP_LOOP_C_486 = 10'd865,
    COMP_LOOP_C_487 = 10'd866,
    COMP_LOOP_C_488 = 10'd867,
    COMP_LOOP_C_489 = 10'd868,
    COMP_LOOP_C_490 = 10'd869,
    COMP_LOOP_C_491 = 10'd870,
    COMP_LOOP_C_492 = 10'd871,
    COMP_LOOP_C_493 = 10'd872,
    COMP_LOOP_C_494 = 10'd873,
    COMP_LOOP_C_495 = 10'd874,
    COMP_LOOP_C_496 = 10'd875,
    COMP_LOOP_C_497 = 10'd876,
    COMP_LOOP_C_498 = 10'd877,
    COMP_LOOP_C_499 = 10'd878,
    COMP_LOOP_C_500 = 10'd879,
    COMP_LOOP_C_501 = 10'd880,
    COMP_LOOP_C_502 = 10'd881,
    COMP_LOOP_C_503 = 10'd882,
    COMP_LOOP_C_504 = 10'd883,
    COMP_LOOP_C_505 = 10'd884,
    COMP_LOOP_C_506 = 10'd885,
    COMP_LOOP_C_507 = 10'd886,
    COMP_LOOP_C_508 = 10'd887,
    COMP_LOOP_C_509 = 10'd888,
    COMP_LOOP_C_510 = 10'd889,
    COMP_LOOP_C_511 = 10'd890,
    COMP_LOOP_C_512 = 10'd891,
    COMP_LOOP_C_513 = 10'd892,
    COMP_LOOP_C_514 = 10'd893,
    COMP_LOOP_C_515 = 10'd894,
    COMP_LOOP_C_516 = 10'd895,
    COMP_LOOP_C_517 = 10'd896,
    COMP_LOOP_C_518 = 10'd897,
    COMP_LOOP_C_519 = 10'd898,
    COMP_LOOP_C_520 = 10'd899,
    VEC_LOOP_C_0 = 10'd900,
    STAGE_LOOP_C_9 = 10'd901,
    main_C_1 = 10'd902;

  reg [9:0] state_var;
  reg [9:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 10'b0000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 10'b0000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 10'b0000000100;
        state_var_NS = STAGE_LOOP_C_4;
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 10'b0000000101;
        state_var_NS = STAGE_LOOP_C_5;
      end
      STAGE_LOOP_C_5 : begin
        fsm_output = 10'b0000000110;
        state_var_NS = STAGE_LOOP_C_6;
      end
      STAGE_LOOP_C_6 : begin
        fsm_output = 10'b0000000111;
        state_var_NS = STAGE_LOOP_C_7;
      end
      STAGE_LOOP_C_7 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = STAGE_LOOP_C_8;
      end
      STAGE_LOOP_C_8 : begin
        fsm_output = 10'b0000001001;
        if ( STAGE_LOOP_C_8_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      modExp_while_C_0 : begin
        fsm_output = 10'b0000001010;
        state_var_NS = modExp_while_C_1;
      end
      modExp_while_C_1 : begin
        fsm_output = 10'b0000001011;
        state_var_NS = modExp_while_C_2;
      end
      modExp_while_C_2 : begin
        fsm_output = 10'b0000001100;
        state_var_NS = modExp_while_C_3;
      end
      modExp_while_C_3 : begin
        fsm_output = 10'b0000001101;
        state_var_NS = modExp_while_C_4;
      end
      modExp_while_C_4 : begin
        fsm_output = 10'b0000001110;
        state_var_NS = modExp_while_C_5;
      end
      modExp_while_C_5 : begin
        fsm_output = 10'b0000001111;
        state_var_NS = modExp_while_C_6;
      end
      modExp_while_C_6 : begin
        fsm_output = 10'b0000010000;
        state_var_NS = modExp_while_C_7;
      end
      modExp_while_C_7 : begin
        fsm_output = 10'b0000010001;
        state_var_NS = modExp_while_C_8;
      end
      modExp_while_C_8 : begin
        fsm_output = 10'b0000010010;
        state_var_NS = modExp_while_C_9;
      end
      modExp_while_C_9 : begin
        fsm_output = 10'b0000010011;
        state_var_NS = modExp_while_C_10;
      end
      modExp_while_C_10 : begin
        fsm_output = 10'b0000010100;
        state_var_NS = modExp_while_C_11;
      end
      modExp_while_C_11 : begin
        fsm_output = 10'b0000010101;
        state_var_NS = modExp_while_C_12;
      end
      modExp_while_C_12 : begin
        fsm_output = 10'b0000010110;
        state_var_NS = modExp_while_C_13;
      end
      modExp_while_C_13 : begin
        fsm_output = 10'b0000010111;
        state_var_NS = modExp_while_C_14;
      end
      modExp_while_C_14 : begin
        fsm_output = 10'b0000011000;
        state_var_NS = modExp_while_C_15;
      end
      modExp_while_C_15 : begin
        fsm_output = 10'b0000011001;
        state_var_NS = modExp_while_C_16;
      end
      modExp_while_C_16 : begin
        fsm_output = 10'b0000011010;
        state_var_NS = modExp_while_C_17;
      end
      modExp_while_C_17 : begin
        fsm_output = 10'b0000011011;
        state_var_NS = modExp_while_C_18;
      end
      modExp_while_C_18 : begin
        fsm_output = 10'b0000011100;
        state_var_NS = modExp_while_C_19;
      end
      modExp_while_C_19 : begin
        fsm_output = 10'b0000011101;
        state_var_NS = modExp_while_C_20;
      end
      modExp_while_C_20 : begin
        fsm_output = 10'b0000011110;
        state_var_NS = modExp_while_C_21;
      end
      modExp_while_C_21 : begin
        fsm_output = 10'b0000011111;
        state_var_NS = modExp_while_C_22;
      end
      modExp_while_C_22 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = modExp_while_C_23;
      end
      modExp_while_C_23 : begin
        fsm_output = 10'b0000100001;
        state_var_NS = modExp_while_C_24;
      end
      modExp_while_C_24 : begin
        fsm_output = 10'b0000100010;
        state_var_NS = modExp_while_C_25;
      end
      modExp_while_C_25 : begin
        fsm_output = 10'b0000100011;
        state_var_NS = modExp_while_C_26;
      end
      modExp_while_C_26 : begin
        fsm_output = 10'b0000100100;
        state_var_NS = modExp_while_C_27;
      end
      modExp_while_C_27 : begin
        fsm_output = 10'b0000100101;
        state_var_NS = modExp_while_C_28;
      end
      modExp_while_C_28 : begin
        fsm_output = 10'b0000100110;
        state_var_NS = modExp_while_C_29;
      end
      modExp_while_C_29 : begin
        fsm_output = 10'b0000100111;
        state_var_NS = modExp_while_C_30;
      end
      modExp_while_C_30 : begin
        fsm_output = 10'b0000101000;
        state_var_NS = modExp_while_C_31;
      end
      modExp_while_C_31 : begin
        fsm_output = 10'b0000101001;
        state_var_NS = modExp_while_C_32;
      end
      modExp_while_C_32 : begin
        fsm_output = 10'b0000101010;
        state_var_NS = modExp_while_C_33;
      end
      modExp_while_C_33 : begin
        fsm_output = 10'b0000101011;
        state_var_NS = modExp_while_C_34;
      end
      modExp_while_C_34 : begin
        fsm_output = 10'b0000101100;
        state_var_NS = modExp_while_C_35;
      end
      modExp_while_C_35 : begin
        fsm_output = 10'b0000101101;
        state_var_NS = modExp_while_C_36;
      end
      modExp_while_C_36 : begin
        fsm_output = 10'b0000101110;
        state_var_NS = modExp_while_C_37;
      end
      modExp_while_C_37 : begin
        fsm_output = 10'b0000101111;
        state_var_NS = modExp_while_C_38;
      end
      modExp_while_C_38 : begin
        fsm_output = 10'b0000110000;
        state_var_NS = modExp_while_C_39;
      end
      modExp_while_C_39 : begin
        fsm_output = 10'b0000110001;
        state_var_NS = modExp_while_C_40;
      end
      modExp_while_C_40 : begin
        fsm_output = 10'b0000110010;
        if ( modExp_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 10'b0000110011;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 10'b0000110100;
        if ( COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 10'b0000110101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_1;
      end
      COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 10'b0000110110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_2;
      end
      COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 10'b0000110111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_3;
      end
      COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 10'b0000111000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_4;
      end
      COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 10'b0000111001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_5;
      end
      COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 10'b0000111010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_6;
      end
      COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 10'b0000111011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_7;
      end
      COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 10'b0000111100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_8;
      end
      COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 10'b0000111101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_9;
      end
      COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 10'b0000111110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_10;
      end
      COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 10'b0000111111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_11;
      end
      COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_12;
      end
      COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 10'b0001000001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_13;
      end
      COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 10'b0001000010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_14;
      end
      COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 10'b0001000011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_15;
      end
      COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 10'b0001000100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_16;
      end
      COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 10'b0001000101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_17;
      end
      COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 10'b0001000110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_18;
      end
      COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 10'b0001000111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_19;
      end
      COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 10'b0001001000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_20;
      end
      COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 10'b0001001001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_21;
      end
      COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 10'b0001001010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_22;
      end
      COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 10'b0001001011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_23;
      end
      COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 10'b0001001100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_24;
      end
      COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 10'b0001001101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_25;
      end
      COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 10'b0001001110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_26;
      end
      COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 10'b0001001111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_27;
      end
      COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 10'b0001010000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_28;
      end
      COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 10'b0001010001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_29;
      end
      COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 10'b0001010010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_30;
      end
      COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 10'b0001010011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_31;
      end
      COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 10'b0001010100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_32;
      end
      COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 10'b0001010101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_33;
      end
      COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 10'b0001010110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_34;
      end
      COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 10'b0001010111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_35;
      end
      COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 10'b0001011000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_36;
      end
      COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 10'b0001011001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_37;
      end
      COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 10'b0001011010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_38;
      end
      COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 10'b0001011011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_39;
      end
      COMP_LOOP_1_modExp_1_while_C_39 : begin
        fsm_output = 10'b0001011100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_40;
      end
      COMP_LOOP_1_modExp_1_while_C_40 : begin
        fsm_output = 10'b0001011101;
        if ( COMP_LOOP_1_modExp_1_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 10'b0001011110;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 10'b0001011111;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 10'b0001100000;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 10'b0001100001;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 10'b0001100010;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 10'b0001100011;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 10'b0001100100;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 10'b0001100101;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 10'b0001100110;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 10'b0001100111;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 10'b0001101000;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 10'b0001101001;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 10'b0001101010;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 10'b0001101011;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 10'b0001101100;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 10'b0001101101;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 10'b0001101110;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 10'b0001101111;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 10'b0001110000;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 10'b0001110001;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 10'b0001110010;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 10'b0001110011;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 10'b0001110100;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 10'b0001110101;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 10'b0001110110;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 10'b0001110111;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 10'b0001111000;
        state_var_NS = COMP_LOOP_C_29;
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 10'b0001111001;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 10'b0001111010;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 10'b0001111011;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 10'b0001111100;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 10'b0001111101;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 10'b0001111110;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 10'b0001111111;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 10'b0010000000;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 10'b0010000001;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 10'b0010000010;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 10'b0010000011;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 10'b0010000100;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 10'b0010000101;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 10'b0010000110;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 10'b0010000111;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 10'b0010001000;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 10'b0010001001;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 10'b0010001010;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 10'b0010001011;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 10'b0010001100;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 10'b0010001101;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 10'b0010001110;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 10'b0010001111;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 10'b0010010000;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 10'b0010010001;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 10'b0010010010;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 10'b0010010011;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 10'b0010010100;
        state_var_NS = COMP_LOOP_C_57;
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 10'b0010010101;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 10'b0010010110;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 10'b0010010111;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 10'b0010011000;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 10'b0010011001;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 10'b0010011010;
        state_var_NS = COMP_LOOP_C_63;
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 10'b0010011011;
        state_var_NS = COMP_LOOP_C_64;
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 10'b0010011100;
        state_var_NS = COMP_LOOP_C_65;
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 10'b0010011101;
        if ( COMP_LOOP_C_65_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_66;
        end
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 10'b0010011110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
      end
      COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 10'b0010011111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_1;
      end
      COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 10'b0010100000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_2;
      end
      COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 10'b0010100001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_3;
      end
      COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 10'b0010100010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_4;
      end
      COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 10'b0010100011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_5;
      end
      COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 10'b0010100100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_6;
      end
      COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 10'b0010100101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_7;
      end
      COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 10'b0010100110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_8;
      end
      COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 10'b0010100111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_9;
      end
      COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 10'b0010101000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_10;
      end
      COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 10'b0010101001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_11;
      end
      COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 10'b0010101010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_12;
      end
      COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 10'b0010101011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_13;
      end
      COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 10'b0010101100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_14;
      end
      COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 10'b0010101101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_15;
      end
      COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 10'b0010101110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_16;
      end
      COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 10'b0010101111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_17;
      end
      COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 10'b0010110000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_18;
      end
      COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 10'b0010110001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_19;
      end
      COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 10'b0010110010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_20;
      end
      COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 10'b0010110011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_21;
      end
      COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 10'b0010110100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_22;
      end
      COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 10'b0010110101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_23;
      end
      COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 10'b0010110110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_24;
      end
      COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 10'b0010110111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_25;
      end
      COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 10'b0010111000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_26;
      end
      COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 10'b0010111001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_27;
      end
      COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 10'b0010111010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_28;
      end
      COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 10'b0010111011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_29;
      end
      COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 10'b0010111100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_30;
      end
      COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 10'b0010111101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_31;
      end
      COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 10'b0010111110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_32;
      end
      COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 10'b0010111111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_33;
      end
      COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 10'b0011000000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_34;
      end
      COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 10'b0011000001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_35;
      end
      COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 10'b0011000010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_36;
      end
      COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 10'b0011000011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_37;
      end
      COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 10'b0011000100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_38;
      end
      COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 10'b0011000101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_39;
      end
      COMP_LOOP_2_modExp_1_while_C_39 : begin
        fsm_output = 10'b0011000110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_40;
      end
      COMP_LOOP_2_modExp_1_while_C_40 : begin
        fsm_output = 10'b0011000111;
        if ( COMP_LOOP_2_modExp_1_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_67;
        end
        else begin
          state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 10'b0011001000;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 10'b0011001001;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 10'b0011001010;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 10'b0011001011;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 10'b0011001100;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 10'b0011001101;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 10'b0011001110;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 10'b0011001111;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 10'b0011010000;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 10'b0011010001;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 10'b0011010010;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 10'b0011010011;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 10'b0011010100;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 10'b0011010101;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 10'b0011010110;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 10'b0011010111;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 10'b0011011000;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 10'b0011011001;
        state_var_NS = COMP_LOOP_C_85;
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 10'b0011011010;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 10'b0011011011;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 10'b0011011100;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 10'b0011011101;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 10'b0011011110;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 10'b0011011111;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 10'b0011100000;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 10'b0011100001;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 10'b0011100010;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 10'b0011100011;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 10'b0011100100;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 10'b0011100101;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 10'b0011100110;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 10'b0011100111;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 10'b0011101000;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 10'b0011101001;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 10'b0011101010;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 10'b0011101011;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 10'b0011101100;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 10'b0011101101;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 10'b0011101110;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 10'b0011101111;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 10'b0011110000;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 10'b0011110001;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 10'b0011110010;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 10'b0011110011;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 10'b0011110100;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 10'b0011110101;
        state_var_NS = COMP_LOOP_C_113;
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 10'b0011110110;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 10'b0011110111;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 10'b0011111000;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 10'b0011111001;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 10'b0011111010;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 10'b0011111011;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 10'b0011111100;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 10'b0011111101;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 10'b0011111110;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 10'b0011111111;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 10'b0100000001;
        state_var_NS = COMP_LOOP_C_125;
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 10'b0100000010;
        state_var_NS = COMP_LOOP_C_126;
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 10'b0100000011;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 10'b0100000100;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 10'b0100000101;
        state_var_NS = COMP_LOOP_C_129;
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 10'b0100000110;
        state_var_NS = COMP_LOOP_C_130;
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 10'b0100000111;
        if ( COMP_LOOP_C_130_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_131;
        end
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 10'b0100001000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
      end
      COMP_LOOP_3_modExp_1_while_C_0 : begin
        fsm_output = 10'b0100001001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_1;
      end
      COMP_LOOP_3_modExp_1_while_C_1 : begin
        fsm_output = 10'b0100001010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_2;
      end
      COMP_LOOP_3_modExp_1_while_C_2 : begin
        fsm_output = 10'b0100001011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_3;
      end
      COMP_LOOP_3_modExp_1_while_C_3 : begin
        fsm_output = 10'b0100001100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_4;
      end
      COMP_LOOP_3_modExp_1_while_C_4 : begin
        fsm_output = 10'b0100001101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_5;
      end
      COMP_LOOP_3_modExp_1_while_C_5 : begin
        fsm_output = 10'b0100001110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_6;
      end
      COMP_LOOP_3_modExp_1_while_C_6 : begin
        fsm_output = 10'b0100001111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_7;
      end
      COMP_LOOP_3_modExp_1_while_C_7 : begin
        fsm_output = 10'b0100010000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_8;
      end
      COMP_LOOP_3_modExp_1_while_C_8 : begin
        fsm_output = 10'b0100010001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_9;
      end
      COMP_LOOP_3_modExp_1_while_C_9 : begin
        fsm_output = 10'b0100010010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_10;
      end
      COMP_LOOP_3_modExp_1_while_C_10 : begin
        fsm_output = 10'b0100010011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_11;
      end
      COMP_LOOP_3_modExp_1_while_C_11 : begin
        fsm_output = 10'b0100010100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_12;
      end
      COMP_LOOP_3_modExp_1_while_C_12 : begin
        fsm_output = 10'b0100010101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_13;
      end
      COMP_LOOP_3_modExp_1_while_C_13 : begin
        fsm_output = 10'b0100010110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_14;
      end
      COMP_LOOP_3_modExp_1_while_C_14 : begin
        fsm_output = 10'b0100010111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_15;
      end
      COMP_LOOP_3_modExp_1_while_C_15 : begin
        fsm_output = 10'b0100011000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_16;
      end
      COMP_LOOP_3_modExp_1_while_C_16 : begin
        fsm_output = 10'b0100011001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_17;
      end
      COMP_LOOP_3_modExp_1_while_C_17 : begin
        fsm_output = 10'b0100011010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_18;
      end
      COMP_LOOP_3_modExp_1_while_C_18 : begin
        fsm_output = 10'b0100011011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_19;
      end
      COMP_LOOP_3_modExp_1_while_C_19 : begin
        fsm_output = 10'b0100011100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_20;
      end
      COMP_LOOP_3_modExp_1_while_C_20 : begin
        fsm_output = 10'b0100011101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_21;
      end
      COMP_LOOP_3_modExp_1_while_C_21 : begin
        fsm_output = 10'b0100011110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_22;
      end
      COMP_LOOP_3_modExp_1_while_C_22 : begin
        fsm_output = 10'b0100011111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_23;
      end
      COMP_LOOP_3_modExp_1_while_C_23 : begin
        fsm_output = 10'b0100100000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_24;
      end
      COMP_LOOP_3_modExp_1_while_C_24 : begin
        fsm_output = 10'b0100100001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_25;
      end
      COMP_LOOP_3_modExp_1_while_C_25 : begin
        fsm_output = 10'b0100100010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_26;
      end
      COMP_LOOP_3_modExp_1_while_C_26 : begin
        fsm_output = 10'b0100100011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_27;
      end
      COMP_LOOP_3_modExp_1_while_C_27 : begin
        fsm_output = 10'b0100100100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_28;
      end
      COMP_LOOP_3_modExp_1_while_C_28 : begin
        fsm_output = 10'b0100100101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_29;
      end
      COMP_LOOP_3_modExp_1_while_C_29 : begin
        fsm_output = 10'b0100100110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_30;
      end
      COMP_LOOP_3_modExp_1_while_C_30 : begin
        fsm_output = 10'b0100100111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_31;
      end
      COMP_LOOP_3_modExp_1_while_C_31 : begin
        fsm_output = 10'b0100101000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_32;
      end
      COMP_LOOP_3_modExp_1_while_C_32 : begin
        fsm_output = 10'b0100101001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_33;
      end
      COMP_LOOP_3_modExp_1_while_C_33 : begin
        fsm_output = 10'b0100101010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_34;
      end
      COMP_LOOP_3_modExp_1_while_C_34 : begin
        fsm_output = 10'b0100101011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_35;
      end
      COMP_LOOP_3_modExp_1_while_C_35 : begin
        fsm_output = 10'b0100101100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_36;
      end
      COMP_LOOP_3_modExp_1_while_C_36 : begin
        fsm_output = 10'b0100101101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_37;
      end
      COMP_LOOP_3_modExp_1_while_C_37 : begin
        fsm_output = 10'b0100101110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_38;
      end
      COMP_LOOP_3_modExp_1_while_C_38 : begin
        fsm_output = 10'b0100101111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_39;
      end
      COMP_LOOP_3_modExp_1_while_C_39 : begin
        fsm_output = 10'b0100110000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_40;
      end
      COMP_LOOP_3_modExp_1_while_C_40 : begin
        fsm_output = 10'b0100110001;
        if ( COMP_LOOP_3_modExp_1_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_132;
        end
        else begin
          state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 10'b0100110010;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 10'b0100110011;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 10'b0100110100;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 10'b0100110101;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 10'b0100110110;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 10'b0100110111;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 10'b0100111000;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 10'b0100111001;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 10'b0100111010;
        state_var_NS = COMP_LOOP_C_141;
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 10'b0100111011;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 10'b0100111100;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 10'b0100111101;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 10'b0100111110;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 10'b0100111111;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 10'b0101000000;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 10'b0101000001;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 10'b0101000010;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 10'b0101000011;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 10'b0101000100;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 10'b0101000101;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 10'b0101000110;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 10'b0101000111;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 10'b0101001000;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 10'b0101001001;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 10'b0101001010;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 10'b0101001011;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 10'b0101001100;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 10'b0101001101;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 10'b0101001110;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 10'b0101001111;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 10'b0101010000;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 10'b0101010001;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 10'b0101010010;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 10'b0101010011;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 10'b0101010100;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 10'b0101010101;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 10'b0101010110;
        state_var_NS = COMP_LOOP_C_169;
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 10'b0101010111;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 10'b0101011000;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 10'b0101011001;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 10'b0101011010;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 10'b0101011011;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 10'b0101011100;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 10'b0101011101;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 10'b0101011110;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 10'b0101011111;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 10'b0101100000;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 10'b0101100001;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 10'b0101100010;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 10'b0101100011;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 10'b0101100100;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 10'b0101100101;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 10'b0101100110;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 10'b0101100111;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 10'b0101101000;
        state_var_NS = COMP_LOOP_C_187;
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 10'b0101101001;
        state_var_NS = COMP_LOOP_C_188;
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 10'b0101101010;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 10'b0101101011;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 10'b0101101100;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 10'b0101101101;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 10'b0101101110;
        state_var_NS = COMP_LOOP_C_193;
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 10'b0101101111;
        state_var_NS = COMP_LOOP_C_194;
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 10'b0101110000;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 10'b0101110001;
        if ( COMP_LOOP_C_195_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_196;
        end
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 10'b0101110010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
      end
      COMP_LOOP_4_modExp_1_while_C_0 : begin
        fsm_output = 10'b0101110011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_1;
      end
      COMP_LOOP_4_modExp_1_while_C_1 : begin
        fsm_output = 10'b0101110100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_2;
      end
      COMP_LOOP_4_modExp_1_while_C_2 : begin
        fsm_output = 10'b0101110101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_3;
      end
      COMP_LOOP_4_modExp_1_while_C_3 : begin
        fsm_output = 10'b0101110110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_4;
      end
      COMP_LOOP_4_modExp_1_while_C_4 : begin
        fsm_output = 10'b0101110111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_5;
      end
      COMP_LOOP_4_modExp_1_while_C_5 : begin
        fsm_output = 10'b0101111000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_6;
      end
      COMP_LOOP_4_modExp_1_while_C_6 : begin
        fsm_output = 10'b0101111001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_7;
      end
      COMP_LOOP_4_modExp_1_while_C_7 : begin
        fsm_output = 10'b0101111010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_8;
      end
      COMP_LOOP_4_modExp_1_while_C_8 : begin
        fsm_output = 10'b0101111011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_9;
      end
      COMP_LOOP_4_modExp_1_while_C_9 : begin
        fsm_output = 10'b0101111100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_10;
      end
      COMP_LOOP_4_modExp_1_while_C_10 : begin
        fsm_output = 10'b0101111101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_11;
      end
      COMP_LOOP_4_modExp_1_while_C_11 : begin
        fsm_output = 10'b0101111110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_12;
      end
      COMP_LOOP_4_modExp_1_while_C_12 : begin
        fsm_output = 10'b0101111111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_13;
      end
      COMP_LOOP_4_modExp_1_while_C_13 : begin
        fsm_output = 10'b0110000000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_14;
      end
      COMP_LOOP_4_modExp_1_while_C_14 : begin
        fsm_output = 10'b0110000001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_15;
      end
      COMP_LOOP_4_modExp_1_while_C_15 : begin
        fsm_output = 10'b0110000010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_16;
      end
      COMP_LOOP_4_modExp_1_while_C_16 : begin
        fsm_output = 10'b0110000011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_17;
      end
      COMP_LOOP_4_modExp_1_while_C_17 : begin
        fsm_output = 10'b0110000100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_18;
      end
      COMP_LOOP_4_modExp_1_while_C_18 : begin
        fsm_output = 10'b0110000101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_19;
      end
      COMP_LOOP_4_modExp_1_while_C_19 : begin
        fsm_output = 10'b0110000110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_20;
      end
      COMP_LOOP_4_modExp_1_while_C_20 : begin
        fsm_output = 10'b0110000111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_21;
      end
      COMP_LOOP_4_modExp_1_while_C_21 : begin
        fsm_output = 10'b0110001000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_22;
      end
      COMP_LOOP_4_modExp_1_while_C_22 : begin
        fsm_output = 10'b0110001001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_23;
      end
      COMP_LOOP_4_modExp_1_while_C_23 : begin
        fsm_output = 10'b0110001010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_24;
      end
      COMP_LOOP_4_modExp_1_while_C_24 : begin
        fsm_output = 10'b0110001011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_25;
      end
      COMP_LOOP_4_modExp_1_while_C_25 : begin
        fsm_output = 10'b0110001100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_26;
      end
      COMP_LOOP_4_modExp_1_while_C_26 : begin
        fsm_output = 10'b0110001101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_27;
      end
      COMP_LOOP_4_modExp_1_while_C_27 : begin
        fsm_output = 10'b0110001110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_28;
      end
      COMP_LOOP_4_modExp_1_while_C_28 : begin
        fsm_output = 10'b0110001111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_29;
      end
      COMP_LOOP_4_modExp_1_while_C_29 : begin
        fsm_output = 10'b0110010000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_30;
      end
      COMP_LOOP_4_modExp_1_while_C_30 : begin
        fsm_output = 10'b0110010001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_31;
      end
      COMP_LOOP_4_modExp_1_while_C_31 : begin
        fsm_output = 10'b0110010010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_32;
      end
      COMP_LOOP_4_modExp_1_while_C_32 : begin
        fsm_output = 10'b0110010011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_33;
      end
      COMP_LOOP_4_modExp_1_while_C_33 : begin
        fsm_output = 10'b0110010100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_34;
      end
      COMP_LOOP_4_modExp_1_while_C_34 : begin
        fsm_output = 10'b0110010101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_35;
      end
      COMP_LOOP_4_modExp_1_while_C_35 : begin
        fsm_output = 10'b0110010110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_36;
      end
      COMP_LOOP_4_modExp_1_while_C_36 : begin
        fsm_output = 10'b0110010111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_37;
      end
      COMP_LOOP_4_modExp_1_while_C_37 : begin
        fsm_output = 10'b0110011000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_38;
      end
      COMP_LOOP_4_modExp_1_while_C_38 : begin
        fsm_output = 10'b0110011001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_39;
      end
      COMP_LOOP_4_modExp_1_while_C_39 : begin
        fsm_output = 10'b0110011010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_40;
      end
      COMP_LOOP_4_modExp_1_while_C_40 : begin
        fsm_output = 10'b0110011011;
        if ( COMP_LOOP_4_modExp_1_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_197;
        end
        else begin
          state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 10'b0110011100;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 10'b0110011101;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 10'b0110011110;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 10'b0110011111;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 10'b0110100000;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 10'b0110100001;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 10'b0110100010;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 10'b0110100011;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 10'b0110100100;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 10'b0110100101;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 10'b0110100110;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 10'b0110100111;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 10'b0110101000;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 10'b0110101001;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 10'b0110101010;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 10'b0110101011;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 10'b0110101100;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 10'b0110101101;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 10'b0110101110;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 10'b0110101111;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 10'b0110110000;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 10'b0110110001;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 10'b0110110010;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 10'b0110110011;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 10'b0110110100;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 10'b0110110101;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 10'b0110110110;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 10'b0110110111;
        state_var_NS = COMP_LOOP_C_225;
      end
      COMP_LOOP_C_225 : begin
        fsm_output = 10'b0110111000;
        state_var_NS = COMP_LOOP_C_226;
      end
      COMP_LOOP_C_226 : begin
        fsm_output = 10'b0110111001;
        state_var_NS = COMP_LOOP_C_227;
      end
      COMP_LOOP_C_227 : begin
        fsm_output = 10'b0110111010;
        state_var_NS = COMP_LOOP_C_228;
      end
      COMP_LOOP_C_228 : begin
        fsm_output = 10'b0110111011;
        state_var_NS = COMP_LOOP_C_229;
      end
      COMP_LOOP_C_229 : begin
        fsm_output = 10'b0110111100;
        state_var_NS = COMP_LOOP_C_230;
      end
      COMP_LOOP_C_230 : begin
        fsm_output = 10'b0110111101;
        state_var_NS = COMP_LOOP_C_231;
      end
      COMP_LOOP_C_231 : begin
        fsm_output = 10'b0110111110;
        state_var_NS = COMP_LOOP_C_232;
      end
      COMP_LOOP_C_232 : begin
        fsm_output = 10'b0110111111;
        state_var_NS = COMP_LOOP_C_233;
      end
      COMP_LOOP_C_233 : begin
        fsm_output = 10'b0111000000;
        state_var_NS = COMP_LOOP_C_234;
      end
      COMP_LOOP_C_234 : begin
        fsm_output = 10'b0111000001;
        state_var_NS = COMP_LOOP_C_235;
      end
      COMP_LOOP_C_235 : begin
        fsm_output = 10'b0111000010;
        state_var_NS = COMP_LOOP_C_236;
      end
      COMP_LOOP_C_236 : begin
        fsm_output = 10'b0111000011;
        state_var_NS = COMP_LOOP_C_237;
      end
      COMP_LOOP_C_237 : begin
        fsm_output = 10'b0111000100;
        state_var_NS = COMP_LOOP_C_238;
      end
      COMP_LOOP_C_238 : begin
        fsm_output = 10'b0111000101;
        state_var_NS = COMP_LOOP_C_239;
      end
      COMP_LOOP_C_239 : begin
        fsm_output = 10'b0111000110;
        state_var_NS = COMP_LOOP_C_240;
      end
      COMP_LOOP_C_240 : begin
        fsm_output = 10'b0111000111;
        state_var_NS = COMP_LOOP_C_241;
      end
      COMP_LOOP_C_241 : begin
        fsm_output = 10'b0111001000;
        state_var_NS = COMP_LOOP_C_242;
      end
      COMP_LOOP_C_242 : begin
        fsm_output = 10'b0111001001;
        state_var_NS = COMP_LOOP_C_243;
      end
      COMP_LOOP_C_243 : begin
        fsm_output = 10'b0111001010;
        state_var_NS = COMP_LOOP_C_244;
      end
      COMP_LOOP_C_244 : begin
        fsm_output = 10'b0111001011;
        state_var_NS = COMP_LOOP_C_245;
      end
      COMP_LOOP_C_245 : begin
        fsm_output = 10'b0111001100;
        state_var_NS = COMP_LOOP_C_246;
      end
      COMP_LOOP_C_246 : begin
        fsm_output = 10'b0111001101;
        state_var_NS = COMP_LOOP_C_247;
      end
      COMP_LOOP_C_247 : begin
        fsm_output = 10'b0111001110;
        state_var_NS = COMP_LOOP_C_248;
      end
      COMP_LOOP_C_248 : begin
        fsm_output = 10'b0111001111;
        state_var_NS = COMP_LOOP_C_249;
      end
      COMP_LOOP_C_249 : begin
        fsm_output = 10'b0111010000;
        state_var_NS = COMP_LOOP_C_250;
      end
      COMP_LOOP_C_250 : begin
        fsm_output = 10'b0111010001;
        state_var_NS = COMP_LOOP_C_251;
      end
      COMP_LOOP_C_251 : begin
        fsm_output = 10'b0111010010;
        state_var_NS = COMP_LOOP_C_252;
      end
      COMP_LOOP_C_252 : begin
        fsm_output = 10'b0111010011;
        state_var_NS = COMP_LOOP_C_253;
      end
      COMP_LOOP_C_253 : begin
        fsm_output = 10'b0111010100;
        state_var_NS = COMP_LOOP_C_254;
      end
      COMP_LOOP_C_254 : begin
        fsm_output = 10'b0111010101;
        state_var_NS = COMP_LOOP_C_255;
      end
      COMP_LOOP_C_255 : begin
        fsm_output = 10'b0111010110;
        state_var_NS = COMP_LOOP_C_256;
      end
      COMP_LOOP_C_256 : begin
        fsm_output = 10'b0111010111;
        state_var_NS = COMP_LOOP_C_257;
      end
      COMP_LOOP_C_257 : begin
        fsm_output = 10'b0111011000;
        state_var_NS = COMP_LOOP_C_258;
      end
      COMP_LOOP_C_258 : begin
        fsm_output = 10'b0111011001;
        state_var_NS = COMP_LOOP_C_259;
      end
      COMP_LOOP_C_259 : begin
        fsm_output = 10'b0111011010;
        state_var_NS = COMP_LOOP_C_260;
      end
      COMP_LOOP_C_260 : begin
        fsm_output = 10'b0111011011;
        if ( COMP_LOOP_C_260_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_261;
        end
      end
      COMP_LOOP_C_261 : begin
        fsm_output = 10'b0111011100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_0;
      end
      COMP_LOOP_5_modExp_1_while_C_0 : begin
        fsm_output = 10'b0111011101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_1;
      end
      COMP_LOOP_5_modExp_1_while_C_1 : begin
        fsm_output = 10'b0111011110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_2;
      end
      COMP_LOOP_5_modExp_1_while_C_2 : begin
        fsm_output = 10'b0111011111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_3;
      end
      COMP_LOOP_5_modExp_1_while_C_3 : begin
        fsm_output = 10'b0111100000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_4;
      end
      COMP_LOOP_5_modExp_1_while_C_4 : begin
        fsm_output = 10'b0111100001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_5;
      end
      COMP_LOOP_5_modExp_1_while_C_5 : begin
        fsm_output = 10'b0111100010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_6;
      end
      COMP_LOOP_5_modExp_1_while_C_6 : begin
        fsm_output = 10'b0111100011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_7;
      end
      COMP_LOOP_5_modExp_1_while_C_7 : begin
        fsm_output = 10'b0111100100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_8;
      end
      COMP_LOOP_5_modExp_1_while_C_8 : begin
        fsm_output = 10'b0111100101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_9;
      end
      COMP_LOOP_5_modExp_1_while_C_9 : begin
        fsm_output = 10'b0111100110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_10;
      end
      COMP_LOOP_5_modExp_1_while_C_10 : begin
        fsm_output = 10'b0111100111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_11;
      end
      COMP_LOOP_5_modExp_1_while_C_11 : begin
        fsm_output = 10'b0111101000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_12;
      end
      COMP_LOOP_5_modExp_1_while_C_12 : begin
        fsm_output = 10'b0111101001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_13;
      end
      COMP_LOOP_5_modExp_1_while_C_13 : begin
        fsm_output = 10'b0111101010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_14;
      end
      COMP_LOOP_5_modExp_1_while_C_14 : begin
        fsm_output = 10'b0111101011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_15;
      end
      COMP_LOOP_5_modExp_1_while_C_15 : begin
        fsm_output = 10'b0111101100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_16;
      end
      COMP_LOOP_5_modExp_1_while_C_16 : begin
        fsm_output = 10'b0111101101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_17;
      end
      COMP_LOOP_5_modExp_1_while_C_17 : begin
        fsm_output = 10'b0111101110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_18;
      end
      COMP_LOOP_5_modExp_1_while_C_18 : begin
        fsm_output = 10'b0111101111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_19;
      end
      COMP_LOOP_5_modExp_1_while_C_19 : begin
        fsm_output = 10'b0111110000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_20;
      end
      COMP_LOOP_5_modExp_1_while_C_20 : begin
        fsm_output = 10'b0111110001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_21;
      end
      COMP_LOOP_5_modExp_1_while_C_21 : begin
        fsm_output = 10'b0111110010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_22;
      end
      COMP_LOOP_5_modExp_1_while_C_22 : begin
        fsm_output = 10'b0111110011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_23;
      end
      COMP_LOOP_5_modExp_1_while_C_23 : begin
        fsm_output = 10'b0111110100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_24;
      end
      COMP_LOOP_5_modExp_1_while_C_24 : begin
        fsm_output = 10'b0111110101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_25;
      end
      COMP_LOOP_5_modExp_1_while_C_25 : begin
        fsm_output = 10'b0111110110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_26;
      end
      COMP_LOOP_5_modExp_1_while_C_26 : begin
        fsm_output = 10'b0111110111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_27;
      end
      COMP_LOOP_5_modExp_1_while_C_27 : begin
        fsm_output = 10'b0111111000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_28;
      end
      COMP_LOOP_5_modExp_1_while_C_28 : begin
        fsm_output = 10'b0111111001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_29;
      end
      COMP_LOOP_5_modExp_1_while_C_29 : begin
        fsm_output = 10'b0111111010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_30;
      end
      COMP_LOOP_5_modExp_1_while_C_30 : begin
        fsm_output = 10'b0111111011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_31;
      end
      COMP_LOOP_5_modExp_1_while_C_31 : begin
        fsm_output = 10'b0111111100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_32;
      end
      COMP_LOOP_5_modExp_1_while_C_32 : begin
        fsm_output = 10'b0111111101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_33;
      end
      COMP_LOOP_5_modExp_1_while_C_33 : begin
        fsm_output = 10'b0111111110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_34;
      end
      COMP_LOOP_5_modExp_1_while_C_34 : begin
        fsm_output = 10'b0111111111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_35;
      end
      COMP_LOOP_5_modExp_1_while_C_35 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_36;
      end
      COMP_LOOP_5_modExp_1_while_C_36 : begin
        fsm_output = 10'b1000000001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_37;
      end
      COMP_LOOP_5_modExp_1_while_C_37 : begin
        fsm_output = 10'b1000000010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_38;
      end
      COMP_LOOP_5_modExp_1_while_C_38 : begin
        fsm_output = 10'b1000000011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_39;
      end
      COMP_LOOP_5_modExp_1_while_C_39 : begin
        fsm_output = 10'b1000000100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_40;
      end
      COMP_LOOP_5_modExp_1_while_C_40 : begin
        fsm_output = 10'b1000000101;
        if ( COMP_LOOP_5_modExp_1_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_262;
        end
        else begin
          state_var_NS = COMP_LOOP_5_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_262 : begin
        fsm_output = 10'b1000000110;
        state_var_NS = COMP_LOOP_C_263;
      end
      COMP_LOOP_C_263 : begin
        fsm_output = 10'b1000000111;
        state_var_NS = COMP_LOOP_C_264;
      end
      COMP_LOOP_C_264 : begin
        fsm_output = 10'b1000001000;
        state_var_NS = COMP_LOOP_C_265;
      end
      COMP_LOOP_C_265 : begin
        fsm_output = 10'b1000001001;
        state_var_NS = COMP_LOOP_C_266;
      end
      COMP_LOOP_C_266 : begin
        fsm_output = 10'b1000001010;
        state_var_NS = COMP_LOOP_C_267;
      end
      COMP_LOOP_C_267 : begin
        fsm_output = 10'b1000001011;
        state_var_NS = COMP_LOOP_C_268;
      end
      COMP_LOOP_C_268 : begin
        fsm_output = 10'b1000001100;
        state_var_NS = COMP_LOOP_C_269;
      end
      COMP_LOOP_C_269 : begin
        fsm_output = 10'b1000001101;
        state_var_NS = COMP_LOOP_C_270;
      end
      COMP_LOOP_C_270 : begin
        fsm_output = 10'b1000001110;
        state_var_NS = COMP_LOOP_C_271;
      end
      COMP_LOOP_C_271 : begin
        fsm_output = 10'b1000001111;
        state_var_NS = COMP_LOOP_C_272;
      end
      COMP_LOOP_C_272 : begin
        fsm_output = 10'b1000010000;
        state_var_NS = COMP_LOOP_C_273;
      end
      COMP_LOOP_C_273 : begin
        fsm_output = 10'b1000010001;
        state_var_NS = COMP_LOOP_C_274;
      end
      COMP_LOOP_C_274 : begin
        fsm_output = 10'b1000010010;
        state_var_NS = COMP_LOOP_C_275;
      end
      COMP_LOOP_C_275 : begin
        fsm_output = 10'b1000010011;
        state_var_NS = COMP_LOOP_C_276;
      end
      COMP_LOOP_C_276 : begin
        fsm_output = 10'b1000010100;
        state_var_NS = COMP_LOOP_C_277;
      end
      COMP_LOOP_C_277 : begin
        fsm_output = 10'b1000010101;
        state_var_NS = COMP_LOOP_C_278;
      end
      COMP_LOOP_C_278 : begin
        fsm_output = 10'b1000010110;
        state_var_NS = COMP_LOOP_C_279;
      end
      COMP_LOOP_C_279 : begin
        fsm_output = 10'b1000010111;
        state_var_NS = COMP_LOOP_C_280;
      end
      COMP_LOOP_C_280 : begin
        fsm_output = 10'b1000011000;
        state_var_NS = COMP_LOOP_C_281;
      end
      COMP_LOOP_C_281 : begin
        fsm_output = 10'b1000011001;
        state_var_NS = COMP_LOOP_C_282;
      end
      COMP_LOOP_C_282 : begin
        fsm_output = 10'b1000011010;
        state_var_NS = COMP_LOOP_C_283;
      end
      COMP_LOOP_C_283 : begin
        fsm_output = 10'b1000011011;
        state_var_NS = COMP_LOOP_C_284;
      end
      COMP_LOOP_C_284 : begin
        fsm_output = 10'b1000011100;
        state_var_NS = COMP_LOOP_C_285;
      end
      COMP_LOOP_C_285 : begin
        fsm_output = 10'b1000011101;
        state_var_NS = COMP_LOOP_C_286;
      end
      COMP_LOOP_C_286 : begin
        fsm_output = 10'b1000011110;
        state_var_NS = COMP_LOOP_C_287;
      end
      COMP_LOOP_C_287 : begin
        fsm_output = 10'b1000011111;
        state_var_NS = COMP_LOOP_C_288;
      end
      COMP_LOOP_C_288 : begin
        fsm_output = 10'b1000100000;
        state_var_NS = COMP_LOOP_C_289;
      end
      COMP_LOOP_C_289 : begin
        fsm_output = 10'b1000100001;
        state_var_NS = COMP_LOOP_C_290;
      end
      COMP_LOOP_C_290 : begin
        fsm_output = 10'b1000100010;
        state_var_NS = COMP_LOOP_C_291;
      end
      COMP_LOOP_C_291 : begin
        fsm_output = 10'b1000100011;
        state_var_NS = COMP_LOOP_C_292;
      end
      COMP_LOOP_C_292 : begin
        fsm_output = 10'b1000100100;
        state_var_NS = COMP_LOOP_C_293;
      end
      COMP_LOOP_C_293 : begin
        fsm_output = 10'b1000100101;
        state_var_NS = COMP_LOOP_C_294;
      end
      COMP_LOOP_C_294 : begin
        fsm_output = 10'b1000100110;
        state_var_NS = COMP_LOOP_C_295;
      end
      COMP_LOOP_C_295 : begin
        fsm_output = 10'b1000100111;
        state_var_NS = COMP_LOOP_C_296;
      end
      COMP_LOOP_C_296 : begin
        fsm_output = 10'b1000101000;
        state_var_NS = COMP_LOOP_C_297;
      end
      COMP_LOOP_C_297 : begin
        fsm_output = 10'b1000101001;
        state_var_NS = COMP_LOOP_C_298;
      end
      COMP_LOOP_C_298 : begin
        fsm_output = 10'b1000101010;
        state_var_NS = COMP_LOOP_C_299;
      end
      COMP_LOOP_C_299 : begin
        fsm_output = 10'b1000101011;
        state_var_NS = COMP_LOOP_C_300;
      end
      COMP_LOOP_C_300 : begin
        fsm_output = 10'b1000101100;
        state_var_NS = COMP_LOOP_C_301;
      end
      COMP_LOOP_C_301 : begin
        fsm_output = 10'b1000101101;
        state_var_NS = COMP_LOOP_C_302;
      end
      COMP_LOOP_C_302 : begin
        fsm_output = 10'b1000101110;
        state_var_NS = COMP_LOOP_C_303;
      end
      COMP_LOOP_C_303 : begin
        fsm_output = 10'b1000101111;
        state_var_NS = COMP_LOOP_C_304;
      end
      COMP_LOOP_C_304 : begin
        fsm_output = 10'b1000110000;
        state_var_NS = COMP_LOOP_C_305;
      end
      COMP_LOOP_C_305 : begin
        fsm_output = 10'b1000110001;
        state_var_NS = COMP_LOOP_C_306;
      end
      COMP_LOOP_C_306 : begin
        fsm_output = 10'b1000110010;
        state_var_NS = COMP_LOOP_C_307;
      end
      COMP_LOOP_C_307 : begin
        fsm_output = 10'b1000110011;
        state_var_NS = COMP_LOOP_C_308;
      end
      COMP_LOOP_C_308 : begin
        fsm_output = 10'b1000110100;
        state_var_NS = COMP_LOOP_C_309;
      end
      COMP_LOOP_C_309 : begin
        fsm_output = 10'b1000110101;
        state_var_NS = COMP_LOOP_C_310;
      end
      COMP_LOOP_C_310 : begin
        fsm_output = 10'b1000110110;
        state_var_NS = COMP_LOOP_C_311;
      end
      COMP_LOOP_C_311 : begin
        fsm_output = 10'b1000110111;
        state_var_NS = COMP_LOOP_C_312;
      end
      COMP_LOOP_C_312 : begin
        fsm_output = 10'b1000111000;
        state_var_NS = COMP_LOOP_C_313;
      end
      COMP_LOOP_C_313 : begin
        fsm_output = 10'b1000111001;
        state_var_NS = COMP_LOOP_C_314;
      end
      COMP_LOOP_C_314 : begin
        fsm_output = 10'b1000111010;
        state_var_NS = COMP_LOOP_C_315;
      end
      COMP_LOOP_C_315 : begin
        fsm_output = 10'b1000111011;
        state_var_NS = COMP_LOOP_C_316;
      end
      COMP_LOOP_C_316 : begin
        fsm_output = 10'b1000111100;
        state_var_NS = COMP_LOOP_C_317;
      end
      COMP_LOOP_C_317 : begin
        fsm_output = 10'b1000111101;
        state_var_NS = COMP_LOOP_C_318;
      end
      COMP_LOOP_C_318 : begin
        fsm_output = 10'b1000111110;
        state_var_NS = COMP_LOOP_C_319;
      end
      COMP_LOOP_C_319 : begin
        fsm_output = 10'b1000111111;
        state_var_NS = COMP_LOOP_C_320;
      end
      COMP_LOOP_C_320 : begin
        fsm_output = 10'b1001000000;
        state_var_NS = COMP_LOOP_C_321;
      end
      COMP_LOOP_C_321 : begin
        fsm_output = 10'b1001000001;
        state_var_NS = COMP_LOOP_C_322;
      end
      COMP_LOOP_C_322 : begin
        fsm_output = 10'b1001000010;
        state_var_NS = COMP_LOOP_C_323;
      end
      COMP_LOOP_C_323 : begin
        fsm_output = 10'b1001000011;
        state_var_NS = COMP_LOOP_C_324;
      end
      COMP_LOOP_C_324 : begin
        fsm_output = 10'b1001000100;
        state_var_NS = COMP_LOOP_C_325;
      end
      COMP_LOOP_C_325 : begin
        fsm_output = 10'b1001000101;
        if ( COMP_LOOP_C_325_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_326;
        end
      end
      COMP_LOOP_C_326 : begin
        fsm_output = 10'b1001000110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_0;
      end
      COMP_LOOP_6_modExp_1_while_C_0 : begin
        fsm_output = 10'b1001000111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_1;
      end
      COMP_LOOP_6_modExp_1_while_C_1 : begin
        fsm_output = 10'b1001001000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_2;
      end
      COMP_LOOP_6_modExp_1_while_C_2 : begin
        fsm_output = 10'b1001001001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_3;
      end
      COMP_LOOP_6_modExp_1_while_C_3 : begin
        fsm_output = 10'b1001001010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_4;
      end
      COMP_LOOP_6_modExp_1_while_C_4 : begin
        fsm_output = 10'b1001001011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_5;
      end
      COMP_LOOP_6_modExp_1_while_C_5 : begin
        fsm_output = 10'b1001001100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_6;
      end
      COMP_LOOP_6_modExp_1_while_C_6 : begin
        fsm_output = 10'b1001001101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_7;
      end
      COMP_LOOP_6_modExp_1_while_C_7 : begin
        fsm_output = 10'b1001001110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_8;
      end
      COMP_LOOP_6_modExp_1_while_C_8 : begin
        fsm_output = 10'b1001001111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_9;
      end
      COMP_LOOP_6_modExp_1_while_C_9 : begin
        fsm_output = 10'b1001010000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_10;
      end
      COMP_LOOP_6_modExp_1_while_C_10 : begin
        fsm_output = 10'b1001010001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_11;
      end
      COMP_LOOP_6_modExp_1_while_C_11 : begin
        fsm_output = 10'b1001010010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_12;
      end
      COMP_LOOP_6_modExp_1_while_C_12 : begin
        fsm_output = 10'b1001010011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_13;
      end
      COMP_LOOP_6_modExp_1_while_C_13 : begin
        fsm_output = 10'b1001010100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_14;
      end
      COMP_LOOP_6_modExp_1_while_C_14 : begin
        fsm_output = 10'b1001010101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_15;
      end
      COMP_LOOP_6_modExp_1_while_C_15 : begin
        fsm_output = 10'b1001010110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_16;
      end
      COMP_LOOP_6_modExp_1_while_C_16 : begin
        fsm_output = 10'b1001010111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_17;
      end
      COMP_LOOP_6_modExp_1_while_C_17 : begin
        fsm_output = 10'b1001011000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_18;
      end
      COMP_LOOP_6_modExp_1_while_C_18 : begin
        fsm_output = 10'b1001011001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_19;
      end
      COMP_LOOP_6_modExp_1_while_C_19 : begin
        fsm_output = 10'b1001011010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_20;
      end
      COMP_LOOP_6_modExp_1_while_C_20 : begin
        fsm_output = 10'b1001011011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_21;
      end
      COMP_LOOP_6_modExp_1_while_C_21 : begin
        fsm_output = 10'b1001011100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_22;
      end
      COMP_LOOP_6_modExp_1_while_C_22 : begin
        fsm_output = 10'b1001011101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_23;
      end
      COMP_LOOP_6_modExp_1_while_C_23 : begin
        fsm_output = 10'b1001011110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_24;
      end
      COMP_LOOP_6_modExp_1_while_C_24 : begin
        fsm_output = 10'b1001011111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_25;
      end
      COMP_LOOP_6_modExp_1_while_C_25 : begin
        fsm_output = 10'b1001100000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_26;
      end
      COMP_LOOP_6_modExp_1_while_C_26 : begin
        fsm_output = 10'b1001100001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_27;
      end
      COMP_LOOP_6_modExp_1_while_C_27 : begin
        fsm_output = 10'b1001100010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_28;
      end
      COMP_LOOP_6_modExp_1_while_C_28 : begin
        fsm_output = 10'b1001100011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_29;
      end
      COMP_LOOP_6_modExp_1_while_C_29 : begin
        fsm_output = 10'b1001100100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_30;
      end
      COMP_LOOP_6_modExp_1_while_C_30 : begin
        fsm_output = 10'b1001100101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_31;
      end
      COMP_LOOP_6_modExp_1_while_C_31 : begin
        fsm_output = 10'b1001100110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_32;
      end
      COMP_LOOP_6_modExp_1_while_C_32 : begin
        fsm_output = 10'b1001100111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_33;
      end
      COMP_LOOP_6_modExp_1_while_C_33 : begin
        fsm_output = 10'b1001101000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_34;
      end
      COMP_LOOP_6_modExp_1_while_C_34 : begin
        fsm_output = 10'b1001101001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_35;
      end
      COMP_LOOP_6_modExp_1_while_C_35 : begin
        fsm_output = 10'b1001101010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_36;
      end
      COMP_LOOP_6_modExp_1_while_C_36 : begin
        fsm_output = 10'b1001101011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_37;
      end
      COMP_LOOP_6_modExp_1_while_C_37 : begin
        fsm_output = 10'b1001101100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_38;
      end
      COMP_LOOP_6_modExp_1_while_C_38 : begin
        fsm_output = 10'b1001101101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_39;
      end
      COMP_LOOP_6_modExp_1_while_C_39 : begin
        fsm_output = 10'b1001101110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_40;
      end
      COMP_LOOP_6_modExp_1_while_C_40 : begin
        fsm_output = 10'b1001101111;
        if ( COMP_LOOP_6_modExp_1_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_327;
        end
        else begin
          state_var_NS = COMP_LOOP_6_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_327 : begin
        fsm_output = 10'b1001110000;
        state_var_NS = COMP_LOOP_C_328;
      end
      COMP_LOOP_C_328 : begin
        fsm_output = 10'b1001110001;
        state_var_NS = COMP_LOOP_C_329;
      end
      COMP_LOOP_C_329 : begin
        fsm_output = 10'b1001110010;
        state_var_NS = COMP_LOOP_C_330;
      end
      COMP_LOOP_C_330 : begin
        fsm_output = 10'b1001110011;
        state_var_NS = COMP_LOOP_C_331;
      end
      COMP_LOOP_C_331 : begin
        fsm_output = 10'b1001110100;
        state_var_NS = COMP_LOOP_C_332;
      end
      COMP_LOOP_C_332 : begin
        fsm_output = 10'b1001110101;
        state_var_NS = COMP_LOOP_C_333;
      end
      COMP_LOOP_C_333 : begin
        fsm_output = 10'b1001110110;
        state_var_NS = COMP_LOOP_C_334;
      end
      COMP_LOOP_C_334 : begin
        fsm_output = 10'b1001110111;
        state_var_NS = COMP_LOOP_C_335;
      end
      COMP_LOOP_C_335 : begin
        fsm_output = 10'b1001111000;
        state_var_NS = COMP_LOOP_C_336;
      end
      COMP_LOOP_C_336 : begin
        fsm_output = 10'b1001111001;
        state_var_NS = COMP_LOOP_C_337;
      end
      COMP_LOOP_C_337 : begin
        fsm_output = 10'b1001111010;
        state_var_NS = COMP_LOOP_C_338;
      end
      COMP_LOOP_C_338 : begin
        fsm_output = 10'b1001111011;
        state_var_NS = COMP_LOOP_C_339;
      end
      COMP_LOOP_C_339 : begin
        fsm_output = 10'b1001111100;
        state_var_NS = COMP_LOOP_C_340;
      end
      COMP_LOOP_C_340 : begin
        fsm_output = 10'b1001111101;
        state_var_NS = COMP_LOOP_C_341;
      end
      COMP_LOOP_C_341 : begin
        fsm_output = 10'b1001111110;
        state_var_NS = COMP_LOOP_C_342;
      end
      COMP_LOOP_C_342 : begin
        fsm_output = 10'b1001111111;
        state_var_NS = COMP_LOOP_C_343;
      end
      COMP_LOOP_C_343 : begin
        fsm_output = 10'b1010000000;
        state_var_NS = COMP_LOOP_C_344;
      end
      COMP_LOOP_C_344 : begin
        fsm_output = 10'b1010000001;
        state_var_NS = COMP_LOOP_C_345;
      end
      COMP_LOOP_C_345 : begin
        fsm_output = 10'b1010000010;
        state_var_NS = COMP_LOOP_C_346;
      end
      COMP_LOOP_C_346 : begin
        fsm_output = 10'b1010000011;
        state_var_NS = COMP_LOOP_C_347;
      end
      COMP_LOOP_C_347 : begin
        fsm_output = 10'b1010000100;
        state_var_NS = COMP_LOOP_C_348;
      end
      COMP_LOOP_C_348 : begin
        fsm_output = 10'b1010000101;
        state_var_NS = COMP_LOOP_C_349;
      end
      COMP_LOOP_C_349 : begin
        fsm_output = 10'b1010000110;
        state_var_NS = COMP_LOOP_C_350;
      end
      COMP_LOOP_C_350 : begin
        fsm_output = 10'b1010000111;
        state_var_NS = COMP_LOOP_C_351;
      end
      COMP_LOOP_C_351 : begin
        fsm_output = 10'b1010001000;
        state_var_NS = COMP_LOOP_C_352;
      end
      COMP_LOOP_C_352 : begin
        fsm_output = 10'b1010001001;
        state_var_NS = COMP_LOOP_C_353;
      end
      COMP_LOOP_C_353 : begin
        fsm_output = 10'b1010001010;
        state_var_NS = COMP_LOOP_C_354;
      end
      COMP_LOOP_C_354 : begin
        fsm_output = 10'b1010001011;
        state_var_NS = COMP_LOOP_C_355;
      end
      COMP_LOOP_C_355 : begin
        fsm_output = 10'b1010001100;
        state_var_NS = COMP_LOOP_C_356;
      end
      COMP_LOOP_C_356 : begin
        fsm_output = 10'b1010001101;
        state_var_NS = COMP_LOOP_C_357;
      end
      COMP_LOOP_C_357 : begin
        fsm_output = 10'b1010001110;
        state_var_NS = COMP_LOOP_C_358;
      end
      COMP_LOOP_C_358 : begin
        fsm_output = 10'b1010001111;
        state_var_NS = COMP_LOOP_C_359;
      end
      COMP_LOOP_C_359 : begin
        fsm_output = 10'b1010010000;
        state_var_NS = COMP_LOOP_C_360;
      end
      COMP_LOOP_C_360 : begin
        fsm_output = 10'b1010010001;
        state_var_NS = COMP_LOOP_C_361;
      end
      COMP_LOOP_C_361 : begin
        fsm_output = 10'b1010010010;
        state_var_NS = COMP_LOOP_C_362;
      end
      COMP_LOOP_C_362 : begin
        fsm_output = 10'b1010010011;
        state_var_NS = COMP_LOOP_C_363;
      end
      COMP_LOOP_C_363 : begin
        fsm_output = 10'b1010010100;
        state_var_NS = COMP_LOOP_C_364;
      end
      COMP_LOOP_C_364 : begin
        fsm_output = 10'b1010010101;
        state_var_NS = COMP_LOOP_C_365;
      end
      COMP_LOOP_C_365 : begin
        fsm_output = 10'b1010010110;
        state_var_NS = COMP_LOOP_C_366;
      end
      COMP_LOOP_C_366 : begin
        fsm_output = 10'b1010010111;
        state_var_NS = COMP_LOOP_C_367;
      end
      COMP_LOOP_C_367 : begin
        fsm_output = 10'b1010011000;
        state_var_NS = COMP_LOOP_C_368;
      end
      COMP_LOOP_C_368 : begin
        fsm_output = 10'b1010011001;
        state_var_NS = COMP_LOOP_C_369;
      end
      COMP_LOOP_C_369 : begin
        fsm_output = 10'b1010011010;
        state_var_NS = COMP_LOOP_C_370;
      end
      COMP_LOOP_C_370 : begin
        fsm_output = 10'b1010011011;
        state_var_NS = COMP_LOOP_C_371;
      end
      COMP_LOOP_C_371 : begin
        fsm_output = 10'b1010011100;
        state_var_NS = COMP_LOOP_C_372;
      end
      COMP_LOOP_C_372 : begin
        fsm_output = 10'b1010011101;
        state_var_NS = COMP_LOOP_C_373;
      end
      COMP_LOOP_C_373 : begin
        fsm_output = 10'b1010011110;
        state_var_NS = COMP_LOOP_C_374;
      end
      COMP_LOOP_C_374 : begin
        fsm_output = 10'b1010011111;
        state_var_NS = COMP_LOOP_C_375;
      end
      COMP_LOOP_C_375 : begin
        fsm_output = 10'b1010100000;
        state_var_NS = COMP_LOOP_C_376;
      end
      COMP_LOOP_C_376 : begin
        fsm_output = 10'b1010100001;
        state_var_NS = COMP_LOOP_C_377;
      end
      COMP_LOOP_C_377 : begin
        fsm_output = 10'b1010100010;
        state_var_NS = COMP_LOOP_C_378;
      end
      COMP_LOOP_C_378 : begin
        fsm_output = 10'b1010100011;
        state_var_NS = COMP_LOOP_C_379;
      end
      COMP_LOOP_C_379 : begin
        fsm_output = 10'b1010100100;
        state_var_NS = COMP_LOOP_C_380;
      end
      COMP_LOOP_C_380 : begin
        fsm_output = 10'b1010100101;
        state_var_NS = COMP_LOOP_C_381;
      end
      COMP_LOOP_C_381 : begin
        fsm_output = 10'b1010100110;
        state_var_NS = COMP_LOOP_C_382;
      end
      COMP_LOOP_C_382 : begin
        fsm_output = 10'b1010100111;
        state_var_NS = COMP_LOOP_C_383;
      end
      COMP_LOOP_C_383 : begin
        fsm_output = 10'b1010101000;
        state_var_NS = COMP_LOOP_C_384;
      end
      COMP_LOOP_C_384 : begin
        fsm_output = 10'b1010101001;
        state_var_NS = COMP_LOOP_C_385;
      end
      COMP_LOOP_C_385 : begin
        fsm_output = 10'b1010101010;
        state_var_NS = COMP_LOOP_C_386;
      end
      COMP_LOOP_C_386 : begin
        fsm_output = 10'b1010101011;
        state_var_NS = COMP_LOOP_C_387;
      end
      COMP_LOOP_C_387 : begin
        fsm_output = 10'b1010101100;
        state_var_NS = COMP_LOOP_C_388;
      end
      COMP_LOOP_C_388 : begin
        fsm_output = 10'b1010101101;
        state_var_NS = COMP_LOOP_C_389;
      end
      COMP_LOOP_C_389 : begin
        fsm_output = 10'b1010101110;
        state_var_NS = COMP_LOOP_C_390;
      end
      COMP_LOOP_C_390 : begin
        fsm_output = 10'b1010101111;
        if ( COMP_LOOP_C_390_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_391;
        end
      end
      COMP_LOOP_C_391 : begin
        fsm_output = 10'b1010110000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_0;
      end
      COMP_LOOP_7_modExp_1_while_C_0 : begin
        fsm_output = 10'b1010110001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_1;
      end
      COMP_LOOP_7_modExp_1_while_C_1 : begin
        fsm_output = 10'b1010110010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_2;
      end
      COMP_LOOP_7_modExp_1_while_C_2 : begin
        fsm_output = 10'b1010110011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_3;
      end
      COMP_LOOP_7_modExp_1_while_C_3 : begin
        fsm_output = 10'b1010110100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_4;
      end
      COMP_LOOP_7_modExp_1_while_C_4 : begin
        fsm_output = 10'b1010110101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_5;
      end
      COMP_LOOP_7_modExp_1_while_C_5 : begin
        fsm_output = 10'b1010110110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_6;
      end
      COMP_LOOP_7_modExp_1_while_C_6 : begin
        fsm_output = 10'b1010110111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_7;
      end
      COMP_LOOP_7_modExp_1_while_C_7 : begin
        fsm_output = 10'b1010111000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_8;
      end
      COMP_LOOP_7_modExp_1_while_C_8 : begin
        fsm_output = 10'b1010111001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_9;
      end
      COMP_LOOP_7_modExp_1_while_C_9 : begin
        fsm_output = 10'b1010111010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_10;
      end
      COMP_LOOP_7_modExp_1_while_C_10 : begin
        fsm_output = 10'b1010111011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_11;
      end
      COMP_LOOP_7_modExp_1_while_C_11 : begin
        fsm_output = 10'b1010111100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_12;
      end
      COMP_LOOP_7_modExp_1_while_C_12 : begin
        fsm_output = 10'b1010111101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_13;
      end
      COMP_LOOP_7_modExp_1_while_C_13 : begin
        fsm_output = 10'b1010111110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_14;
      end
      COMP_LOOP_7_modExp_1_while_C_14 : begin
        fsm_output = 10'b1010111111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_15;
      end
      COMP_LOOP_7_modExp_1_while_C_15 : begin
        fsm_output = 10'b1011000000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_16;
      end
      COMP_LOOP_7_modExp_1_while_C_16 : begin
        fsm_output = 10'b1011000001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_17;
      end
      COMP_LOOP_7_modExp_1_while_C_17 : begin
        fsm_output = 10'b1011000010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_18;
      end
      COMP_LOOP_7_modExp_1_while_C_18 : begin
        fsm_output = 10'b1011000011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_19;
      end
      COMP_LOOP_7_modExp_1_while_C_19 : begin
        fsm_output = 10'b1011000100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_20;
      end
      COMP_LOOP_7_modExp_1_while_C_20 : begin
        fsm_output = 10'b1011000101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_21;
      end
      COMP_LOOP_7_modExp_1_while_C_21 : begin
        fsm_output = 10'b1011000110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_22;
      end
      COMP_LOOP_7_modExp_1_while_C_22 : begin
        fsm_output = 10'b1011000111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_23;
      end
      COMP_LOOP_7_modExp_1_while_C_23 : begin
        fsm_output = 10'b1011001000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_24;
      end
      COMP_LOOP_7_modExp_1_while_C_24 : begin
        fsm_output = 10'b1011001001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_25;
      end
      COMP_LOOP_7_modExp_1_while_C_25 : begin
        fsm_output = 10'b1011001010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_26;
      end
      COMP_LOOP_7_modExp_1_while_C_26 : begin
        fsm_output = 10'b1011001011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_27;
      end
      COMP_LOOP_7_modExp_1_while_C_27 : begin
        fsm_output = 10'b1011001100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_28;
      end
      COMP_LOOP_7_modExp_1_while_C_28 : begin
        fsm_output = 10'b1011001101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_29;
      end
      COMP_LOOP_7_modExp_1_while_C_29 : begin
        fsm_output = 10'b1011001110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_30;
      end
      COMP_LOOP_7_modExp_1_while_C_30 : begin
        fsm_output = 10'b1011001111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_31;
      end
      COMP_LOOP_7_modExp_1_while_C_31 : begin
        fsm_output = 10'b1011010000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_32;
      end
      COMP_LOOP_7_modExp_1_while_C_32 : begin
        fsm_output = 10'b1011010001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_33;
      end
      COMP_LOOP_7_modExp_1_while_C_33 : begin
        fsm_output = 10'b1011010010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_34;
      end
      COMP_LOOP_7_modExp_1_while_C_34 : begin
        fsm_output = 10'b1011010011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_35;
      end
      COMP_LOOP_7_modExp_1_while_C_35 : begin
        fsm_output = 10'b1011010100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_36;
      end
      COMP_LOOP_7_modExp_1_while_C_36 : begin
        fsm_output = 10'b1011010101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_37;
      end
      COMP_LOOP_7_modExp_1_while_C_37 : begin
        fsm_output = 10'b1011010110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_38;
      end
      COMP_LOOP_7_modExp_1_while_C_38 : begin
        fsm_output = 10'b1011010111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_39;
      end
      COMP_LOOP_7_modExp_1_while_C_39 : begin
        fsm_output = 10'b1011011000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_40;
      end
      COMP_LOOP_7_modExp_1_while_C_40 : begin
        fsm_output = 10'b1011011001;
        if ( COMP_LOOP_7_modExp_1_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_392;
        end
        else begin
          state_var_NS = COMP_LOOP_7_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_392 : begin
        fsm_output = 10'b1011011010;
        state_var_NS = COMP_LOOP_C_393;
      end
      COMP_LOOP_C_393 : begin
        fsm_output = 10'b1011011011;
        state_var_NS = COMP_LOOP_C_394;
      end
      COMP_LOOP_C_394 : begin
        fsm_output = 10'b1011011100;
        state_var_NS = COMP_LOOP_C_395;
      end
      COMP_LOOP_C_395 : begin
        fsm_output = 10'b1011011101;
        state_var_NS = COMP_LOOP_C_396;
      end
      COMP_LOOP_C_396 : begin
        fsm_output = 10'b1011011110;
        state_var_NS = COMP_LOOP_C_397;
      end
      COMP_LOOP_C_397 : begin
        fsm_output = 10'b1011011111;
        state_var_NS = COMP_LOOP_C_398;
      end
      COMP_LOOP_C_398 : begin
        fsm_output = 10'b1011100000;
        state_var_NS = COMP_LOOP_C_399;
      end
      COMP_LOOP_C_399 : begin
        fsm_output = 10'b1011100001;
        state_var_NS = COMP_LOOP_C_400;
      end
      COMP_LOOP_C_400 : begin
        fsm_output = 10'b1011100010;
        state_var_NS = COMP_LOOP_C_401;
      end
      COMP_LOOP_C_401 : begin
        fsm_output = 10'b1011100011;
        state_var_NS = COMP_LOOP_C_402;
      end
      COMP_LOOP_C_402 : begin
        fsm_output = 10'b1011100100;
        state_var_NS = COMP_LOOP_C_403;
      end
      COMP_LOOP_C_403 : begin
        fsm_output = 10'b1011100101;
        state_var_NS = COMP_LOOP_C_404;
      end
      COMP_LOOP_C_404 : begin
        fsm_output = 10'b1011100110;
        state_var_NS = COMP_LOOP_C_405;
      end
      COMP_LOOP_C_405 : begin
        fsm_output = 10'b1011100111;
        state_var_NS = COMP_LOOP_C_406;
      end
      COMP_LOOP_C_406 : begin
        fsm_output = 10'b1011101000;
        state_var_NS = COMP_LOOP_C_407;
      end
      COMP_LOOP_C_407 : begin
        fsm_output = 10'b1011101001;
        state_var_NS = COMP_LOOP_C_408;
      end
      COMP_LOOP_C_408 : begin
        fsm_output = 10'b1011101010;
        state_var_NS = COMP_LOOP_C_409;
      end
      COMP_LOOP_C_409 : begin
        fsm_output = 10'b1011101011;
        state_var_NS = COMP_LOOP_C_410;
      end
      COMP_LOOP_C_410 : begin
        fsm_output = 10'b1011101100;
        state_var_NS = COMP_LOOP_C_411;
      end
      COMP_LOOP_C_411 : begin
        fsm_output = 10'b1011101101;
        state_var_NS = COMP_LOOP_C_412;
      end
      COMP_LOOP_C_412 : begin
        fsm_output = 10'b1011101110;
        state_var_NS = COMP_LOOP_C_413;
      end
      COMP_LOOP_C_413 : begin
        fsm_output = 10'b1011101111;
        state_var_NS = COMP_LOOP_C_414;
      end
      COMP_LOOP_C_414 : begin
        fsm_output = 10'b1011110000;
        state_var_NS = COMP_LOOP_C_415;
      end
      COMP_LOOP_C_415 : begin
        fsm_output = 10'b1011110001;
        state_var_NS = COMP_LOOP_C_416;
      end
      COMP_LOOP_C_416 : begin
        fsm_output = 10'b1011110010;
        state_var_NS = COMP_LOOP_C_417;
      end
      COMP_LOOP_C_417 : begin
        fsm_output = 10'b1011110011;
        state_var_NS = COMP_LOOP_C_418;
      end
      COMP_LOOP_C_418 : begin
        fsm_output = 10'b1011110100;
        state_var_NS = COMP_LOOP_C_419;
      end
      COMP_LOOP_C_419 : begin
        fsm_output = 10'b1011110101;
        state_var_NS = COMP_LOOP_C_420;
      end
      COMP_LOOP_C_420 : begin
        fsm_output = 10'b1011110110;
        state_var_NS = COMP_LOOP_C_421;
      end
      COMP_LOOP_C_421 : begin
        fsm_output = 10'b1011110111;
        state_var_NS = COMP_LOOP_C_422;
      end
      COMP_LOOP_C_422 : begin
        fsm_output = 10'b1011111000;
        state_var_NS = COMP_LOOP_C_423;
      end
      COMP_LOOP_C_423 : begin
        fsm_output = 10'b1011111001;
        state_var_NS = COMP_LOOP_C_424;
      end
      COMP_LOOP_C_424 : begin
        fsm_output = 10'b1011111010;
        state_var_NS = COMP_LOOP_C_425;
      end
      COMP_LOOP_C_425 : begin
        fsm_output = 10'b1011111011;
        state_var_NS = COMP_LOOP_C_426;
      end
      COMP_LOOP_C_426 : begin
        fsm_output = 10'b1011111100;
        state_var_NS = COMP_LOOP_C_427;
      end
      COMP_LOOP_C_427 : begin
        fsm_output = 10'b1011111101;
        state_var_NS = COMP_LOOP_C_428;
      end
      COMP_LOOP_C_428 : begin
        fsm_output = 10'b1011111110;
        state_var_NS = COMP_LOOP_C_429;
      end
      COMP_LOOP_C_429 : begin
        fsm_output = 10'b1011111111;
        state_var_NS = COMP_LOOP_C_430;
      end
      COMP_LOOP_C_430 : begin
        fsm_output = 10'b1100000000;
        state_var_NS = COMP_LOOP_C_431;
      end
      COMP_LOOP_C_431 : begin
        fsm_output = 10'b1100000001;
        state_var_NS = COMP_LOOP_C_432;
      end
      COMP_LOOP_C_432 : begin
        fsm_output = 10'b1100000010;
        state_var_NS = COMP_LOOP_C_433;
      end
      COMP_LOOP_C_433 : begin
        fsm_output = 10'b1100000011;
        state_var_NS = COMP_LOOP_C_434;
      end
      COMP_LOOP_C_434 : begin
        fsm_output = 10'b1100000100;
        state_var_NS = COMP_LOOP_C_435;
      end
      COMP_LOOP_C_435 : begin
        fsm_output = 10'b1100000101;
        state_var_NS = COMP_LOOP_C_436;
      end
      COMP_LOOP_C_436 : begin
        fsm_output = 10'b1100000110;
        state_var_NS = COMP_LOOP_C_437;
      end
      COMP_LOOP_C_437 : begin
        fsm_output = 10'b1100000111;
        state_var_NS = COMP_LOOP_C_438;
      end
      COMP_LOOP_C_438 : begin
        fsm_output = 10'b1100001000;
        state_var_NS = COMP_LOOP_C_439;
      end
      COMP_LOOP_C_439 : begin
        fsm_output = 10'b1100001001;
        state_var_NS = COMP_LOOP_C_440;
      end
      COMP_LOOP_C_440 : begin
        fsm_output = 10'b1100001010;
        state_var_NS = COMP_LOOP_C_441;
      end
      COMP_LOOP_C_441 : begin
        fsm_output = 10'b1100001011;
        state_var_NS = COMP_LOOP_C_442;
      end
      COMP_LOOP_C_442 : begin
        fsm_output = 10'b1100001100;
        state_var_NS = COMP_LOOP_C_443;
      end
      COMP_LOOP_C_443 : begin
        fsm_output = 10'b1100001101;
        state_var_NS = COMP_LOOP_C_444;
      end
      COMP_LOOP_C_444 : begin
        fsm_output = 10'b1100001110;
        state_var_NS = COMP_LOOP_C_445;
      end
      COMP_LOOP_C_445 : begin
        fsm_output = 10'b1100001111;
        state_var_NS = COMP_LOOP_C_446;
      end
      COMP_LOOP_C_446 : begin
        fsm_output = 10'b1100010000;
        state_var_NS = COMP_LOOP_C_447;
      end
      COMP_LOOP_C_447 : begin
        fsm_output = 10'b1100010001;
        state_var_NS = COMP_LOOP_C_448;
      end
      COMP_LOOP_C_448 : begin
        fsm_output = 10'b1100010010;
        state_var_NS = COMP_LOOP_C_449;
      end
      COMP_LOOP_C_449 : begin
        fsm_output = 10'b1100010011;
        state_var_NS = COMP_LOOP_C_450;
      end
      COMP_LOOP_C_450 : begin
        fsm_output = 10'b1100010100;
        state_var_NS = COMP_LOOP_C_451;
      end
      COMP_LOOP_C_451 : begin
        fsm_output = 10'b1100010101;
        state_var_NS = COMP_LOOP_C_452;
      end
      COMP_LOOP_C_452 : begin
        fsm_output = 10'b1100010110;
        state_var_NS = COMP_LOOP_C_453;
      end
      COMP_LOOP_C_453 : begin
        fsm_output = 10'b1100010111;
        state_var_NS = COMP_LOOP_C_454;
      end
      COMP_LOOP_C_454 : begin
        fsm_output = 10'b1100011000;
        state_var_NS = COMP_LOOP_C_455;
      end
      COMP_LOOP_C_455 : begin
        fsm_output = 10'b1100011001;
        if ( COMP_LOOP_C_455_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_456;
        end
      end
      COMP_LOOP_C_456 : begin
        fsm_output = 10'b1100011010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_0;
      end
      COMP_LOOP_8_modExp_1_while_C_0 : begin
        fsm_output = 10'b1100011011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_1;
      end
      COMP_LOOP_8_modExp_1_while_C_1 : begin
        fsm_output = 10'b1100011100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_2;
      end
      COMP_LOOP_8_modExp_1_while_C_2 : begin
        fsm_output = 10'b1100011101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_3;
      end
      COMP_LOOP_8_modExp_1_while_C_3 : begin
        fsm_output = 10'b1100011110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_4;
      end
      COMP_LOOP_8_modExp_1_while_C_4 : begin
        fsm_output = 10'b1100011111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_5;
      end
      COMP_LOOP_8_modExp_1_while_C_5 : begin
        fsm_output = 10'b1100100000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_6;
      end
      COMP_LOOP_8_modExp_1_while_C_6 : begin
        fsm_output = 10'b1100100001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_7;
      end
      COMP_LOOP_8_modExp_1_while_C_7 : begin
        fsm_output = 10'b1100100010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_8;
      end
      COMP_LOOP_8_modExp_1_while_C_8 : begin
        fsm_output = 10'b1100100011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_9;
      end
      COMP_LOOP_8_modExp_1_while_C_9 : begin
        fsm_output = 10'b1100100100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_10;
      end
      COMP_LOOP_8_modExp_1_while_C_10 : begin
        fsm_output = 10'b1100100101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_11;
      end
      COMP_LOOP_8_modExp_1_while_C_11 : begin
        fsm_output = 10'b1100100110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_12;
      end
      COMP_LOOP_8_modExp_1_while_C_12 : begin
        fsm_output = 10'b1100100111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_13;
      end
      COMP_LOOP_8_modExp_1_while_C_13 : begin
        fsm_output = 10'b1100101000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_14;
      end
      COMP_LOOP_8_modExp_1_while_C_14 : begin
        fsm_output = 10'b1100101001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_15;
      end
      COMP_LOOP_8_modExp_1_while_C_15 : begin
        fsm_output = 10'b1100101010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_16;
      end
      COMP_LOOP_8_modExp_1_while_C_16 : begin
        fsm_output = 10'b1100101011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_17;
      end
      COMP_LOOP_8_modExp_1_while_C_17 : begin
        fsm_output = 10'b1100101100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_18;
      end
      COMP_LOOP_8_modExp_1_while_C_18 : begin
        fsm_output = 10'b1100101101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_19;
      end
      COMP_LOOP_8_modExp_1_while_C_19 : begin
        fsm_output = 10'b1100101110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_20;
      end
      COMP_LOOP_8_modExp_1_while_C_20 : begin
        fsm_output = 10'b1100101111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_21;
      end
      COMP_LOOP_8_modExp_1_while_C_21 : begin
        fsm_output = 10'b1100110000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_22;
      end
      COMP_LOOP_8_modExp_1_while_C_22 : begin
        fsm_output = 10'b1100110001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_23;
      end
      COMP_LOOP_8_modExp_1_while_C_23 : begin
        fsm_output = 10'b1100110010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_24;
      end
      COMP_LOOP_8_modExp_1_while_C_24 : begin
        fsm_output = 10'b1100110011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_25;
      end
      COMP_LOOP_8_modExp_1_while_C_25 : begin
        fsm_output = 10'b1100110100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_26;
      end
      COMP_LOOP_8_modExp_1_while_C_26 : begin
        fsm_output = 10'b1100110101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_27;
      end
      COMP_LOOP_8_modExp_1_while_C_27 : begin
        fsm_output = 10'b1100110110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_28;
      end
      COMP_LOOP_8_modExp_1_while_C_28 : begin
        fsm_output = 10'b1100110111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_29;
      end
      COMP_LOOP_8_modExp_1_while_C_29 : begin
        fsm_output = 10'b1100111000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_30;
      end
      COMP_LOOP_8_modExp_1_while_C_30 : begin
        fsm_output = 10'b1100111001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_31;
      end
      COMP_LOOP_8_modExp_1_while_C_31 : begin
        fsm_output = 10'b1100111010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_32;
      end
      COMP_LOOP_8_modExp_1_while_C_32 : begin
        fsm_output = 10'b1100111011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_33;
      end
      COMP_LOOP_8_modExp_1_while_C_33 : begin
        fsm_output = 10'b1100111100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_34;
      end
      COMP_LOOP_8_modExp_1_while_C_34 : begin
        fsm_output = 10'b1100111101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_35;
      end
      COMP_LOOP_8_modExp_1_while_C_35 : begin
        fsm_output = 10'b1100111110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_36;
      end
      COMP_LOOP_8_modExp_1_while_C_36 : begin
        fsm_output = 10'b1100111111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_37;
      end
      COMP_LOOP_8_modExp_1_while_C_37 : begin
        fsm_output = 10'b1101000000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_38;
      end
      COMP_LOOP_8_modExp_1_while_C_38 : begin
        fsm_output = 10'b1101000001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_39;
      end
      COMP_LOOP_8_modExp_1_while_C_39 : begin
        fsm_output = 10'b1101000010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_40;
      end
      COMP_LOOP_8_modExp_1_while_C_40 : begin
        fsm_output = 10'b1101000011;
        if ( COMP_LOOP_8_modExp_1_while_C_40_tr0 ) begin
          state_var_NS = COMP_LOOP_C_457;
        end
        else begin
          state_var_NS = COMP_LOOP_8_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_457 : begin
        fsm_output = 10'b1101000100;
        state_var_NS = COMP_LOOP_C_458;
      end
      COMP_LOOP_C_458 : begin
        fsm_output = 10'b1101000101;
        state_var_NS = COMP_LOOP_C_459;
      end
      COMP_LOOP_C_459 : begin
        fsm_output = 10'b1101000110;
        state_var_NS = COMP_LOOP_C_460;
      end
      COMP_LOOP_C_460 : begin
        fsm_output = 10'b1101000111;
        state_var_NS = COMP_LOOP_C_461;
      end
      COMP_LOOP_C_461 : begin
        fsm_output = 10'b1101001000;
        state_var_NS = COMP_LOOP_C_462;
      end
      COMP_LOOP_C_462 : begin
        fsm_output = 10'b1101001001;
        state_var_NS = COMP_LOOP_C_463;
      end
      COMP_LOOP_C_463 : begin
        fsm_output = 10'b1101001010;
        state_var_NS = COMP_LOOP_C_464;
      end
      COMP_LOOP_C_464 : begin
        fsm_output = 10'b1101001011;
        state_var_NS = COMP_LOOP_C_465;
      end
      COMP_LOOP_C_465 : begin
        fsm_output = 10'b1101001100;
        state_var_NS = COMP_LOOP_C_466;
      end
      COMP_LOOP_C_466 : begin
        fsm_output = 10'b1101001101;
        state_var_NS = COMP_LOOP_C_467;
      end
      COMP_LOOP_C_467 : begin
        fsm_output = 10'b1101001110;
        state_var_NS = COMP_LOOP_C_468;
      end
      COMP_LOOP_C_468 : begin
        fsm_output = 10'b1101001111;
        state_var_NS = COMP_LOOP_C_469;
      end
      COMP_LOOP_C_469 : begin
        fsm_output = 10'b1101010000;
        state_var_NS = COMP_LOOP_C_470;
      end
      COMP_LOOP_C_470 : begin
        fsm_output = 10'b1101010001;
        state_var_NS = COMP_LOOP_C_471;
      end
      COMP_LOOP_C_471 : begin
        fsm_output = 10'b1101010010;
        state_var_NS = COMP_LOOP_C_472;
      end
      COMP_LOOP_C_472 : begin
        fsm_output = 10'b1101010011;
        state_var_NS = COMP_LOOP_C_473;
      end
      COMP_LOOP_C_473 : begin
        fsm_output = 10'b1101010100;
        state_var_NS = COMP_LOOP_C_474;
      end
      COMP_LOOP_C_474 : begin
        fsm_output = 10'b1101010101;
        state_var_NS = COMP_LOOP_C_475;
      end
      COMP_LOOP_C_475 : begin
        fsm_output = 10'b1101010110;
        state_var_NS = COMP_LOOP_C_476;
      end
      COMP_LOOP_C_476 : begin
        fsm_output = 10'b1101010111;
        state_var_NS = COMP_LOOP_C_477;
      end
      COMP_LOOP_C_477 : begin
        fsm_output = 10'b1101011000;
        state_var_NS = COMP_LOOP_C_478;
      end
      COMP_LOOP_C_478 : begin
        fsm_output = 10'b1101011001;
        state_var_NS = COMP_LOOP_C_479;
      end
      COMP_LOOP_C_479 : begin
        fsm_output = 10'b1101011010;
        state_var_NS = COMP_LOOP_C_480;
      end
      COMP_LOOP_C_480 : begin
        fsm_output = 10'b1101011011;
        state_var_NS = COMP_LOOP_C_481;
      end
      COMP_LOOP_C_481 : begin
        fsm_output = 10'b1101011100;
        state_var_NS = COMP_LOOP_C_482;
      end
      COMP_LOOP_C_482 : begin
        fsm_output = 10'b1101011101;
        state_var_NS = COMP_LOOP_C_483;
      end
      COMP_LOOP_C_483 : begin
        fsm_output = 10'b1101011110;
        state_var_NS = COMP_LOOP_C_484;
      end
      COMP_LOOP_C_484 : begin
        fsm_output = 10'b1101011111;
        state_var_NS = COMP_LOOP_C_485;
      end
      COMP_LOOP_C_485 : begin
        fsm_output = 10'b1101100000;
        state_var_NS = COMP_LOOP_C_486;
      end
      COMP_LOOP_C_486 : begin
        fsm_output = 10'b1101100001;
        state_var_NS = COMP_LOOP_C_487;
      end
      COMP_LOOP_C_487 : begin
        fsm_output = 10'b1101100010;
        state_var_NS = COMP_LOOP_C_488;
      end
      COMP_LOOP_C_488 : begin
        fsm_output = 10'b1101100011;
        state_var_NS = COMP_LOOP_C_489;
      end
      COMP_LOOP_C_489 : begin
        fsm_output = 10'b1101100100;
        state_var_NS = COMP_LOOP_C_490;
      end
      COMP_LOOP_C_490 : begin
        fsm_output = 10'b1101100101;
        state_var_NS = COMP_LOOP_C_491;
      end
      COMP_LOOP_C_491 : begin
        fsm_output = 10'b1101100110;
        state_var_NS = COMP_LOOP_C_492;
      end
      COMP_LOOP_C_492 : begin
        fsm_output = 10'b1101100111;
        state_var_NS = COMP_LOOP_C_493;
      end
      COMP_LOOP_C_493 : begin
        fsm_output = 10'b1101101000;
        state_var_NS = COMP_LOOP_C_494;
      end
      COMP_LOOP_C_494 : begin
        fsm_output = 10'b1101101001;
        state_var_NS = COMP_LOOP_C_495;
      end
      COMP_LOOP_C_495 : begin
        fsm_output = 10'b1101101010;
        state_var_NS = COMP_LOOP_C_496;
      end
      COMP_LOOP_C_496 : begin
        fsm_output = 10'b1101101011;
        state_var_NS = COMP_LOOP_C_497;
      end
      COMP_LOOP_C_497 : begin
        fsm_output = 10'b1101101100;
        state_var_NS = COMP_LOOP_C_498;
      end
      COMP_LOOP_C_498 : begin
        fsm_output = 10'b1101101101;
        state_var_NS = COMP_LOOP_C_499;
      end
      COMP_LOOP_C_499 : begin
        fsm_output = 10'b1101101110;
        state_var_NS = COMP_LOOP_C_500;
      end
      COMP_LOOP_C_500 : begin
        fsm_output = 10'b1101101111;
        state_var_NS = COMP_LOOP_C_501;
      end
      COMP_LOOP_C_501 : begin
        fsm_output = 10'b1101110000;
        state_var_NS = COMP_LOOP_C_502;
      end
      COMP_LOOP_C_502 : begin
        fsm_output = 10'b1101110001;
        state_var_NS = COMP_LOOP_C_503;
      end
      COMP_LOOP_C_503 : begin
        fsm_output = 10'b1101110010;
        state_var_NS = COMP_LOOP_C_504;
      end
      COMP_LOOP_C_504 : begin
        fsm_output = 10'b1101110011;
        state_var_NS = COMP_LOOP_C_505;
      end
      COMP_LOOP_C_505 : begin
        fsm_output = 10'b1101110100;
        state_var_NS = COMP_LOOP_C_506;
      end
      COMP_LOOP_C_506 : begin
        fsm_output = 10'b1101110101;
        state_var_NS = COMP_LOOP_C_507;
      end
      COMP_LOOP_C_507 : begin
        fsm_output = 10'b1101110110;
        state_var_NS = COMP_LOOP_C_508;
      end
      COMP_LOOP_C_508 : begin
        fsm_output = 10'b1101110111;
        state_var_NS = COMP_LOOP_C_509;
      end
      COMP_LOOP_C_509 : begin
        fsm_output = 10'b1101111000;
        state_var_NS = COMP_LOOP_C_510;
      end
      COMP_LOOP_C_510 : begin
        fsm_output = 10'b1101111001;
        state_var_NS = COMP_LOOP_C_511;
      end
      COMP_LOOP_C_511 : begin
        fsm_output = 10'b1101111010;
        state_var_NS = COMP_LOOP_C_512;
      end
      COMP_LOOP_C_512 : begin
        fsm_output = 10'b1101111011;
        state_var_NS = COMP_LOOP_C_513;
      end
      COMP_LOOP_C_513 : begin
        fsm_output = 10'b1101111100;
        state_var_NS = COMP_LOOP_C_514;
      end
      COMP_LOOP_C_514 : begin
        fsm_output = 10'b1101111101;
        state_var_NS = COMP_LOOP_C_515;
      end
      COMP_LOOP_C_515 : begin
        fsm_output = 10'b1101111110;
        state_var_NS = COMP_LOOP_C_516;
      end
      COMP_LOOP_C_516 : begin
        fsm_output = 10'b1101111111;
        state_var_NS = COMP_LOOP_C_517;
      end
      COMP_LOOP_C_517 : begin
        fsm_output = 10'b1110000000;
        state_var_NS = COMP_LOOP_C_518;
      end
      COMP_LOOP_C_518 : begin
        fsm_output = 10'b1110000001;
        state_var_NS = COMP_LOOP_C_519;
      end
      COMP_LOOP_C_519 : begin
        fsm_output = 10'b1110000010;
        state_var_NS = COMP_LOOP_C_520;
      end
      COMP_LOOP_C_520 : begin
        fsm_output = 10'b1110000011;
        if ( COMP_LOOP_C_520_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 10'b1110000100;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_9;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_9 : begin
        fsm_output = 10'b1110000101;
        if ( STAGE_LOOP_C_9_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 10'b1110000110;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 10'b0000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d, vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_adra_d_pff, vec_rsc_0_0_i_da_d_pff,
      vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff, vec_rsc_0_2_i_wea_d_pff,
      vec_rsc_0_3_i_wea_d_pff, vec_rsc_0_4_i_wea_d_pff, vec_rsc_0_5_i_wea_d_pff,
      vec_rsc_0_6_i_wea_d_pff, vec_rsc_0_7_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_qa_d;
  output vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_qa_d;
  output vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_qa_d;
  output vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_qa_d;
  output vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_qa_d;
  output vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_qa_d;
  output vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [8:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;
  output vec_rsc_0_2_i_wea_d_pff;
  output vec_rsc_0_3_i_wea_d_pff;
  output vec_rsc_0_4_i_wea_d_pff;
  output vec_rsc_0_5_i_wea_d_pff;
  output vec_rsc_0_6_i_wea_d_pff;
  output vec_rsc_0_7_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  reg [63:0] modulo_result_rem_cmp_a;
  reg [63:0] modulo_result_rem_cmp_b;
  wire [63:0] modulo_result_rem_cmp_z;
  reg [64:0] operator_66_true_div_cmp_a;
  wire [64:0] operator_66_true_div_cmp_z;
  reg [9:0] operator_66_true_div_cmp_b_9_0;
  wire [9:0] fsm_output;
  wire or_dcpl_3;
  wire or_tmp_5;
  wire or_tmp_9;
  wire or_tmp_13;
  wire not_tmp_29;
  wire or_tmp_58;
  wire or_tmp_60;
  wire mux_tmp_77;
  wire or_tmp_63;
  wire not_tmp_46;
  wire mux_tmp_81;
  wire mux_tmp_83;
  wire nor_tmp_12;
  wire and_tmp_2;
  wire or_tmp_71;
  wire or_tmp_72;
  wire or_tmp_73;
  wire nor_tmp_13;
  wire mux_tmp_164;
  wire nor_tmp_21;
  wire not_tmp_82;
  wire mux_tmp_229;
  wire mux_tmp_390;
  wire not_tmp_121;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire and_dcpl_18;
  wire and_dcpl_23;
  wire and_dcpl_26;
  wire and_dcpl_33;
  wire not_tmp_129;
  wire and_dcpl_49;
  wire and_dcpl_50;
  wire and_dcpl_53;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_61;
  wire or_dcpl_39;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire and_dcpl_75;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_98;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_122;
  wire and_dcpl_124;
  wire and_dcpl_126;
  wire and_dcpl_133;
  wire and_dcpl_134;
  wire mux_tmp_469;
  wire not_tmp_166;
  wire mux_tmp_472;
  wire mux_tmp_473;
  wire mux_tmp_488;
  wire not_tmp_170;
  wire not_tmp_171;
  wire mux_tmp_504;
  wire not_tmp_177;
  wire not_tmp_178;
  wire mux_tmp_523;
  wire mux_tmp_539;
  wire not_tmp_189;
  wire mux_tmp_542;
  wire not_tmp_190;
  wire mux_tmp_558;
  wire mux_tmp_574;
  wire not_tmp_201;
  wire not_tmp_202;
  wire mux_tmp_593;
  wire mux_tmp_609;
  wire not_tmp_214;
  wire mux_tmp_616;
  wire mux_tmp_620;
  wire mux_tmp_628;
  wire mux_tmp_644;
  wire not_tmp_225;
  wire not_tmp_226;
  wire mux_tmp_663;
  wire mux_tmp_679;
  wire not_tmp_237;
  wire mux_tmp_686;
  wire not_tmp_239;
  wire mux_tmp_698;
  wire mux_tmp_714;
  wire not_tmp_249;
  wire not_tmp_250;
  wire mux_tmp_733;
  wire and_dcpl_150;
  wire or_tmp_672;
  wire or_tmp_677;
  wire or_tmp_679;
  wire nor_tmp_166;
  wire or_tmp_681;
  wire mux_tmp_760;
  wire or_tmp_682;
  wire mux_tmp_773;
  wire mux_tmp_777;
  wire nor_tmp_168;
  wire not_tmp_276;
  wire mux_tmp_814;
  wire mux_tmp_823;
  wire mux_tmp_825;
  wire mux_tmp_833;
  wire or_tmp_737;
  wire mux_tmp_860;
  wire or_tmp_738;
  wire mux_tmp_865;
  wire and_dcpl_151;
  wire not_tmp_309;
  wire and_dcpl_152;
  wire and_dcpl_156;
  wire and_dcpl_157;
  wire mux_tmp_898;
  wire mux_tmp_899;
  wire mux_tmp_900;
  wire or_tmp_783;
  wire mux_tmp_912;
  wire mux_tmp_1013;
  wire or_dcpl_56;
  wire mux_tmp_1037;
  wire nor_tmp_223;
  wire and_dcpl_174;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire not_tmp_375;
  wire or_dcpl_62;
  wire not_tmp_384;
  wire or_tmp_966;
  wire not_tmp_390;
  wire or_tmp_970;
  wire or_tmp_992;
  wire or_tmp_993;
  wire mux_tmp_1175;
  wire mux_tmp_1179;
  wire mux_tmp_1182;
  wire mux_tmp_1184;
  wire mux_tmp_1187;
  wire mux_tmp_1189;
  wire mux_tmp_1190;
  wire mux_tmp_1191;
  wire mux_tmp_1192;
  wire mux_tmp_1199;
  wire mux_tmp_1203;
  wire not_tmp_414;
  wire mux_tmp_1208;
  wire or_tmp_1034;
  wire and_dcpl_191;
  wire or_tmp_1050;
  wire mux_tmp_1272;
  wire mux_tmp_1276;
  wire mux_tmp_1277;
  wire mux_tmp_1288;
  wire and_dcpl_192;
  wire and_dcpl_194;
  wire not_tmp_458;
  wire mux_tmp_1329;
  wire mux_tmp_1331;
  wire mux_tmp_1332;
  wire or_tmp_1128;
  wire mux_tmp_1341;
  wire mux_tmp_1345;
  wire mux_tmp_1348;
  wire mux_tmp_1351;
  wire or_tmp_1137;
  wire mux_tmp_1353;
  wire mux_tmp_1355;
  wire or_tmp_1142;
  wire not_tmp_496;
  wire or_tmp_1157;
  reg COMP_LOOP_COMP_LOOP_and_11_itm;
  reg COMP_LOOP_COMP_LOOP_and_2_itm;
  reg [5:0] COMP_LOOP_k_9_3_sva_5_0;
  reg [11:0] VEC_LOOP_j_sva_11_0;
  reg COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  reg operator_64_false_slc_modExp_exp_0_1_itm;
  reg [11:0] COMP_LOOP_acc_10_cse_12_1_1_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_4_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_6_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_6_sva;
  reg [10:0] COMP_LOOP_acc_11_psp_sva;
  reg [10:0] COMP_LOOP_acc_14_psp_sva;
  reg [9:0] COMP_LOOP_acc_13_psp_sva;
  wire [11:0] COMP_LOOP_acc_1_cse_2_sva_1;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_2_sva_1;
  wire modExp_while_and_1_rgt;
  wire and_244_m1c;
  wire and_250_m1c;
  wire and_185_m1c;
  wire or_294_cse;
  wire nor_115_cse;
  wire or_521_cse;
  wire and_336_cse;
  reg reg_vec_rsc_triosy_0_7_obj_ld_cse;
  wire and_316_cse;
  wire or_722_cse;
  wire or_730_cse;
  wire nor_397_cse;
  wire nor_398_cse;
  wire or_857_cse;
  wire nand_82_cse;
  wire or_1161_cse;
  wire nor_400_cse;
  wire [63:0] modulo_result_mux_1_cse;
  wire and_293_cse;
  wire and_398_cse;
  wire and_292_cse;
  wire or_831_cse;
  wire or_91_cse;
  wire or_90_cse;
  wire nor_401_cse;
  wire or_5_cse;
  wire or_217_cse;
  wire or_157_cse;
  wire nand_245_cse;
  wire nor_265_cse;
  wire mux_483_cse;
  wire nand_232_cse;
  wire or_1379_cse;
  wire or_277_cse;
  wire nor_112_cse;
  wire nor_114_cse;
  wire nor_122_cse;
  wire mux_995_cse;
  wire and_434_cse;
  wire or_29_cse;
  wire and_312_cse;
  wire or_823_cse;
  wire or_843_cse;
  wire nor_692_cse;
  wire or_1275_cse;
  wire and_433_cse;
  wire or_1156_cse;
  wire or_119_cse;
  wire nand_240_cse;
  wire or_731_cse;
  wire nor_365_cse;
  wire mux_477_cse;
  wire nor_624_cse;
  wire nor_594_cse;
  wire mux_445_cse;
  wire nand_244_cse;
  wire mux_417_cse;
  wire mux_903_cse;
  wire mux_919_cse;
  wire mux_923_cse;
  wire mux_929_cse;
  wire mux_937_cse;
  wire COMP_LOOP_nor_97_cse;
  wire mux_446_cse;
  wire mux_438_cse;
  wire mux_928_cse;
  wire mux_82_cse;
  wire mux_1026_cse;
  wire [8:0] COMP_LOOP_acc_psp_sva_1;
  wire [9:0] nl_COMP_LOOP_acc_psp_sva_1;
  reg [8:0] COMP_LOOP_acc_psp_sva;
  wire mux_453_itm;
  wire mux_1151_itm;
  wire mux_1209_itm;
  wire mux_1289_itm;
  wire and_dcpl_218;
  wire and_dcpl_223;
  wire not_tmp_519;
  wire mux_tmp_1422;
  wire mux_tmp_1425;
  wire not_tmp_524;
  wire [63:0] z_out;
  wire [127:0] nl_z_out;
  wire [12:0] z_out_1;
  wire [13:0] nl_z_out_1;
  wire and_dcpl_246;
  wire nor_tmp_272;
  wire and_dcpl_247;
  wire and_dcpl_248;
  wire and_dcpl_256;
  wire and_dcpl_262;
  wire [64:0] z_out_2;
  wire and_dcpl_265;
  wire and_dcpl_267;
  wire and_dcpl_271;
  wire and_dcpl_277;
  wire and_dcpl_278;
  wire and_dcpl_280;
  wire and_dcpl_284;
  wire and_dcpl_289;
  wire [7:0] z_out_3;
  wire and_dcpl_291;
  wire and_dcpl_298;
  wire and_dcpl_300;
  wire and_dcpl_305;
  wire and_dcpl_309;
  wire and_dcpl_312;
  wire and_dcpl_313;
  wire and_dcpl_318;
  wire and_dcpl_324;
  wire and_dcpl_326;
  wire and_dcpl_330;
  wire [9:0] z_out_4;
  wire and_dcpl_342;
  wire and_dcpl_355;
  wire and_dcpl_359;
  wire and_dcpl_360;
  wire and_dcpl_410;
  wire and_dcpl_411;
  wire and_dcpl_442;
  wire [64:0] z_out_7;
  wire [65:0] nl_z_out_7;
  wire and_dcpl_451;
  wire and_dcpl_460;
  wire and_dcpl_467;
  wire [63:0] z_out_8;
  wire [64:0] nl_z_out_8;
  reg [63:0] p_sva;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg [63:0] modExp_base_sva;
  reg [63:0] modExp_result_sva;
  reg modExp_exp_1_7_1_sva;
  reg modExp_exp_1_6_1_sva;
  reg modExp_exp_1_5_1_sva;
  reg modExp_exp_1_4_1_sva;
  reg modExp_exp_1_3_1_sva;
  reg modExp_exp_1_2_1_sva;
  reg modExp_exp_1_1_1_sva;
  reg modExp_exp_1_0_1_sva_1;
  reg [63:0] tmp_10_lpi_4_dfm;
  reg [63:0] COMP_LOOP_1_mul_mut;
  reg [62:0] operator_64_false_slc_modExp_exp_63_1_itm;
  reg COMP_LOOP_COMP_LOOP_nor_itm;
  reg COMP_LOOP_COMP_LOOP_and_4_itm;
  reg COMP_LOOP_COMP_LOOP_and_5_itm;
  reg COMP_LOOP_COMP_LOOP_and_6_itm;
  reg COMP_LOOP_COMP_LOOP_nor_1_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg [63:0] COMP_LOOP_1_acc_8_itm;
  reg COMP_LOOP_COMP_LOOP_and_30_itm;
  reg COMP_LOOP_COMP_LOOP_and_32_itm;
  reg COMP_LOOP_COMP_LOOP_and_58_itm;
  reg COMP_LOOP_COMP_LOOP_and_124_itm;
  reg COMP_LOOP_COMP_LOOP_and_125_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [3:0] STAGE_LOOP_i_3_0_sva_2;
  wire [4:0] nl_STAGE_LOOP_i_3_0_sva_2;
  wire [63:0] COMP_LOOP_1_acc_5_mut_mx0w5;
  wire [64:0] nl_COMP_LOOP_1_acc_5_mut_mx0w5;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire VEC_LOOP_j_sva_11_0_mx0c1;
  wire modExp_result_sva_mx0c0;
  wire modExp_base_sva_mx0c1;
  wire [63:0] modulo_qr_sva_1_mx1w1;
  wire [64:0] nl_modulo_qr_sva_1_mx1w1;
  wire [62:0] operator_64_false_slc_modExp_exp_63_1_3;
  wire tmp_10_lpi_4_dfm_mx0c1;
  wire tmp_10_lpi_4_dfm_mx0c2;
  wire tmp_10_lpi_4_dfm_mx0c3;
  wire tmp_10_lpi_4_dfm_mx0c4;
  wire tmp_10_lpi_4_dfm_mx0c5;
  wire tmp_10_lpi_4_dfm_mx0c6;
  wire tmp_10_lpi_4_dfm_mx0c7;
  wire COMP_LOOP_COMP_LOOP_and_211;
  wire COMP_LOOP_COMP_LOOP_and_213;
  wire COMP_LOOP_COMP_LOOP_and_215;
  wire and_243_m1c;
  wire modExp_result_and_rgt;
  wire modExp_result_and_1_rgt;
  reg [62:0] modExp_exp_sva_rsp_1;
  wire COMP_LOOP_COMP_LOOP_and_11_cse;
  wire modExp_while_or_1_cse;
  wire COMP_LOOP_COMP_LOOP_and_12_cse;
  wire COMP_LOOP_COMP_LOOP_and_37_cse;
  wire COMP_LOOP_COMP_LOOP_and_13_cse;
  wire COMP_LOOP_or_3_cse;
  wire or_718_cse;
  wire or_1312_cse;
  wire or_798_cse;
  wire nor_tmp_273;
  wire mux_tmp_1456;
  wire or_tmp_1262;
  wire or_tmp_1267;
  wire or_tmp_1269;
  wire or_tmp_1273;
  wire or_tmp_1274;
  wire not_tmp_621;
  wire [64:0] operator_64_false_operator_64_false_mux_rgt;
  reg operator_64_false_acc_mut_64;
  reg [63:0] operator_64_false_acc_mut_63_0;
  wire or_1470_cse;
  wire or_1516_cse;
  wire and_721_cse;
  wire or_1483_cse;
  wire nor_813_cse;
  wire and_303_cse;
  wire or_750_cse;
  wire nor_820_cse;
  wire mux_1001_cse;
  wire mux_1014_cse;
  wire mux_1460_cse;
  wire mux_936_cse;
  wire mux_1447_cse;
  wire COMP_LOOP_or_39_itm;
  wire operator_64_false_1_nor_1_itm;
  wire COMP_LOOP_or_43_itm;
  wire STAGE_LOOP_acc_itm_2_1;
  wire [11:0] z_out_6_12_1;
  wire nor_379_cse;
  wire nor_797_cse;

  wire[0:0] or_1380_nl;
  wire[0:0] or_1381_nl;
  wire[0:0] modulo_result_or_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] or_767_nl;
  wire[0:0] or_766_nl;
  wire[0:0] or_764_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] mux_851_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] mux_850_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] mux_849_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] mux_802_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] or_733_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] mux_793_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] mux_787_nl;
  wire[0:0] mux_786_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] mux_783_nl;
  wire[0:0] mux_782_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] mux_780_nl;
  wire[0:0] mux_779_nl;
  wire[0:0] mux_778_nl;
  wire[0:0] mux_776_nl;
  wire[0:0] mux_775_nl;
  wire[0:0] or_728_nl;
  wire[0:0] mux_774_nl;
  wire[0:0] or_727_nl;
  wire[0:0] mux_771_nl;
  wire[0:0] mux_770_nl;
  wire[0:0] mux_769_nl;
  wire[0:0] mux_768_nl;
  wire[0:0] mux_767_nl;
  wire[0:0] or_726_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] mux_765_nl;
  wire[0:0] mux_764_nl;
  wire[0:0] mux_763_nl;
  wire[0:0] mux_762_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] mux_759_nl;
  wire[0:0] mux_758_nl;
  wire[0:0] mux_757_nl;
  wire[0:0] mux_756_nl;
  wire[0:0] mux_755_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] mux_753_nl;
  wire[0:0] mux_752_nl;
  wire[0:0] or_716_nl;
  wire[0:0] mux_751_nl;
  wire[0:0] mux_750_nl;
  wire[0:0] or_715_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] mux_845_nl;
  wire[0:0] mux_844_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] mux_842_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] or_754_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] or_753_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] mux_836_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] or_751_nl;
  wire[0:0] mux_832_nl;
  wire[0:0] or_748_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] mux_829_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] mux_826_nl;
  wire[0:0] or_745_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] mux_818_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] mux_813_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] or_740_nl;
  wire[0:0] mux_811_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] mux_809_nl;
  wire[0:0] nand_127_nl;
  wire[0:0] or_737_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] mux_879_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] mux_877_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] mux_876_nl;
  wire[0:0] mux_875_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] mux_874_nl;
  wire[0:0] mux_873_nl;
  wire[0:0] mux_872_nl;
  wire[0:0] or_789_nl;
  wire[0:0] or_788_nl;
  wire[0:0] mux_871_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] mux_868_nl;
  wire[0:0] mux_867_nl;
  wire[0:0] nor_383_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] mux_861_nl;
  wire[0:0] and_304_nl;
  wire[0:0] and_305_nl;
  wire[0:0] and_306_nl;
  wire[0:0] and_307_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] and_446_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] and_56_nl;
  wire[0:0] and_55_nl;
  wire[0:0] and_57_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] and_54_nl;
  wire[63:0] modExp_while_if_mux1h_nl;
  wire[0:0] modExp_while_if_or_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] nor_333_nl;
  wire[0:0] nor_335_nl;
  wire[0:0] nor_336_nl;
  wire[0:0] and_274_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] and_275_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] nor_337_nl;
  wire[0:0] nor_338_nl;
  wire[0:0] nor_339_nl;
  wire[0:0] modExp_1_while_and_16_nl;
  wire[0:0] modExp_1_while_and_18_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] mux_1005_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] mux_1000_nl;
  wire[0:0] mux_999_nl;
  wire[0:0] mux_998_nl;
  wire[0:0] mux_997_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] mux_992_nl;
  wire[0:0] mux_991_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] mux_989_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] and_176_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] mux_978_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] mux_973_nl;
  wire[0:0] mux_972_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] mux_968_nl;
  wire[0:0] mux_967_nl;
  wire[0:0] mux_966_nl;
  wire[0:0] mux_965_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] mux_963_nl;
  wire[0:0] mux_962_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] or_1466_nl;
  wire[0:0] mux_1493_nl;
  wire[0:0] mux_1492_nl;
  wire[0:0] mux_1491_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] mux_1489_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] mux_1487_nl;
  wire[0:0] nor_815_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] mux_1485_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] mux_1483_nl;
  wire[0:0] nor_835_nl;
  wire[0:0] or_1473_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] nor_836_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] and_720_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] mux_1459_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] mux_1519_nl;
  wire[0:0] mux_1518_nl;
  wire[0:0] mux_1517_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] nor_828_nl;
  wire[0:0] and_715_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] nor_829_nl;
  wire[0:0] nor_830_nl;
  wire[0:0] and_716_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] or_1504_nl;
  wire[0:0] nor_831_nl;
  wire[0:0] mux_1512_nl;
  wire[0:0] mux_1511_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] mux_1509_nl;
  wire[0:0] and_717_nl;
  wire[0:0] or_1502_nl;
  wire[0:0] and_718_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] nand_268_nl;
  wire[0:0] or_1498_nl;
  wire[0:0] mux_1506_nl;
  wire[0:0] mux_1505_nl;
  wire[0:0] or_1494_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] or_1492_nl;
  wire[0:0] mux_1503_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] nor_832_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] nor_834_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] mux_1500_nl;
  wire[0:0] mux_1499_nl;
  wire[0:0] or_1485_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] or_1484_nl;
  wire[0:0] or_1481_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] or_1478_nl;
  wire[0:0] mux_1495_nl;
  wire[0:0] mux_1494_nl;
  wire[0:0] or_1476_nl;
  wire[0:0] or_844_nl;
  wire[0:0] or_1460_nl;
  wire[0:0] mux_1015_nl;
  wire[0:0] or_845_nl;
  wire[0:0] or_841_nl;
  wire[0:0] mux_1522_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] nor_826_nl;
  wire[0:0] nor_827_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] mux_1029_nl;
  wire[0:0] and_286_nl;
  wire[0:0] or_864_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] nor_327_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] nor_329_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] or_982_nl;
  wire[0:0] or_980_nl;
  wire[0:0] nor_330_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] mux_56_nl;
  wire[0:0] nand_238_nl;
  wire[0:0] mux_55_nl;
  wire[0:0] nor_721_nl;
  wire[0:0] nor_722_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_2_nl;
  wire[9:0] COMP_LOOP_1_acc_nl;
  wire[10:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] nor_808_nl;
  wire[0:0] and_714_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] or_1266_nl;
  wire[0:0] nor_323_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] or_1025_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] or_1032_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] nand_112_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] and_208_nl;
  wire[0:0] and_207_nl;
  wire[0:0] or_1038_nl;
  wire[0:0] or_1043_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] and_211_nl;
  wire[0:0] and_210_nl;
  wire[0:0] and_212_nl;
  wire[0:0] and_214_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] or_1046_nl;
  wire[0:0] or_1045_nl;
  wire[0:0] operator_64_false_1_mux1h_nl;
  wire[0:0] operator_64_false_1_or_2_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] or_1066_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] or_1064_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] or_1063_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] nor_318_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] or_1401_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] or_964_nl;
  wire[0:0] or_1052_nl;
  wire[0:0] nand_243_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] nor_320_nl;
  wire[0:0] nor_321_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] and_267_nl;
  wire[0:0] mux_1214_nl;
  wire[0:0] nor_314_nl;
  wire[0:0] nor_315_nl;
  wire[0:0] and_268_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] nor_316_nl;
  wire[0:0] nor_317_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] nor_308_nl;
  wire[0:0] nor_309_nl;
  wire[0:0] COMP_LOOP_mux_42_nl;
  wire[0:0] and_222_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] nand_109_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] or_1103_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] or_1101_nl;
  wire[0:0] or_1100_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] or_1098_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] nor_312_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] or_1078_nl;
  wire[0:0] or_1077_nl;
  wire[0:0] nor_313_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] or_1074_nl;
  wire[0:0] or_1073_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] nand_242_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] nor_305_nl;
  wire[0:0] nor_306_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] or_1109_nl;
  wire[0:0] or_1108_nl;
  wire[0:0] or_1400_nl;
  wire[0:0] COMP_LOOP_mux1h_32_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] and_259_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] nor_299_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] nor_300_nl;
  wire[0:0] nor_301_nl;
  wire[0:0] nor_302_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] or_1119_nl;
  wire[0:0] COMP_LOOP_mux1h_46_nl;
  wire[0:0] COMP_LOOP_mux1h_48_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] mux_1307_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] nand_192_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] nor_296_nl;
  wire[0:0] nor_297_nl;
  wire[0:0] or_1300_nl;
  wire[0:0] mux_1309_nl;
  wire[0:0] nand_106_nl;
  wire[0:0] or_1140_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] or_1308_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] or_1154_nl;
  wire[0:0] or_1152_nl;
  wire[0:0] or_1309_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] or_1150_nl;
  wire[0:0] or_1148_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] or_1168_nl;
  wire[0:0] nand_86_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] nor_292_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] or_1166_nl;
  wire[0:0] or_1165_nl;
  wire[0:0] nor_293_nl;
  wire[0:0] or_1162_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] mux_1316_nl;
  wire[0:0] or_1160_nl;
  wire[0:0] or_1158_nl;
  wire[0:0] mux_1315_nl;
  wire[0:0] or_1157_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_or_17_nl;
  wire[0:0] COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_or_19_nl;
  wire[0:0] COMP_LOOP_or_20_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire[0:0] COMP_LOOP_or_26_nl;
  wire[0:0] COMP_LOOP_or_27_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] nor_746_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] mux_71_nl;
  wire[0:0] or_1391_nl;
  wire[0:0] or_1392_nl;
  wire[0:0] or_1393_nl;
  wire[0:0] or_1394_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] or_1395_nl;
  wire[0:0] mux_69_nl;
  wire[0:0] or_1396_nl;
  wire[0:0] or_1397_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] or_56_nl;
  wire[0:0] or_54_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] mux_1380_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] mux_1378_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] mux_1375_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] mux_1370_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] mux_1368_nl;
  wire[0:0] mux_1367_nl;
  wire[0:0] and_253_nl;
  wire[0:0] mux_1366_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] mux_1364_nl;
  wire[0:0] or_1207_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] or_1206_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] mux_1356_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] or_1201_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] or_1196_nl;
  wire[0:0] nand_98_nl;
  wire[0:0] or_1192_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] or_1191_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] nand_183_nl;
  wire[0:0] and_432_nl;
  wire[0:0] and_60_nl;
  wire[0:0] or_263_nl;
  wire[0:0] or_261_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] or_270_nl;
  wire[0:0] or_269_nl;
  wire[0:0] or_275_nl;
  wire[0:0] or_273_nl;
  wire[0:0] or_1376_nl;
  wire[0:0] or_1377_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] nor_630_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] or_297_nl;
  wire[0:0] or_296_nl;
  wire[0:0] or_324_nl;
  wire[0:0] or_322_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] nor_609_nl;
  wire[0:0] or_355_nl;
  wire[0:0] or_354_nl;
  wire[0:0] or_382_nl;
  wire[0:0] or_380_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] or_389_nl;
  wire[0:0] or_388_nl;
  wire[0:0] nor_578_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] or_412_nl;
  wire[0:0] or_411_nl;
  wire[0:0] or_438_nl;
  wire[0:0] or_436_nl;
  wire[0:0] nor_550_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] or_465_nl;
  wire[0:0] or_464_nl;
  wire[0:0] or_490_nl;
  wire[0:0] or_488_nl;
  wire[0:0] nor_520_nl;
  wire[0:0] nor_521_nl;
  wire[0:0] or_504_nl;
  wire[0:0] or_503_nl;
  wire[0:0] or_514_nl;
  wire[0:0] or_512_nl;
  wire[0:0] or_524_nl;
  wire[0:0] or_523_nl;
  wire[0:0] or_550_nl;
  wire[0:0] or_548_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] or_581_nl;
  wire[0:0] or_580_nl;
  wire[0:0] or_607_nl;
  wire[0:0] or_605_nl;
  wire[0:0] nor_460_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] or_621_nl;
  wire[0:0] or_620_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] or_637_nl;
  wire[0:0] or_636_nl;
  wire[0:0] or_662_nl;
  wire[0:0] nand_136_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] and_447_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] nand_131_nl;
  wire[0:0] or_688_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] and_310_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] nand_194_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] and_301_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] or_1313_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] or_797_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] nor_375_nl;
  wire[0:0] nor_376_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] and_298_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] or_811_nl;
  wire[0:0] nand_69_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] and_299_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] mux_894_nl;
  wire[0:0] nor_750_nl;
  wire[0:0] and_296_nl;
  wire[0:0] nand_191_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] or_953_nl;
  wire[0:0] or_952_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] nor_670_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] or_946_nl;
  wire[0:0] or_945_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] and_198_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] or_1017_nl;
  wire[0:0] or_1015_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] or_1062_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] mux_1206_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] or_73_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] mux_1302_nl;
  wire[0:0] mux_1301_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] or_1132_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] or_1199_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] nor_282_nl;
  wire[0:0] and_256_nl;
  wire[0:0] and_251_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] and_252_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] nor_277_nl;
  wire[0:0] nor_278_nl;
  wire[0:0] nor_279_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] or_1215_nl;
  wire[0:0] or_1214_nl;
  wire[0:0] nor_280_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] or_1212_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] nand_182_nl;
  wire[0:0] or_1209_nl;
  wire[0:0] mux_1025_nl;
  wire[0:0] mux_1024_nl;
  wire[0:0] mux_1023_nl;
  wire[0:0] or_859_nl;
  wire[2:0] STAGE_LOOP_acc_nl;
  wire[3:0] nl_STAGE_LOOP_acc_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] nor_273_nl;
  wire[0:0] mux_1395_nl;
  wire[0:0] nand_89_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] nor_274_nl;
  wire[0:0] nor_275_nl;
  wire[0:0] or_1228_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] or_1227_nl;
  wire[0:0] nor_276_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] or_1224_nl;
  wire[0:0] or_1222_nl;
  wire[0:0] and_98_nl;
  wire[0:0] nor_740_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] nand_235_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] or_1386_nl;
  wire[0:0] or_1387_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] or_1388_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] or_234_nl;
  wire[0:0] or_233_nl;
  wire[0:0] or_232_nl;
  wire[0:0] or_1389_nl;
  wire[0:0] and_103_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] and_110_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] and_116_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] and_121_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] and_449_nl;
  wire[0:0] and_127_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] and_135_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] and_145_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] and_382_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] mux_487_nl;
  wire[0:0] mux_486_nl;
  wire[0:0] mux_485_nl;
  wire[0:0] mux_484_nl;
  wire[0:0] or_1375_nl;
  wire[0:0] mux_482_nl;
  wire[0:0] or_1378_nl;
  wire[0:0] mux_480_nl;
  wire[0:0] mux_479_nl;
  wire[0:0] nand_233_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] or_1382_nl;
  wire[0:0] mux_476_nl;
  wire[0:0] mux_475_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] or_1383_nl;
  wire[0:0] or_1384_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] nand_234_nl;
  wire[0:0] or_1385_nl;
  wire[0:0] or_260_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] mux_501_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] nor_612_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] and_377_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] mux_497_nl;
  wire[0:0] nor_617_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] or_311_nl;
  wire[0:0] or_309_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] and_378_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] mux_491_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] or_1366_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] nand_228_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] nand_229_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] or_1372_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] mux_509_nl;
  wire[0:0] or_1373_nl;
  wire[0:0] nand_230_nl;
  wire[0:0] mux_506_nl;
  wire[0:0] nand_231_nl;
  wire[0:0] or_1374_nl;
  wire[0:0] or_321_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] mux_535_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] and_370_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] nor_588_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] or_369_nl;
  wire[0:0] or_367_nl;
  wire[0:0] mux_530_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] and_371_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] nor_590_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] mux_554_nl;
  wire[0:0] nand_222_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] or_1359_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] nand_224_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] or_1363_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] nand_225_nl;
  wire[0:0] or_1364_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] nand_226_nl;
  wire[0:0] or_1365_nl;
  wire[0:0] or_379_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] mux_570_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] nor_553_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] and_363_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] mux_566_nl;
  wire[0:0] or_425_nl;
  wire[0:0] or_423_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] mux_564_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] and_364_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] nor_560_nl;
  wire[0:0] nor_561_nl;
  wire[0:0] nor_562_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] nor_564_nl;
  wire[0:0] nor_566_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] mux_590_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] nand_215_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] nand_217_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] nand_218_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] or_1355_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] mux_579_nl;
  wire[0:0] nand_219_nl;
  wire[0:0] nand_220_nl;
  wire[0:0] mux_576_nl;
  wire[0:0] nand_221_nl;
  wire[0:0] or_1356_nl;
  wire[0:0] or_435_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] nor_522_nl;
  wire[0:0] nor_523_nl;
  wire[0:0] nor_524_nl;
  wire[0:0] and_354_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] nor_525_nl;
  wire[0:0] nor_526_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] nor_527_nl;
  wire[0:0] nor_528_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] or_478_nl;
  wire[0:0] or_476_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] and_355_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] nor_530_nl;
  wire[0:0] nor_531_nl;
  wire[0:0] nor_532_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] nor_533_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] nor_534_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] or_1339_nl;
  wire[0:0] or_1340_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] nand_212_nl;
  wire[0:0] or_1341_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] or_1342_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] or_1345_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] nand_214_nl;
  wire[0:0] mux_612_nl;
  wire[0:0] or_1349_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] nor_128_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] and_349_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] or_538_nl;
  wire[0:0] or_536_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] and_350_nl;
  wire[0:0] mux_633_nl;
  wire[0:0] mux_632_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] or_1330_nl;
  wire[0:0] nand_207_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] nand_208_nl;
  wire[0:0] or_1331_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] mux_656_nl;
  wire[0:0] or_1332_nl;
  wire[0:0] mux_653_nl;
  wire[0:0] nand_210_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] nand_211_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] or_1338_nl;
  wire[0:0] mux_645_nl;
  wire[0:0] nor_135_nl;
  wire[0:0] mux_677_nl;
  wire[0:0] mux_676_nl;
  wire[0:0] mux_675_nl;
  wire[0:0] mux_674_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] and_342_nl;
  wire[0:0] mux_673_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] or_595_nl;
  wire[0:0] or_593_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] and_343_nl;
  wire[0:0] mux_668_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] mux_666_nl;
  wire[0:0] mux_665_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] mux_697_nl;
  wire[0:0] mux_696_nl;
  wire[0:0] mux_695_nl;
  wire[0:0] nand_202_nl;
  wire[0:0] or_1321_nl;
  wire[0:0] mux_694_nl;
  wire[0:0] nand_203_nl;
  wire[0:0] or_1322_nl;
  wire[0:0] mux_693_nl;
  wire[0:0] mux_692_nl;
  wire[0:0] mux_691_nl;
  wire[0:0] nand_204_nl;
  wire[0:0] mux_688_nl;
  wire[0:0] or_1325_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] nand_206_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] or_1329_nl;
  wire[0:0] mux_680_nl;
  wire[0:0] nor_143_nl;
  wire[0:0] mux_712_nl;
  wire[0:0] mux_711_nl;
  wire[0:0] mux_710_nl;
  wire[0:0] mux_709_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] and_334_nl;
  wire[0:0] mux_708_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] mux_707_nl;
  wire[0:0] nor_437_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] mux_706_nl;
  wire[0:0] or_650_nl;
  wire[0:0] or_648_nl;
  wire[0:0] mux_705_nl;
  wire[0:0] mux_704_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] and_335_nl;
  wire[0:0] mux_703_nl;
  wire[0:0] mux_702_nl;
  wire[0:0] nor_440_nl;
  wire[0:0] nor_441_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] mux_701_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] nor_443_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] mux_732_nl;
  wire[0:0] mux_731_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] nand_195_nl;
  wire[0:0] nand_196_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] nand_197_nl;
  wire[0:0] or_1314_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] mux_727_nl;
  wire[0:0] mux_726_nl;
  wire[0:0] nand_198_nl;
  wire[0:0] mux_723_nl;
  wire[0:0] nand_200_nl;
  wire[0:0] mux_720_nl;
  wire[0:0] mux_719_nl;
  wire[0:0] nand_201_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] or_1320_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] and_333_nl;
  wire[0:0] mux_747_nl;
  wire[0:0] mux_746_nl;
  wire[0:0] mux_745_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] and_321_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] and_322_nl;
  wire[0:0] mux_743_nl;
  wire[0:0] and_323_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] mux_742_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] mux_741_nl;
  wire[0:0] or_702_nl;
  wire[0:0] or_700_nl;
  wire[0:0] mux_740_nl;
  wire[0:0] mux_739_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] and_324_nl;
  wire[0:0] mux_738_nl;
  wire[0:0] mux_737_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] mux_736_nl;
  wire[0:0] mux_735_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] mux_734_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] nor_789_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] or_1409_nl;
  wire[0:0] or_1407_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] and_709_nl;
  wire[0:0] and_710_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] and_711_nl;
  wire[0:0] nor_790_nl;
  wire[0:0] and_712_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] nor_791_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] nand_259_nl;
  wire[0:0] or_1403_nl;
  wire[0:0] nor_792_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] nor_784_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] nor_785_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] nand_249_nl;
  wire[0:0] or_1425_nl;
  wire[0:0] and_708_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] and_713_nl;
  wire[0:0] nor_787_nl;
  wire[0:0] nor_788_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] or_1420_nl;
  wire[0:0] nand_247_nl;
  wire[0:0] or_1415_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] or_1456_nl;
  wire[0:0] nand_nl;
  wire[0:0] or_1457_nl;
  wire[0:0] nand_256_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] nor_775_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] nor_777_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] nor_779_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] nor_780_nl;
  wire[0:0] and_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] nor_781_nl;
  wire[0:0] nor_782_nl;
  wire[0:0] nor_783_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] nand_262_nl;
  wire[0:0] or_1442_nl;
  wire[0:0] mux_1038_nl;
  wire[63:0] modExp_while_mux1h_3_nl;
  wire[0:0] and_725_nl;
  wire[0:0] and_726_nl;
  wire[63:0] modExp_while_mux_1_nl;
  wire[0:0] modExp_while_or_2_nl;
  wire[9:0] COMP_LOOP_mux_45_nl;
  wire[0:0] and_727_nl;
  wire[65:0] acc_1_nl;
  wire[66:0] nl_acc_1_nl;
  wire[55:0] COMP_LOOP_COMP_LOOP_or_6_nl;
  wire[55:0] COMP_LOOP_mux_46_nl;
  wire[0:0] COMP_LOOP_mux1h_268_nl;
  wire[0:0] COMP_LOOP_mux1h_269_nl;
  wire[0:0] COMP_LOOP_mux1h_270_nl;
  wire[0:0] COMP_LOOP_mux1h_271_nl;
  wire[0:0] COMP_LOOP_mux1h_272_nl;
  wire[0:0] COMP_LOOP_mux1h_273_nl;
  wire[0:0] COMP_LOOP_mux1h_274_nl;
  wire[0:0] COMP_LOOP_mux1h_275_nl;
  wire[0:0] COMP_LOOP_or_48_nl;
  wire[63:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nand_1_nl;
  wire[63:0] COMP_LOOP_mux_47_nl;
  wire[0:0] COMP_LOOP_not_199_nl;
  wire[8:0] acc_2_nl;
  wire[9:0] nl_acc_2_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_2_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_or_3_nl;
  wire[0:0] operator_64_false_1_mux_1_nl;
  wire[5:0] operator_64_false_1_mux1h_3_nl;
  wire[0:0] operator_64_false_1_or_4_nl;
  wire[0:0] operator_64_false_1_operator_64_false_1_and_1_nl;
  wire[5:0] operator_64_false_1_mux1h_4_nl;
  wire[0:0] operator_64_false_1_or_5_nl;
  wire[10:0] acc_3_nl;
  wire[11:0] nl_acc_3_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_7_nl;
  wire[8:0] COMP_LOOP_COMP_LOOP_mux_9_nl;
  wire[0:0] COMP_LOOP_or_49_nl;
  wire[5:0] COMP_LOOP_COMP_LOOP_mux_10_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_10_nl;
  wire[12:0] COMP_LOOP_acc_58_nl;
  wire[13:0] nl_COMP_LOOP_acc_58_nl;
  wire[9:0] COMP_LOOP_COMP_LOOP_mux_11_nl;
  wire[9:0] COMP_LOOP_acc_59_nl;
  wire[10:0] nl_COMP_LOOP_acc_59_nl;
  wire[2:0] COMP_LOOP_or_50_nl;
  wire[2:0] COMP_LOOP_mux1h_276_nl;
  wire[0:0] and_728_nl;
  wire[0:0] and_729_nl;
  wire[0:0] and_730_nl;
  wire[0:0] and_731_nl;
  wire[0:0] and_732_nl;
  wire[0:0] and_733_nl;
  wire[0:0] and_734_nl;
  wire[0:0] COMP_LOOP_or_51_nl;
  wire[52:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_2_nl;
  wire[0:0] COMP_LOOP_not_200_nl;
  wire[10:0] COMP_LOOP_mux_48_nl;
  wire[5:0] COMP_LOOP_COMP_LOOP_and_220_nl;
  wire[0:0] not_2902_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_11_nl;
  wire[51:0] COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_3_nl;
  wire[0:0] COMP_LOOP_or_52_nl;
  wire[10:0] COMP_LOOP_mux1h_277_nl;
  wire[5:0] COMP_LOOP_COMP_LOOP_and_221_nl;
  wire[0:0] COMP_LOOP_nor_109_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_operator_66_true_div_cmp_b;
  assign nl_operator_66_true_div_cmp_b = {1'b0, operator_66_true_div_cmp_b_9_0};
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 = ~ (z_out_7[64]);
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_65_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_65_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_40_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_130_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_130_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_40_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_195_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_195_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_40_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_260_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_260_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_40_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_325_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_325_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_40_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_390_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_390_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_40_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_455_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_455_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_40_tr0
      = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_1[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 = ~ STAGE_LOOP_acc_itm_2_1;
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_7_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd1)) modulo_result_rem_cmp (
      .a(modulo_result_rem_cmp_a),
      .b(modulo_result_rem_cmp_b),
      .z(modulo_result_rem_cmp_z)
    );
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(nl_operator_66_true_div_cmp_b[10:0]),
      .z(operator_66_true_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_8_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0[0:0]),
      .modExp_while_C_40_tr0(COMP_LOOP_COMP_LOOP_and_11_itm),
      .COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0[0:0]),
      .COMP_LOOP_1_modExp_1_while_C_40_tr0(COMP_LOOP_COMP_LOOP_and_11_itm),
      .COMP_LOOP_C_65_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_65_tr0[0:0]),
      .COMP_LOOP_2_modExp_1_while_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_40_tr0[0:0]),
      .COMP_LOOP_C_130_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_130_tr0[0:0]),
      .COMP_LOOP_3_modExp_1_while_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_40_tr0[0:0]),
      .COMP_LOOP_C_195_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_195_tr0[0:0]),
      .COMP_LOOP_4_modExp_1_while_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_40_tr0[0:0]),
      .COMP_LOOP_C_260_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_260_tr0[0:0]),
      .COMP_LOOP_5_modExp_1_while_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_40_tr0[0:0]),
      .COMP_LOOP_C_325_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_325_tr0[0:0]),
      .COMP_LOOP_6_modExp_1_while_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_40_tr0[0:0]),
      .COMP_LOOP_C_390_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_390_tr0[0:0]),
      .COMP_LOOP_7_modExp_1_while_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_40_tr0[0:0]),
      .COMP_LOOP_C_455_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_455_tr0[0:0]),
      .COMP_LOOP_8_modExp_1_while_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_40_tr0[0:0]),
      .COMP_LOOP_C_520_tr0(COMP_LOOP_COMP_LOOP_and_2_itm),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_9_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0[0:0])
    );
  assign or_1380_nl = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[5]) | nand_245_cse;
  assign or_1381_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[5])
      | (fsm_output[9]) | (~ (fsm_output[7]));
  assign mux_477_cse = MUX_s_1_2_2(or_1380_nl, or_1381_nl, fsm_output[4]);
  assign or_294_cse = (COMP_LOOP_acc_13_psp_sva[0]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]);
  assign nor_624_cse = ~((fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[6:5]!=2'b10)
      | not_tmp_170);
  assign nor_594_cse = ~((fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[6:5]!=2'b10)
      | not_tmp_170);
  assign nor_115_cse = ~((COMP_LOOP_acc_13_psp_sva[0]) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (VEC_LOOP_j_sva_11_0[1])));
  assign or_521_cse = (~ (COMP_LOOP_acc_13_psp_sva[0])) | (~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (VEC_LOOP_j_sva_11_0[1]);
  assign and_336_cse = (COMP_LOOP_acc_13_psp_sva[0]) & COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm
      & (VEC_LOOP_j_sva_11_0[1]);
  assign and_316_cse = (fsm_output[2:1]==2'b11);
  assign or_722_cse = (fsm_output[2:1]!=2'b00);
  assign or_730_cse = (fsm_output[0]) | (fsm_output[7]);
  assign nor_397_cse = ~((fsm_output[6]) | (fsm_output[9]) | (~ (fsm_output[1]))
      | (~ (fsm_output[3])) | (fsm_output[5]));
  assign nor_398_cse = ~((fsm_output[9:1]!=9'b000011010));
  assign nor_400_cse = ~((~ (fsm_output[7])) | (fsm_output[0]));
  assign nor_401_cse = ~((fsm_output[0]) | (fsm_output[9]));
  assign and_312_cse = (fsm_output[7]) & (fsm_output[9]);
  assign or_1275_cse = (~ (fsm_output[0])) | (fsm_output[9]);
  assign or_731_cse = (~ (fsm_output[6])) | (fsm_output[8]);
  assign or_718_cse = (fsm_output[8]) | (fsm_output[0]) | (~ (fsm_output[7]));
  assign and_303_cse = (fsm_output[1:0]==2'b11);
  assign nor_379_cse = ~((fsm_output[0]) | (fsm_output[4]));
  assign or_217_cse = (fsm_output[6:3]!=4'b0000);
  assign and_56_nl = (fsm_output[7]) & or_217_cse;
  assign and_55_nl = (fsm_output[7]) & or_5_cse;
  assign mux_445_cse = MUX_s_1_2_2(and_56_nl, and_55_nl, fsm_output[1]);
  assign and_57_nl = (fsm_output[8]) & mux_445_cse;
  assign mux_446_cse = MUX_s_1_2_2(not_tmp_129, and_57_nl, fsm_output[9]);
  assign or_831_cse = (fsm_output[9:8]!=2'b01);
  assign mux_995_cse = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[8]);
  assign mux_1001_cse = MUX_s_1_2_2(mux_tmp_898, or_tmp_71, fsm_output[0]);
  assign nor_333_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[3])) | (fsm_output[5]));
  assign mux_1107_nl = MUX_s_1_2_2(nor_333_nl, nor_397_cse, fsm_output[8]);
  assign nor_335_nl = ~((fsm_output[8]) | (fsm_output[6]) | (fsm_output[9]) | (fsm_output[1])
      | (fsm_output[3]) | (~ (fsm_output[5])));
  assign mux_1108_nl = MUX_s_1_2_2(mux_1107_nl, nor_335_nl, fsm_output[7]);
  assign nor_336_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (fsm_output[6]) |
      (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[3]) | (~ (fsm_output[5])));
  assign mux_1109_nl = MUX_s_1_2_2(mux_1108_nl, nor_336_nl, fsm_output[4]);
  assign nor_337_nl = ~((~ (fsm_output[9])) | (fsm_output[1]) | (~ (fsm_output[3]))
      | (fsm_output[5]));
  assign nor_338_nl = ~((fsm_output[9]) | (fsm_output[1]) | (fsm_output[3]) | (~
      (fsm_output[5])));
  assign mux_1105_nl = MUX_s_1_2_2(nor_337_nl, nor_338_nl, fsm_output[6]);
  assign and_275_nl = (fsm_output[8]) & mux_1105_nl;
  assign nor_339_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (~ (fsm_output[3])) | (fsm_output[5]));
  assign mux_1106_nl = MUX_s_1_2_2(and_275_nl, nor_339_nl, fsm_output[7]);
  assign and_274_nl = (fsm_output[4]) & mux_1106_nl;
  assign mux_1110_nl = MUX_s_1_2_2(mux_1109_nl, and_274_nl, fsm_output[2]);
  assign mux_1111_nl = MUX_s_1_2_2(mux_1110_nl, nor_398_cse, fsm_output[0]);
  assign modExp_while_if_or_nl = and_dcpl_150 | (mux_1111_nl & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign modExp_1_while_and_16_nl = (~ (modulo_result_rem_cmp_z[63])) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & and_dcpl_174;
  assign modExp_1_while_and_18_nl = (modulo_result_rem_cmp_z[63]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & and_dcpl_174;
  assign modExp_while_if_mux1h_nl = MUX1HOT_v_64_5_2(z_out, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      modulo_result_rem_cmp_z, modulo_qr_sva_1_mx1w1, COMP_LOOP_1_acc_5_mut_mx0w5,
      {modExp_while_if_or_nl , COMP_LOOP_nor_97_cse , modExp_1_while_and_16_nl ,
      modExp_1_while_and_18_nl , and_dcpl_151});
  assign mux_949_nl = MUX_s_1_2_2((~ or_tmp_71), mux_tmp_898, or_731_cse);
  assign mux_1005_nl = MUX_s_1_2_2(mux_923_cse, mux_tmp_900, fsm_output[6]);
  assign mux_950_nl = MUX_s_1_2_2(mux_949_nl, mux_1005_nl, fsm_output[1]);
  assign mux_1002_nl = MUX_s_1_2_2((~ or_tmp_71), mux_1001_cse, fsm_output[8]);
  assign mux_1003_nl = MUX_s_1_2_2(mux_919_cse, mux_1002_nl, fsm_output[6]);
  assign mux_1000_nl = MUX_s_1_2_2(mux_937_cse, (fsm_output[8]), fsm_output[6]);
  assign mux_1004_nl = MUX_s_1_2_2(mux_1003_nl, mux_1000_nl, fsm_output[1]);
  assign mux_951_nl = MUX_s_1_2_2(mux_950_nl, mux_1004_nl, fsm_output[2]);
  assign mux_952_nl = MUX_s_1_2_2(mux_951_nl, mux_1460_cse, fsm_output[5]);
  assign mux_996_nl = MUX_s_1_2_2(mux_995_cse, mux_937_cse, fsm_output[6]);
  assign mux_991_nl = MUX_s_1_2_2((~ (fsm_output[7])), and_312_cse, fsm_output[8]);
  assign mux_992_nl = MUX_s_1_2_2(mux_991_nl, mux_929_cse, fsm_output[6]);
  assign mux_997_nl = MUX_s_1_2_2(mux_996_nl, mux_992_nl, fsm_output[1]);
  assign mux_998_nl = MUX_s_1_2_2(mux_997_nl, mux_1447_cse, fsm_output[2]);
  assign mux_999_nl = MUX_s_1_2_2(mux_928_cse, mux_998_nl, fsm_output[5]);
  assign mux_953_nl = MUX_s_1_2_2(mux_952_nl, mux_999_nl, fsm_output[4]);
  assign and_176_nl = (fsm_output[8]) & or_tmp_783;
  assign mux_987_nl = MUX_s_1_2_2(mux_929_cse, and_176_nl, fsm_output[6]);
  assign mux_988_nl = MUX_s_1_2_2(mux_987_nl, mux_928_cse, or_722_cse);
  assign mux_981_nl = MUX_s_1_2_2(mux_903_cse, mux_923_cse, fsm_output[6]);
  assign mux_977_nl = MUX_s_1_2_2(mux_tmp_898, or_tmp_72, fsm_output[0]);
  assign mux_978_nl = MUX_s_1_2_2(mux_977_nl, (fsm_output[7]), fsm_output[8]);
  assign mux_979_nl = MUX_s_1_2_2(mux_978_nl, mux_919_cse, fsm_output[6]);
  assign mux_982_nl = MUX_s_1_2_2(mux_981_nl, mux_979_nl, fsm_output[1]);
  assign mux_984_nl = MUX_s_1_2_2(mux_1460_cse, mux_982_nl, fsm_output[2]);
  assign mux_989_nl = MUX_s_1_2_2(mux_988_nl, mux_984_nl, fsm_output[5]);
  assign mux_970_nl = MUX_s_1_2_2((~ mux_tmp_898), or_tmp_783, fsm_output[0]);
  assign mux_971_nl = MUX_s_1_2_2(mux_970_nl, (fsm_output[9]), fsm_output[8]);
  assign mux_972_nl = MUX_s_1_2_2(mux_971_nl, mux_tmp_912, fsm_output[6]);
  assign mux_967_nl = MUX_s_1_2_2(or_tmp_783, and_312_cse, fsm_output[8]);
  assign mux_966_nl = MUX_s_1_2_2((~ or_tmp_72), or_823_cse, fsm_output[8]);
  assign mux_968_nl = MUX_s_1_2_2(mux_967_nl, mux_966_nl, fsm_output[6]);
  assign mux_973_nl = MUX_s_1_2_2(mux_972_nl, mux_968_nl, fsm_output[1]);
  assign mux_963_nl = MUX_s_1_2_2(or_823_cse, and_312_cse, fsm_output[8]);
  assign mux_962_nl = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_831_cse);
  assign mux_964_nl = MUX_s_1_2_2(mux_963_nl, mux_962_nl, fsm_output[6]);
  assign mux_959_nl = MUX_s_1_2_2(and_312_cse, mux_tmp_898, fsm_output[8]);
  assign mux_961_nl = MUX_s_1_2_2(mux_903_cse, mux_959_nl, fsm_output[6]);
  assign mux_965_nl = MUX_s_1_2_2(mux_964_nl, mux_961_nl, fsm_output[1]);
  assign mux_974_nl = MUX_s_1_2_2(mux_973_nl, mux_965_nl, fsm_output[2]);
  assign mux_975_nl = MUX_s_1_2_2(mux_974_nl, mux_1447_cse, fsm_output[5]);
  assign mux_990_nl = MUX_s_1_2_2(mux_989_nl, mux_975_nl, fsm_output[4]);
  assign mux_954_nl = MUX_s_1_2_2(mux_953_nl, mux_990_nl, fsm_output[3]);
  assign operator_64_false_operator_64_false_mux_rgt = MUX_v_65_2_2(({1'b0 , modExp_while_if_mux1h_nl}),
      z_out_2, mux_954_nl);
  assign or_1470_cse = (fsm_output[1:0]!=2'b00);
  assign or_1516_cse = (fsm_output[3:2]!=2'b00);
  assign and_721_cse = (fsm_output[3:2]==2'b11);
  assign nor_813_cse = ~((fsm_output[6]) | (~ (fsm_output[8])));
  assign or_1466_nl = nor_813_cse | (fsm_output[9]);
  assign mux_1460_cse = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_1466_nl);
  assign mux_1447_cse = MUX_s_1_2_2(mux_tmp_900, mux_tmp_899, fsm_output[6]);
  assign or_1483_cse = (fsm_output[9:8]!=2'b00);
  assign nor_820_cse = ~(COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm | (~ (fsm_output[8])));
  assign or_843_cse = (~ (fsm_output[3])) | (fsm_output[1]) | (fsm_output[4]) | (fsm_output[5]);
  assign or_857_cse = (fsm_output[7:6]!=2'b00);
  assign and_293_cse = (fsm_output[7:6]==2'b11);
  assign and_292_cse = (fsm_output[5:4]==2'b11);
  assign or_844_nl = (fsm_output[3]) | (~((fsm_output[1]) & (fsm_output[4]) & (fsm_output[5])));
  assign mux_1014_cse = MUX_s_1_2_2(or_844_nl, or_843_cse, fsm_output[0]);
  assign and_185_m1c = and_dcpl_103 & and_dcpl_72;
  assign or_5_cse = (fsm_output[6:2]!=5'b00000);
  assign modExp_result_and_rgt = (~ modExp_while_and_1_rgt) & and_185_m1c;
  assign modExp_result_and_1_rgt = modExp_while_and_1_rgt & and_185_m1c;
  assign COMP_LOOP_COMP_LOOP_and_11_cse = (z_out_6_12_1[2:0]==3'b101);
  assign modExp_while_or_1_cse = and_dcpl_90 | and_dcpl_98 | and_dcpl_104 | and_dcpl_109
      | and_dcpl_116 | and_dcpl_126 | and_dcpl_134;
  assign COMP_LOOP_COMP_LOOP_and_37_cse = (z_out_6_12_1[2:0]==3'b011);
  assign nor_692_cse = ~((fsm_output[9:7]!=3'b000));
  assign or_157_cse = (fsm_output[4:3]!=2'b00);
  assign and_398_cse = (fsm_output[4:3]==2'b11);
  assign nor_308_nl = ~((fsm_output[4]) | (fsm_output[3]) | (~ (fsm_output[7])) |
      (fsm_output[5]));
  assign nor_309_nl = ~((fsm_output[4]) | (~ (fsm_output[3])) | (fsm_output[7]) |
      (~ (fsm_output[5])));
  assign mux_1257_nl = MUX_s_1_2_2(nor_308_nl, nor_309_nl, fsm_output[9]);
  assign nand_82_cse = ~((fsm_output[6]) & mux_1257_nl);
  assign or_1161_cse = (fsm_output[1]) | (fsm_output[6]) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[2]) | (fsm_output[7]);
  assign or_1156_cse = (~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[7]);
  assign or_1168_nl = (fsm_output[4]) | (~ (fsm_output[1])) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[2])) | (fsm_output[7]);
  assign or_1166_nl = (fsm_output[8]) | (~ (fsm_output[2])) | (fsm_output[7]);
  assign or_1165_nl = (fsm_output[8]) | (fsm_output[2]) | (~ (fsm_output[7]));
  assign mux_1318_nl = MUX_s_1_2_2(or_1166_nl, or_1165_nl, fsm_output[9]);
  assign nor_292_nl = ~((fsm_output[6]) | mux_1318_nl);
  assign nor_293_nl = ~((~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[2]) | (fsm_output[7]));
  assign mux_1319_nl = MUX_s_1_2_2(nor_292_nl, nor_293_nl, fsm_output[1]);
  assign nand_86_nl = ~((fsm_output[4]) & mux_1319_nl);
  assign mux_1320_nl = MUX_s_1_2_2(or_1168_nl, nand_86_nl, fsm_output[5]);
  assign or_1160_nl = (~ (fsm_output[6])) | (fsm_output[9]) | (~((fsm_output[8])
      & (fsm_output[2]) & (fsm_output[7])));
  assign or_1157_nl = (fsm_output[8]) | (~((fsm_output[2]) & (fsm_output[7])));
  assign mux_1315_nl = MUX_s_1_2_2(or_1157_nl, or_1156_cse, fsm_output[9]);
  assign or_1158_nl = (fsm_output[6]) | mux_1315_nl;
  assign mux_1316_nl = MUX_s_1_2_2(or_1160_nl, or_1158_nl, fsm_output[1]);
  assign mux_1317_nl = MUX_s_1_2_2(or_1161_cse, mux_1316_nl, fsm_output[4]);
  assign or_1162_nl = (fsm_output[5]) | mux_1317_nl;
  assign mux_1321_nl = MUX_s_1_2_2(mux_1320_nl, or_1162_nl, fsm_output[3]);
  assign COMP_LOOP_nor_97_cse = ~(mux_1321_nl | (fsm_output[0]));
  assign modulo_result_mux_1_cse = MUX_v_64_2_2(modulo_result_rem_cmp_z, modulo_qr_sva_1_mx1w1,
      modulo_result_rem_cmp_z[63]);
  assign nand_245_cse = ~((fsm_output[7]) & (fsm_output[9]));
  assign or_29_cse = (fsm_output[7]) | (~ (fsm_output[1])) | (~ (fsm_output[9]))
      | (fsm_output[6]) | (~ (fsm_output[8]));
  assign nand_244_cse = ~(nand_245_cse & (fsm_output[8]));
  assign mux_417_cse = MUX_s_1_2_2(not_tmp_121, or_1483_cse, fsm_output[7]);
  assign mux_438_cse = MUX_s_1_2_2(or_tmp_73, mux_tmp_390, fsm_output[6]);
  assign nor_265_cse = ~((fsm_output[2]) | (~ (fsm_output[4])));
  assign COMP_LOOP_or_3_cse = and_dcpl_77 | and_dcpl_90 | and_dcpl_98 | and_dcpl_104
      | and_dcpl_109 | and_dcpl_116 | and_dcpl_126 | and_dcpl_134;
  assign COMP_LOOP_COMP_LOOP_and_12_cse = (z_out_6_12_1[2:0]==3'b110);
  assign COMP_LOOP_COMP_LOOP_and_13_cse = (z_out_6_12_1[2:0]==3'b111);
  assign nl_STAGE_LOOP_i_3_0_sva_2 = STAGE_LOOP_i_3_0_sva + 4'b0001;
  assign STAGE_LOOP_i_3_0_sva_2 = nl_STAGE_LOOP_i_3_0_sva_2[3:0];
  assign nl_COMP_LOOP_acc_psp_sva_1 = (VEC_LOOP_j_sva_11_0[11:3]) + conv_u2u_6_9(COMP_LOOP_k_9_3_sva_5_0);
  assign COMP_LOOP_acc_psp_sva_1 = nl_COMP_LOOP_acc_psp_sva_1[8:0];
  assign nl_COMP_LOOP_1_acc_5_mut_mx0w5 = tmp_10_lpi_4_dfm + modulo_result_mux_1_cse;
  assign COMP_LOOP_1_acc_5_mut_mx0w5 = nl_COMP_LOOP_1_acc_5_mut_mx0w5[63:0];
  assign modExp_while_and_1_rgt = (modulo_result_rem_cmp_z[63]) & operator_64_false_slc_modExp_exp_0_1_itm;
  assign nl_modulo_qr_sva_1_mx1w1 = modulo_result_rem_cmp_z + p_sva;
  assign modulo_qr_sva_1_mx1w1 = nl_modulo_qr_sva_1_mx1w1[63:0];
  assign operator_64_false_slc_modExp_exp_63_1_3 = MUX_v_63_2_2((operator_66_true_div_cmp_z[63:1]),
      ({1'b0 , (modExp_exp_sva_rsp_1[62:1])}), or_dcpl_56);
  assign nl_COMP_LOOP_acc_1_cse_2_sva_1 = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_3_sva_5_0
      , 3'b001});
  assign COMP_LOOP_acc_1_cse_2_sva_1 = nl_COMP_LOOP_acc_1_cse_2_sva_1[11:0];
  assign COMP_LOOP_COMP_LOOP_and_211 = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b001);
  assign COMP_LOOP_COMP_LOOP_and_213 = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b010);
  assign COMP_LOOP_COMP_LOOP_and_215 = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b100);
  assign or_dcpl_3 = (~ COMP_LOOP_COMP_LOOP_and_11_itm) | (z_out_7[64]);
  assign or_tmp_5 = (fsm_output[7:6]!=2'b01);
  assign or_tmp_9 = (~ (fsm_output[0])) | (fsm_output[7]);
  assign or_tmp_13 = (fsm_output[7:6]!=2'b10);
  assign nand_240_cse = ~((fsm_output[6]) & (fsm_output[0]));
  assign not_tmp_29 = ~((fsm_output[6]) & (fsm_output[8]));
  assign or_tmp_58 = (fsm_output[5]) | and_398_cse;
  assign or_tmp_60 = (fsm_output[5:2]!=4'b0000);
  assign mux_tmp_77 = MUX_s_1_2_2((~ and_292_cse), or_tmp_58, fsm_output[6]);
  assign or_tmp_63 = and_721_cse | (fsm_output[4]);
  assign not_tmp_46 = ~((fsm_output[4:3]!=2'b00));
  assign mux_tmp_81 = MUX_s_1_2_2(not_tmp_46, (fsm_output[4]), fsm_output[5]);
  assign mux_82_cse = MUX_s_1_2_2(or_tmp_60, mux_tmp_81, fsm_output[6]);
  assign mux_tmp_83 = MUX_s_1_2_2(mux_82_cse, mux_tmp_77, fsm_output[7]);
  assign nor_tmp_12 = or_1516_cse & (fsm_output[4]);
  assign and_tmp_2 = (fsm_output[5]) & nor_tmp_12;
  assign or_tmp_71 = (~ (fsm_output[9])) | (fsm_output[7]);
  assign or_tmp_72 = (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_tmp_73 = (fsm_output[9:8]!=2'b10);
  assign or_90_cse = (fsm_output[8:7]!=2'b10);
  assign or_91_cse = (fsm_output[8:7]!=2'b01);
  assign nor_tmp_13 = (fsm_output[8:7]==2'b11);
  assign mux_tmp_164 = MUX_s_1_2_2(or_90_cse, or_91_cse, fsm_output[6]);
  assign and_434_cse = (fsm_output[9]) & (fsm_output[6]);
  assign and_433_cse = (fsm_output[6:4]==3'b111);
  assign nor_tmp_21 = (fsm_output[9:7]==3'b111);
  assign not_tmp_82 = ~((fsm_output[9:8]!=2'b00));
  assign and_432_nl = (fsm_output[9:8]==2'b11);
  assign mux_tmp_229 = MUX_s_1_2_2(not_tmp_82, and_432_nl, fsm_output[7]);
  assign or_119_cse = (fsm_output[6]) | (fsm_output[9]);
  assign mux_tmp_390 = MUX_s_1_2_2((~ (fsm_output[8])), or_1483_cse, fsm_output[7]);
  assign not_tmp_121 = ~((fsm_output[9:8]==2'b11));
  assign and_dcpl_15 = ~((fsm_output[7]) | (fsm_output[1]));
  assign and_dcpl_16 = and_dcpl_15 & (fsm_output[8]);
  assign and_dcpl_18 = (fsm_output[6:5]==2'b10);
  assign and_dcpl_23 = not_tmp_46 & (fsm_output[2]);
  assign and_dcpl_26 = (fsm_output[9]) & (~ (fsm_output[0]));
  assign and_dcpl_33 = ~((fsm_output[6:5]!=2'b00));
  assign not_tmp_129 = ~((fsm_output[8:1]!=8'b00000000));
  assign and_60_nl = (fsm_output[9:8]==2'b11) & mux_445_cse;
  assign mux_453_itm = MUX_s_1_2_2(mux_446_cse, and_60_nl, fsm_output[0]);
  assign and_dcpl_49 = and_dcpl_15 & (~ (fsm_output[8]));
  assign and_dcpl_50 = and_dcpl_49 & nor_401_cse;
  assign and_dcpl_53 = not_tmp_46 & (~ (fsm_output[2]));
  assign and_dcpl_57 = (fsm_output[7]) & (~ (fsm_output[1]));
  assign and_dcpl_58 = and_dcpl_57 & (fsm_output[8]);
  assign and_dcpl_61 = and_dcpl_23 & and_dcpl_33;
  assign or_dcpl_39 = or_157_cse | (fsm_output[5]);
  assign and_dcpl_63 = (~ (fsm_output[9])) & (fsm_output[0]);
  assign and_dcpl_64 = (~ (fsm_output[7])) & (fsm_output[1]);
  assign and_dcpl_65 = and_dcpl_64 & (~ (fsm_output[8]));
  assign and_dcpl_66 = and_dcpl_65 & and_dcpl_63;
  assign and_dcpl_67 = (fsm_output[6:5]==2'b01);
  assign and_dcpl_68 = (fsm_output[4:3]==2'b10);
  assign and_dcpl_69 = and_dcpl_68 & (~ (fsm_output[2]));
  assign and_dcpl_70 = and_dcpl_69 & and_dcpl_67;
  assign and_dcpl_71 = and_dcpl_70 & and_dcpl_66;
  assign and_dcpl_72 = and_dcpl_65 & nor_401_cse;
  assign and_dcpl_75 = and_398_cse & (fsm_output[2]);
  assign and_dcpl_76 = and_dcpl_75 & and_dcpl_18;
  assign and_dcpl_77 = and_dcpl_76 & and_dcpl_72;
  assign and_dcpl_78 = and_dcpl_57 & (~ (fsm_output[8]));
  assign and_dcpl_79 = and_dcpl_78 & nor_401_cse;
  assign and_dcpl_81 = (fsm_output[4:2]==3'b010);
  assign and_dcpl_82 = and_dcpl_81 & and_dcpl_33;
  assign and_dcpl_90 = and_dcpl_81 & and_dcpl_18 & and_dcpl_79;
  assign and_dcpl_91 = (fsm_output[9:8]==2'b01);
  assign and_dcpl_96 = and_dcpl_64 & (fsm_output[8]);
  assign and_dcpl_97 = and_dcpl_96 & nor_401_cse;
  assign and_dcpl_98 = and_dcpl_70 & and_dcpl_97;
  assign and_dcpl_102 = and_dcpl_58 & nor_401_cse;
  assign and_dcpl_103 = and_dcpl_75 & and_dcpl_33;
  assign and_dcpl_104 = and_dcpl_103 & and_dcpl_102;
  assign and_dcpl_108 = and_dcpl_65 & and_dcpl_26;
  assign and_dcpl_109 = and_dcpl_61 & and_dcpl_108;
  assign and_dcpl_115 = and_dcpl_69 & (fsm_output[6:5]==2'b11);
  assign and_dcpl_116 = and_dcpl_115 & and_dcpl_49 & and_dcpl_26;
  assign and_dcpl_122 = (fsm_output[7]) & (fsm_output[1]) & (~ (fsm_output[8]));
  assign and_dcpl_124 = and_398_cse & (~ (fsm_output[2]));
  assign and_dcpl_126 = and_dcpl_124 & and_dcpl_18 & and_dcpl_122 & and_dcpl_26;
  assign and_dcpl_133 = and_dcpl_23 & and_dcpl_18;
  assign and_dcpl_134 = and_dcpl_133 & and_dcpl_16 & and_dcpl_26;
  assign or_263_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b000) | (fsm_output[5]) |
      (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_261_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b000) | (~ (fsm_output[5]))
      | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_469 = MUX_s_1_2_2(or_263_nl, or_261_nl, fsm_output[3]);
  assign nor_640_nl = ~((~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b000)
      | (fsm_output[5]) | nand_245_cse);
  assign nor_641_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b000)
      | (fsm_output[9]) | (~ (fsm_output[7])));
  assign not_tmp_166 = MUX_s_1_2_2(nor_640_nl, nor_641_nl, fsm_output[6]);
  assign or_270_nl = (fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00)
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[7]);
  assign or_269_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00)
      | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]);
  assign mux_tmp_472 = MUX_s_1_2_2(or_270_nl, or_269_nl, fsm_output[4]);
  assign or_275_nl = (VEC_LOOP_j_sva_11_0[2]) | (fsm_output[6]) | (~ (fsm_output[3]))
      | (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_273_nl = (fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_13_psp_sva[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_473 = MUX_s_1_2_2(or_275_nl, or_273_nl, fsm_output[4]);
  assign or_1376_nl = (~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[5]) | (~
      (fsm_output[9])) | (fsm_output[7]);
  assign or_1377_nl = (fsm_output[6]) | (~ (fsm_output[3])) | (fsm_output[5]) | (fsm_output[9])
      | (~ (fsm_output[7]));
  assign mux_483_cse = MUX_s_1_2_2(or_1376_nl, or_1377_nl, fsm_output[4]);
  assign nor_630_nl = ~((~ (fsm_output[3])) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (fsm_output[7]));
  assign nor_631_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[9]) |
      (fsm_output[7]));
  assign mux_481_nl = MUX_s_1_2_2(nor_630_nl, nor_631_nl, fsm_output[6]);
  assign nand_232_cse = ~((fsm_output[4]) & mux_481_nl);
  assign or_1379_cse = (fsm_output[4]) | (fsm_output[6]) | (~((fsm_output[3]) & (fsm_output[5])
      & (fsm_output[9]) & (fsm_output[7])));
  assign or_277_cse = (fsm_output[3]) | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]);
  assign or_297_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b000) | (fsm_output[7:3]!=5'b01110);
  assign or_296_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b000) | (fsm_output[7:3]!=5'b00011);
  assign mux_tmp_488 = MUX_s_1_2_2(or_297_nl, or_296_nl, fsm_output[9]);
  assign not_tmp_170 = ~((fsm_output[4]) & (fsm_output[3]) & (fsm_output[7]));
  assign not_tmp_171 = ~((fsm_output[3]) & (fsm_output[7]));
  assign or_324_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b001) | (fsm_output[5]) |
      (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_322_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b001) | (~ (fsm_output[5]))
      | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_504 = MUX_s_1_2_2(or_324_nl, or_322_nl, fsm_output[3]);
  assign nor_610_nl = ~((~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b001)
      | (fsm_output[5]) | nand_245_cse);
  assign nor_611_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b001)
      | (fsm_output[9]) | (~ (fsm_output[7])));
  assign not_tmp_177 = MUX_s_1_2_2(nor_610_nl, nor_611_nl, fsm_output[6]);
  assign nor_608_nl = ~((fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00)
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[7]));
  assign nor_609_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00)
      | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]));
  assign not_tmp_178 = MUX_s_1_2_2(nor_608_nl, nor_609_nl, fsm_output[4]);
  assign or_355_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b001) | (fsm_output[7:3]!=5'b01110);
  assign or_354_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b001) | (fsm_output[7:3]!=5'b00011);
  assign mux_tmp_523 = MUX_s_1_2_2(or_355_nl, or_354_nl, fsm_output[9]);
  assign or_382_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b010) | (fsm_output[5]) |
      (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_380_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b010) | (~ (fsm_output[5]))
      | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_539 = MUX_s_1_2_2(or_382_nl, or_380_nl, fsm_output[3]);
  assign nor_580_nl = ~((~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b010)
      | (fsm_output[5]) | nand_245_cse);
  assign nor_581_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b010)
      | (fsm_output[9]) | (~ (fsm_output[7])));
  assign not_tmp_189 = MUX_s_1_2_2(nor_580_nl, nor_581_nl, fsm_output[6]);
  assign or_389_nl = (fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01)
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[7]);
  assign or_388_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01)
      | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]);
  assign mux_tmp_542 = MUX_s_1_2_2(or_389_nl, or_388_nl, fsm_output[4]);
  assign nor_578_nl = ~((VEC_LOOP_j_sva_11_0[2]) | (fsm_output[6]) | (~ (fsm_output[3]))
      | (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[7])));
  assign nor_579_nl = ~((fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_13_psp_sva[0])
      | (~ (fsm_output[5])) | (~ (fsm_output[9])) | (fsm_output[7]));
  assign not_tmp_190 = MUX_s_1_2_2(nor_578_nl, nor_579_nl, fsm_output[4]);
  assign nor_112_cse = ~((fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10));
  assign nor_114_cse = ~((VEC_LOOP_j_sva_11_0[1:0]!=2'b10));
  assign or_412_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b010) | (fsm_output[7:3]!=5'b01110);
  assign or_411_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b010) | (fsm_output[7:3]!=5'b00011);
  assign mux_tmp_558 = MUX_s_1_2_2(or_412_nl, or_411_nl, fsm_output[9]);
  assign or_438_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b011) | (fsm_output[5]) |
      (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_436_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b011) | (~ (fsm_output[5]))
      | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_574 = MUX_s_1_2_2(or_438_nl, or_436_nl, fsm_output[3]);
  assign nor_550_nl = ~((~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b011)
      | (fsm_output[5]) | nand_245_cse);
  assign nor_551_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b011)
      | (fsm_output[9]) | (~ (fsm_output[7])));
  assign not_tmp_201 = MUX_s_1_2_2(nor_550_nl, nor_551_nl, fsm_output[6]);
  assign nor_548_nl = ~((fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01)
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[7]));
  assign nor_549_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01)
      | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]));
  assign not_tmp_202 = MUX_s_1_2_2(nor_548_nl, nor_549_nl, fsm_output[4]);
  assign nor_122_cse = ~((fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11));
  assign or_465_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b011) | (fsm_output[7:3]!=5'b01110);
  assign or_464_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b011) | (fsm_output[7:3]!=5'b00011);
  assign mux_tmp_593 = MUX_s_1_2_2(or_465_nl, or_464_nl, fsm_output[9]);
  assign or_490_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b100) | (fsm_output[5]) |
      (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_488_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b100) | (~ (fsm_output[5]))
      | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_609 = MUX_s_1_2_2(or_490_nl, or_488_nl, fsm_output[3]);
  assign nor_520_nl = ~((~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b100)
      | (fsm_output[5]) | nand_245_cse);
  assign nor_521_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b100)
      | (fsm_output[9]) | (~ (fsm_output[7])));
  assign not_tmp_214 = MUX_s_1_2_2(nor_520_nl, nor_521_nl, fsm_output[6]);
  assign or_504_nl = (fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10)
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[7]);
  assign or_503_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10)
      | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]);
  assign mux_tmp_616 = MUX_s_1_2_2(or_504_nl, or_503_nl, fsm_output[4]);
  assign or_514_nl = (~ (VEC_LOOP_j_sva_11_0[2])) | (fsm_output[6]) | (~ (fsm_output[3]))
      | (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_512_nl = (fsm_output[6]) | (fsm_output[3]) | (~ (COMP_LOOP_acc_13_psp_sva[0]))
      | (~ (fsm_output[5])) | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_620 = MUX_s_1_2_2(or_514_nl, or_512_nl, fsm_output[4]);
  assign or_524_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b100) | (fsm_output[7:3]!=5'b01110);
  assign or_523_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b100) | (fsm_output[7:3]!=5'b00011);
  assign mux_tmp_628 = MUX_s_1_2_2(or_524_nl, or_523_nl, fsm_output[9]);
  assign or_550_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b101) | (fsm_output[5]) |
      (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_548_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b101) | (~ (fsm_output[5]))
      | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_644 = MUX_s_1_2_2(or_550_nl, or_548_nl, fsm_output[3]);
  assign nor_490_nl = ~((~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b101)
      | (fsm_output[5]) | nand_245_cse);
  assign nor_491_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b101)
      | (fsm_output[9]) | (~ (fsm_output[7])));
  assign not_tmp_225 = MUX_s_1_2_2(nor_490_nl, nor_491_nl, fsm_output[6]);
  assign nor_488_nl = ~((fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10)
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[7]));
  assign nor_489_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10)
      | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]));
  assign not_tmp_226 = MUX_s_1_2_2(nor_488_nl, nor_489_nl, fsm_output[4]);
  assign or_581_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b101) | (fsm_output[7:3]!=5'b01110);
  assign or_580_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b101) | (fsm_output[7:3]!=5'b00011);
  assign mux_tmp_663 = MUX_s_1_2_2(or_581_nl, or_580_nl, fsm_output[9]);
  assign or_607_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b110) | (fsm_output[5]) |
      (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_605_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b110) | (~ (fsm_output[5]))
      | (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_tmp_679 = MUX_s_1_2_2(or_607_nl, or_605_nl, fsm_output[3]);
  assign nor_460_nl = ~((~ (fsm_output[3])) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b110)
      | (fsm_output[5]) | nand_245_cse);
  assign nor_461_nl = ~((fsm_output[3]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b110)
      | (fsm_output[9]) | (~ (fsm_output[7])));
  assign not_tmp_237 = MUX_s_1_2_2(nor_460_nl, nor_461_nl, fsm_output[6]);
  assign or_621_nl = (fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b11)
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[7]);
  assign or_620_nl = (~ (fsm_output[6])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b11)
      | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]);
  assign mux_tmp_686 = MUX_s_1_2_2(or_621_nl, or_620_nl, fsm_output[4]);
  assign nor_458_nl = ~((~ (VEC_LOOP_j_sva_11_0[2])) | (fsm_output[6]) | (~ (fsm_output[3]))
      | (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[7])));
  assign nor_459_nl = ~((fsm_output[6]) | (fsm_output[3]) | (~ (COMP_LOOP_acc_13_psp_sva[0]))
      | (~ (fsm_output[5])) | (~ (fsm_output[9])) | (fsm_output[7]));
  assign not_tmp_239 = MUX_s_1_2_2(nor_458_nl, nor_459_nl, fsm_output[4]);
  assign or_637_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b110) | (fsm_output[7:3]!=5'b01110);
  assign or_636_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b110) | (fsm_output[7:3]!=5'b00011);
  assign mux_tmp_698 = MUX_s_1_2_2(or_637_nl, or_636_nl, fsm_output[9]);
  assign or_662_nl = (COMP_LOOP_acc_1_cse_4_sva[2:0]!=3'b111) | (fsm_output[5]) |
      (fsm_output[9]) | (~ (fsm_output[7]));
  assign nand_136_nl = ~((COMP_LOOP_acc_1_cse_sva[2:0]==3'b111) & (fsm_output[5])
      & (fsm_output[9]) & (~ (fsm_output[7])));
  assign mux_tmp_714 = MUX_s_1_2_2(or_662_nl, nand_136_nl, fsm_output[3]);
  assign nor_430_nl = ~((~((fsm_output[3]) & (COMP_LOOP_acc_1_cse_6_sva[2:0]==3'b111)
      & (~ (fsm_output[5])))) | nand_245_cse);
  assign and_447_nl = (~ (fsm_output[3])) & (fsm_output[5]) & (COMP_LOOP_acc_1_cse_2_sva[2:0]==3'b111)
      & (~ (fsm_output[9])) & (fsm_output[7]);
  assign not_tmp_249 = MUX_s_1_2_2(nor_430_nl, and_447_nl, fsm_output[6]);
  assign nor_428_nl = ~((fsm_output[6]) | (fsm_output[3]) | (COMP_LOOP_acc_14_psp_sva[1:0]!=2'b11)
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[7]));
  assign nor_429_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[3])) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b11)
      | (fsm_output[5]) | (fsm_output[9]) | (fsm_output[7]));
  assign not_tmp_250 = MUX_s_1_2_2(nor_428_nl, nor_429_nl, fsm_output[4]);
  assign nand_131_nl = ~((COMP_LOOP_acc_1_cse_4_sva[2:0]==3'b111) & (fsm_output[7:3]==5'b01110));
  assign or_688_nl = (COMP_LOOP_acc_1_cse_sva[2:0]!=3'b111) | (fsm_output[7:3]!=5'b00011);
  assign mux_tmp_733 = MUX_s_1_2_2(nand_131_nl, or_688_nl, fsm_output[9]);
  assign and_dcpl_150 = and_dcpl_82 & and_dcpl_72;
  assign or_tmp_672 = nor_813_cse | (fsm_output[7]);
  assign or_tmp_677 = (fsm_output[8]) | (fsm_output[0]) | (fsm_output[7]);
  assign or_tmp_679 = (~((~ (fsm_output[8])) | (fsm_output[0]))) | (fsm_output[7]);
  assign nor_tmp_166 = (fsm_output[0]) & (fsm_output[7]);
  assign or_tmp_681 = (fsm_output[8]) | (~ nor_tmp_166);
  assign mux_tmp_760 = MUX_s_1_2_2(or_90_cse, or_tmp_681, fsm_output[6]);
  assign or_tmp_682 = (~ (fsm_output[8])) | (fsm_output[0]) | (fsm_output[7]);
  assign mux_tmp_773 = MUX_s_1_2_2(or_90_cse, mux_995_cse, fsm_output[6]);
  assign mux_tmp_777 = MUX_s_1_2_2((~ mux_995_cse), or_90_cse, fsm_output[6]);
  assign nor_tmp_168 = ((~ (fsm_output[8])) | (fsm_output[0])) & (fsm_output[7]);
  assign not_tmp_276 = MUX_s_1_2_2((fsm_output[8]), (~ (fsm_output[8])), fsm_output[9]);
  assign mux_tmp_814 = MUX_s_1_2_2((fsm_output[8]), or_831_cse, fsm_output[7]);
  assign mux_822_nl = MUX_s_1_2_2(not_tmp_276, (fsm_output[8]), fsm_output[7]);
  assign mux_tmp_823 = MUX_s_1_2_2(mux_822_nl, or_831_cse, fsm_output[6]);
  assign mux_tmp_825 = MUX_s_1_2_2(mux_tmp_390, mux_tmp_814, fsm_output[6]);
  assign or_750_cse = (fsm_output[0]) | (fsm_output[9]) | (~ (fsm_output[8]));
  assign mux_tmp_833 = MUX_s_1_2_2(not_tmp_121, or_750_cse, fsm_output[7]);
  assign or_tmp_737 = (fsm_output[9]) | (~ (fsm_output[6]));
  assign mux_tmp_860 = MUX_s_1_2_2((~ or_tmp_737), and_434_cse, fsm_output[4]);
  assign or_tmp_738 = (fsm_output[4]) | (~ and_434_cse);
  assign and_310_nl = (fsm_output[0]) & (fsm_output[4]);
  assign mux_tmp_865 = MUX_s_1_2_2((~ or_tmp_737), (fsm_output[6]), and_310_nl);
  assign or_1312_cse = (fsm_output[4]) | (~ (fsm_output[1])) | (fsm_output[6]) |
      (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[7]));
  assign or_798_cse = (fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[2])
      | (~ (fsm_output[8])) | (fsm_output[7]);
  assign nor_371_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[7]));
  assign nor_372_nl = ~((fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign mux_884_nl = MUX_s_1_2_2(nor_371_nl, nor_372_nl, fsm_output[9]);
  assign and_301_nl = (fsm_output[6]) & mux_884_nl;
  assign nor_373_nl = ~((fsm_output[6]) | (fsm_output[9]) | (fsm_output[2]) | (~((fsm_output[8:7]==2'b11))));
  assign mux_885_nl = MUX_s_1_2_2(and_301_nl, nor_373_nl, fsm_output[1]);
  assign nand_194_nl = ~((fsm_output[4]) & mux_885_nl);
  assign mux_886_nl = MUX_s_1_2_2(or_1312_cse, nand_194_nl, fsm_output[5]);
  assign or_797_nl = (fsm_output[6]) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (fsm_output[7]);
  assign nor_375_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[7])));
  assign nor_376_nl = ~((fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[7]));
  assign mux_881_nl = MUX_s_1_2_2(nor_375_nl, nor_376_nl, fsm_output[9]);
  assign nand_66_nl = ~((fsm_output[6]) & mux_881_nl);
  assign mux_882_nl = MUX_s_1_2_2(or_797_nl, nand_66_nl, fsm_output[1]);
  assign mux_883_nl = MUX_s_1_2_2(or_798_cse, mux_882_nl, fsm_output[4]);
  assign or_1313_nl = (fsm_output[5]) | mux_883_nl;
  assign mux_887_nl = MUX_s_1_2_2(mux_886_nl, or_1313_nl, fsm_output[3]);
  assign and_dcpl_151 = ~(mux_887_nl | (fsm_output[0]));
  assign nor_365_cse = ~((~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[9]))
      | (fsm_output[7]) | (~ (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[8]));
  assign nor_366_nl = ~((fsm_output[7]) | (~((fsm_output[1]) & (fsm_output[6]) &
      (fsm_output[8]))));
  assign nor_367_nl = ~((~ (fsm_output[7])) | (fsm_output[1]) | (fsm_output[6]) |
      (fsm_output[8]));
  assign mux_891_nl = MUX_s_1_2_2(nor_366_nl, nor_367_nl, fsm_output[9]);
  assign and_298_nl = nor_265_cse & mux_891_nl;
  assign mux_892_nl = MUX_s_1_2_2(nor_365_cse, and_298_nl, fsm_output[5]);
  assign or_811_nl = (fsm_output[9]) | (fsm_output[7]) | (fsm_output[1]) | (fsm_output[6])
      | (~ (fsm_output[8]));
  assign mux_889_nl = MUX_s_1_2_2(or_811_nl, or_29_cse, fsm_output[4]);
  assign and_299_nl = (fsm_output[6]) & (fsm_output[8]);
  assign nor_369_nl = ~((fsm_output[6]) | (fsm_output[8]));
  assign mux_888_nl = MUX_s_1_2_2(and_299_nl, nor_369_nl, fsm_output[1]);
  assign nand_69_nl = ~((~((~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[7]))))
      & mux_888_nl);
  assign mux_890_nl = MUX_s_1_2_2(mux_889_nl, nand_69_nl, fsm_output[2]);
  assign nor_368_nl = ~((fsm_output[5]) | mux_890_nl);
  assign not_tmp_309 = MUX_s_1_2_2(mux_892_nl, nor_368_nl, fsm_output[3]);
  assign and_dcpl_152 = not_tmp_309 & (fsm_output[0]);
  assign mux_894_nl = MUX_s_1_2_2((fsm_output[3]), (~ (fsm_output[3])), or_722_cse);
  assign nor_750_nl = ~((~((fsm_output[2:1]!=2'b00))) | (fsm_output[3]));
  assign mux_895_nl = MUX_s_1_2_2(mux_894_nl, nor_750_nl, fsm_output[0]);
  assign and_dcpl_156 = mux_895_nl & (~ (fsm_output[4])) & and_dcpl_33 & (~ (fsm_output[7]))
      & not_tmp_82;
  assign and_dcpl_157 = and_dcpl_49 & and_dcpl_63;
  assign mux_tmp_898 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[9]);
  assign mux_tmp_899 = MUX_s_1_2_2((~ mux_tmp_898), (fsm_output[9]), fsm_output[8]);
  assign mux_tmp_900 = MUX_s_1_2_2((~ or_tmp_71), mux_tmp_898, fsm_output[8]);
  assign mux_903_cse = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_1483_cse);
  assign or_823_cse = (~((~ (fsm_output[0])) | (fsm_output[9]))) | (fsm_output[7]);
  assign or_tmp_783 = (fsm_output[9]) | (fsm_output[7]);
  assign mux_tmp_912 = MUX_s_1_2_2((~ or_tmp_72), or_tmp_783, fsm_output[8]);
  assign mux_919_cse = MUX_s_1_2_2(mux_tmp_898, or_tmp_72, fsm_output[8]);
  assign and_296_nl = (fsm_output[8]) & (fsm_output[0]);
  assign mux_923_cse = MUX_s_1_2_2(mux_tmp_898, or_tmp_72, and_296_nl);
  assign mux_928_cse = MUX_s_1_2_2(mux_tmp_899, mux_tmp_912, fsm_output[6]);
  assign mux_929_cse = MUX_s_1_2_2((~ and_312_cse), (fsm_output[9]), fsm_output[8]);
  assign mux_936_cse = MUX_s_1_2_2(or_tmp_783, (fsm_output[9]), fsm_output[0]);
  assign mux_937_cse = MUX_s_1_2_2((~ mux_936_cse), or_tmp_72, fsm_output[8]);
  assign nand_191_nl = ~((fsm_output[1]) & (fsm_output[5]) & (~ (fsm_output[3]))
      & (fsm_output[4]));
  assign mux_tmp_1013 = MUX_s_1_2_2(nand_191_nl, or_843_cse, fsm_output[0]);
  assign or_dcpl_56 = (fsm_output[8:1]!=8'b00000100) | or_1275_cse;
  assign mux_tmp_1037 = MUX_s_1_2_2((~ or_tmp_63), nor_tmp_12, fsm_output[5]);
  assign nor_tmp_223 = (fsm_output[7]) & (fsm_output[4]);
  assign or_953_nl = (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[9]))
      | (fsm_output[7]) | (fsm_output[4]);
  assign or_952_nl = (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[9]) | (fsm_output[7])
      | (~ (fsm_output[4]));
  assign mux_1116_nl = MUX_s_1_2_2(or_953_nl, or_952_nl, fsm_output[5]);
  assign nor_667_nl = ~((fsm_output[6]) | mux_1116_nl);
  assign nor_669_nl = ~((fsm_output[7]) | (fsm_output[4]));
  assign mux_1115_nl = MUX_s_1_2_2(nor_669_nl, nor_tmp_223, fsm_output[9]);
  assign nor_668_nl = ~((~ (fsm_output[6])) | (fsm_output[5]) | (fsm_output[2]) |
      (fsm_output[8]) | (~ mux_1115_nl));
  assign mux_1117_nl = MUX_s_1_2_2(nor_667_nl, nor_668_nl, fsm_output[3]);
  assign or_946_nl = (~ (fsm_output[8])) | (~ (fsm_output[9])) | (fsm_output[7])
      | (fsm_output[4]);
  assign or_945_nl = (fsm_output[8]) | (fsm_output[9]) | (~ (fsm_output[7])) | (fsm_output[4]);
  assign mux_1113_nl = MUX_s_1_2_2(or_946_nl, or_945_nl, fsm_output[2]);
  assign nor_670_nl = ~((fsm_output[6:5]!=2'b10) | mux_1113_nl);
  assign nor_671_nl = ~((fsm_output[5]) | (fsm_output[2]) | (~ (fsm_output[8])) |
      (fsm_output[9]) | (~ nor_tmp_223));
  assign nor_672_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[2])) | (fsm_output[8])
      | (~ (fsm_output[9])) | (fsm_output[7]) | (fsm_output[4]));
  assign mux_1112_nl = MUX_s_1_2_2(nor_671_nl, nor_672_nl, fsm_output[6]);
  assign mux_1114_nl = MUX_s_1_2_2(nor_670_nl, mux_1112_nl, fsm_output[3]);
  assign mux_1118_nl = MUX_s_1_2_2(mux_1117_nl, mux_1114_nl, fsm_output[1]);
  assign and_dcpl_174 = mux_1118_nl & (fsm_output[0]);
  assign and_dcpl_176 = and_dcpl_68 & (fsm_output[2]) & and_dcpl_67;
  assign and_dcpl_177 = and_dcpl_176 & and_dcpl_157;
  assign not_tmp_375 = ~((fsm_output[2]) & (fsm_output[4]));
  assign or_dcpl_62 = (fsm_output[4:2]!=3'b100);
  assign not_tmp_384 = ~((fsm_output[8:6]!=3'b000) | and_tmp_2);
  assign or_1017_nl = (fsm_output[7:5]!=3'b000) | and_dcpl_75;
  assign or_1015_nl = (fsm_output[7:5]!=3'b000) | and_398_cse;
  assign mux_1150_nl = MUX_s_1_2_2(or_1017_nl, or_1015_nl, fsm_output[1]);
  assign and_198_nl = (fsm_output[8]) & mux_1150_nl;
  assign mux_1151_itm = MUX_s_1_2_2(not_tmp_384, and_198_nl, fsm_output[9]);
  assign or_tmp_966 = (fsm_output[5]) | and_dcpl_75;
  assign not_tmp_390 = ~((fsm_output[7:6]!=2'b00) | and_tmp_2);
  assign or_tmp_970 = (fsm_output[6]) | and_tmp_2;
  assign or_tmp_992 = (fsm_output[5]) | (fsm_output[2]) | (~ and_398_cse);
  assign mux_1172_nl = MUX_s_1_2_2((~ or_tmp_992), or_tmp_60, fsm_output[6]);
  assign or_tmp_993 = (fsm_output[7]) | mux_1172_nl;
  assign mux_1174_nl = MUX_s_1_2_2(and_dcpl_53, or_tmp_63, fsm_output[5]);
  assign mux_tmp_1175 = MUX_s_1_2_2(or_tmp_60, mux_1174_nl, fsm_output[6]);
  assign mux_1177_nl = MUX_s_1_2_2(and_292_cse, or_tmp_992, fsm_output[6]);
  assign mux_tmp_1179 = MUX_s_1_2_2((~ mux_82_cse), mux_1177_nl, fsm_output[7]);
  assign mux_tmp_1182 = MUX_s_1_2_2((~ or_tmp_58), or_tmp_966, fsm_output[6]);
  assign mux_tmp_1184 = MUX_s_1_2_2((~ or_tmp_966), or_tmp_966, fsm_output[6]);
  assign mux_1185_nl = MUX_s_1_2_2(or_157_cse, or_dcpl_62, fsm_output[5]);
  assign or_1062_nl = (fsm_output[5:2]!=4'b1100);
  assign mux_1186_nl = MUX_s_1_2_2(mux_1185_nl, or_1062_nl, fsm_output[6]);
  assign mux_tmp_1187 = MUX_s_1_2_2(mux_1186_nl, mux_tmp_1184, fsm_output[7]);
  assign mux_tmp_1189 = MUX_s_1_2_2((~ or_tmp_966), or_tmp_60, fsm_output[6]);
  assign mux_tmp_1190 = MUX_s_1_2_2((~ and_tmp_2), or_tmp_966, fsm_output[6]);
  assign mux_tmp_1191 = MUX_s_1_2_2(mux_tmp_1190, mux_tmp_1189, fsm_output[7]);
  assign mux_tmp_1192 = MUX_s_1_2_2((~ (fsm_output[5])), or_dcpl_39, fsm_output[6]);
  assign mux_tmp_1199 = MUX_s_1_2_2(or_dcpl_39, mux_tmp_81, fsm_output[6]);
  assign mux_tmp_1203 = MUX_s_1_2_2((~ or_tmp_966), (fsm_output[5]), fsm_output[6]);
  assign not_tmp_414 = ~((fsm_output[5:3]==3'b111));
  assign mux_1207_nl = MUX_s_1_2_2(not_tmp_414, (fsm_output[5]), fsm_output[6]);
  assign mux_tmp_1208 = MUX_s_1_2_2(mux_1207_nl, mux_tmp_1192, fsm_output[7]);
  assign mux_1206_nl = MUX_s_1_2_2(mux_tmp_1190, mux_tmp_1192, fsm_output[7]);
  assign mux_1209_itm = MUX_s_1_2_2(mux_tmp_1208, mux_1206_nl, fsm_output[1]);
  assign or_tmp_1034 = (~ (fsm_output[9])) | (fsm_output[4]) | (fsm_output[3]) |
      (fsm_output[7]) | (fsm_output[5]);
  assign and_dcpl_191 = and_dcpl_176 & and_dcpl_50;
  assign or_tmp_1050 = (fsm_output[7]) | mux_tmp_1189;
  assign mux_1269_nl = MUX_s_1_2_2(mux_tmp_1175, mux_tmp_77, fsm_output[7]);
  assign mux_1271_nl = MUX_s_1_2_2(mux_tmp_83, mux_1269_nl, fsm_output[1]);
  assign or_73_nl = (fsm_output[7:6]!=2'b00) | (~ or_tmp_58);
  assign mux_1267_nl = MUX_s_1_2_2(or_tmp_1050, or_73_nl, fsm_output[1]);
  assign mux_tmp_1272 = MUX_s_1_2_2(mux_1271_nl, mux_1267_nl, fsm_output[8]);
  assign mux_90_nl = MUX_s_1_2_2((~ mux_tmp_81), and_tmp_2, fsm_output[6]);
  assign mux_tmp_1276 = MUX_s_1_2_2(mux_90_nl, mux_tmp_1184, fsm_output[7]);
  assign mux_87_nl = MUX_s_1_2_2((~ mux_tmp_81), and_292_cse, fsm_output[6]);
  assign mux_1274_nl = MUX_s_1_2_2(mux_87_nl, mux_tmp_1182, fsm_output[7]);
  assign mux_tmp_1277 = MUX_s_1_2_2(mux_tmp_1276, mux_1274_nl, fsm_output[1]);
  assign mux_1284_nl = MUX_s_1_2_2((~ mux_tmp_1037), and_tmp_2, fsm_output[6]);
  assign mux_1285_nl = MUX_s_1_2_2(mux_1284_nl, mux_tmp_1203, fsm_output[7]);
  assign mux_1286_nl = MUX_s_1_2_2(mux_1285_nl, mux_tmp_1276, fsm_output[1]);
  assign mux_1287_nl = MUX_s_1_2_2(mux_1209_itm, (~ mux_1286_nl), fsm_output[8]);
  assign mux_1281_nl = MUX_s_1_2_2(mux_tmp_1199, mux_tmp_1190, fsm_output[7]);
  assign mux_1282_nl = MUX_s_1_2_2(mux_1281_nl, mux_tmp_83, fsm_output[1]);
  assign mux_1283_nl = MUX_s_1_2_2(mux_1282_nl, or_tmp_1050, fsm_output[8]);
  assign mux_tmp_1288 = MUX_s_1_2_2(mux_1287_nl, mux_1283_nl, fsm_output[9]);
  assign mux_1278_nl = MUX_s_1_2_2(mux_tmp_1208, mux_tmp_1191, fsm_output[1]);
  assign mux_1279_nl = MUX_s_1_2_2(mux_1278_nl, (~ mux_tmp_1277), fsm_output[8]);
  assign mux_1280_nl = MUX_s_1_2_2(mux_1279_nl, mux_tmp_1272, fsm_output[9]);
  assign mux_1289_itm = MUX_s_1_2_2(mux_tmp_1288, mux_1280_nl, fsm_output[0]);
  assign and_dcpl_192 = not_tmp_309 & (~ (fsm_output[0]));
  assign nor_661_nl = ~((fsm_output[6]) | (fsm_output[5]) | (~ (fsm_output[9])) |
      (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[8]));
  assign mux_1299_nl = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[2]);
  assign nor_662_nl = ~((fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[9]) |
      (fsm_output[7]) | mux_1299_nl);
  assign mux_1300_nl = MUX_s_1_2_2(nor_661_nl, nor_662_nl, fsm_output[4]);
  assign nor_663_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[6])) | (fsm_output[5])
      | (~ (fsm_output[9])) | (~ (fsm_output[7])) | (fsm_output[2]) | (fsm_output[8]));
  assign mux_1301_nl = MUX_s_1_2_2(mux_1300_nl, nor_663_nl, fsm_output[3]);
  assign or_1132_nl = (~ (fsm_output[7])) | (~ (fsm_output[2])) | (fsm_output[8]);
  assign mux_1297_nl = MUX_s_1_2_2(or_1132_nl, or_1156_cse, fsm_output[9]);
  assign nor_664_nl = ~((fsm_output[6:4]!=3'b100) | mux_1297_nl);
  assign nor_665_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[8]));
  assign nor_666_nl = ~((fsm_output[6]) | (fsm_output[5]) | (fsm_output[9]) | (~
      (fsm_output[7])) | (fsm_output[2]) | (~ (fsm_output[8])));
  assign mux_1296_nl = MUX_s_1_2_2(nor_665_nl, nor_666_nl, fsm_output[4]);
  assign mux_1298_nl = MUX_s_1_2_2(nor_664_nl, mux_1296_nl, fsm_output[3]);
  assign mux_1302_nl = MUX_s_1_2_2(mux_1301_nl, mux_1298_nl, fsm_output[1]);
  assign and_dcpl_194 = mux_1302_nl & (fsm_output[0]);
  assign not_tmp_458 = ~((fsm_output[1]) & (fsm_output[4]));
  assign mux_tmp_1329 = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[7]);
  assign mux_tmp_1331 = MUX_s_1_2_2(or_tmp_13, or_tmp_5, fsm_output[9]);
  assign mux_1330_nl = MUX_s_1_2_2((~ mux_tmp_1329), or_857_cse, fsm_output[9]);
  assign mux_tmp_1332 = MUX_s_1_2_2(mux_tmp_1331, mux_1330_nl, fsm_output[8]);
  assign or_tmp_1128 = (~ (fsm_output[7])) | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_1340_nl = MUX_s_1_2_2(and_293_cse, mux_tmp_1329, fsm_output[9]);
  assign mux_tmp_1341 = MUX_s_1_2_2((~ mux_1340_nl), mux_tmp_1331, fsm_output[8]);
  assign nor_683_nl = ~((~ (fsm_output[0])) | (fsm_output[6]));
  assign mux_1344_nl = MUX_s_1_2_2(nor_683_nl, (fsm_output[6]), fsm_output[7]);
  assign mux_tmp_1345 = MUX_s_1_2_2(mux_1344_nl, mux_tmp_1329, fsm_output[1]);
  assign or_1199_nl = (~((fsm_output[0]) | (fsm_output[7]))) | (fsm_output[6]);
  assign mux_1347_nl = MUX_s_1_2_2(or_1199_nl, or_tmp_13, fsm_output[1]);
  assign mux_tmp_1348 = MUX_s_1_2_2(mux_1347_nl, or_tmp_5, fsm_output[9]);
  assign mux_1350_nl = MUX_s_1_2_2(or_tmp_5, (~ (fsm_output[6])), fsm_output[9]);
  assign mux_tmp_1351 = MUX_s_1_2_2(mux_1350_nl, or_119_cse, fsm_output[8]);
  assign or_tmp_1137 = (fsm_output[7]) | (fsm_output[0]) | (~ (fsm_output[6]));
  assign mux_tmp_1353 = MUX_s_1_2_2(or_tmp_5, or_tmp_1137, fsm_output[1]);
  assign nor_282_nl = ~(nor_tmp_166 | (fsm_output[6]));
  assign and_256_nl = or_730_cse & (fsm_output[6]);
  assign mux_tmp_1355 = MUX_s_1_2_2(nor_282_nl, and_256_nl, fsm_output[1]);
  assign or_tmp_1142 = (fsm_output[7]) | nand_240_cse;
  assign nor_277_nl = ~((fsm_output[9]) | (~((fsm_output[8]) & (fsm_output[6]) &
      (fsm_output[5]))));
  assign nor_278_nl = ~((fsm_output[9]) | (fsm_output[8]) | (fsm_output[6]) | (~
      (fsm_output[5])));
  assign mux_1388_nl = MUX_s_1_2_2(nor_277_nl, nor_278_nl, fsm_output[1]);
  assign and_252_nl = (fsm_output[4]) & mux_1388_nl;
  assign or_1215_nl = (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[6]))
      | (fsm_output[5]);
  assign or_1214_nl = (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[5]);
  assign mux_1387_nl = MUX_s_1_2_2(or_1215_nl, or_1214_nl, fsm_output[1]);
  assign nor_279_nl = ~((fsm_output[4]) | mux_1387_nl);
  assign mux_1389_nl = MUX_s_1_2_2(and_252_nl, nor_279_nl, fsm_output[2]);
  assign and_251_nl = (fsm_output[7]) & mux_1389_nl;
  assign or_1212_nl = (~ (fsm_output[4])) | (~ (fsm_output[1])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[5]);
  assign nand_182_nl = ~((fsm_output[1]) & (fsm_output[9]) & (fsm_output[8]) & (~
      (fsm_output[6])) & (fsm_output[5]));
  assign or_1209_nl = (fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[6])
      | (fsm_output[5]);
  assign mux_1385_nl = MUX_s_1_2_2(nand_182_nl, or_1209_nl, fsm_output[4]);
  assign mux_1386_nl = MUX_s_1_2_2(or_1212_nl, mux_1385_nl, fsm_output[2]);
  assign nor_280_nl = ~((fsm_output[7]) | mux_1386_nl);
  assign not_tmp_496 = MUX_s_1_2_2(and_251_nl, nor_280_nl, fsm_output[3]);
  assign or_tmp_1157 = ~((fsm_output[9]) & (fsm_output[4]) & (fsm_output[6]) & (~
      (fsm_output[8])));
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_61 & and_dcpl_58 & (fsm_output[9])
      & (fsm_output[0]);
  assign VEC_LOOP_j_sva_11_0_mx0c1 = and_dcpl_61 & and_dcpl_58 & and_dcpl_26;
  assign mux_1024_nl = MUX_s_1_2_2(nor_692_cse, mux_tmp_229, or_1470_cse);
  assign mux_1025_nl = MUX_s_1_2_2(nor_692_cse, mux_1024_nl, fsm_output[2]);
  assign mux_1023_nl = MUX_s_1_2_2(mux_tmp_229, nor_tmp_21, or_722_cse);
  assign mux_1026_cse = MUX_s_1_2_2(mux_1025_nl, mux_1023_nl, fsm_output[3]);
  assign or_859_nl = (fsm_output[6:4]!=3'b000);
  assign modExp_result_sva_mx0c0 = MUX_s_1_2_2(mux_1026_cse, nor_tmp_21, or_859_nl);
  assign modExp_base_sva_mx0c1 = and_dcpl_70 & and_dcpl_72;
  assign tmp_10_lpi_4_dfm_mx0c1 = and_dcpl_103 & and_dcpl_122 & nor_401_cse;
  assign tmp_10_lpi_4_dfm_mx0c2 = and_dcpl_82 & and_dcpl_16 & nor_401_cse;
  assign tmp_10_lpi_4_dfm_mx0c3 = and_dcpl_115 & and_dcpl_97;
  assign tmp_10_lpi_4_dfm_mx0c4 = and_dcpl_76 & and_dcpl_102;
  assign tmp_10_lpi_4_dfm_mx0c5 = and_dcpl_133 & and_dcpl_108;
  assign tmp_10_lpi_4_dfm_mx0c6 = and_dcpl_70 & and_dcpl_78 & and_dcpl_26;
  assign tmp_10_lpi_4_dfm_mx0c7 = and_dcpl_124 & and_dcpl_33 & and_dcpl_96 & and_dcpl_26;
  assign nl_STAGE_LOOP_acc_nl = (STAGE_LOOP_i_3_0_sva_2[3:1]) + 3'b011;
  assign STAGE_LOOP_acc_nl = nl_STAGE_LOOP_acc_nl[2:0];
  assign STAGE_LOOP_acc_itm_2_1 = readslicef_3_1_2(STAGE_LOOP_acc_nl);
  assign and_244_m1c = and_dcpl_76 & and_dcpl_66;
  assign nor_274_nl = ~((~ (fsm_output[9])) | (fsm_output[4]) | not_tmp_29);
  assign nor_275_nl = ~((~ (fsm_output[9])) | (fsm_output[4]) | (fsm_output[6]) |
      (fsm_output[8]));
  assign mux_1394_nl = MUX_s_1_2_2(nor_274_nl, nor_275_nl, fsm_output[1]);
  assign nand_89_nl = ~((fsm_output[2]) & mux_1394_nl);
  assign or_1227_nl = (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[6]) | (~
      (fsm_output[8]));
  assign mux_1393_nl = MUX_s_1_2_2(or_tmp_1157, or_1227_nl, fsm_output[1]);
  assign or_1228_nl = (fsm_output[2]) | mux_1393_nl;
  assign mux_1395_nl = MUX_s_1_2_2(nand_89_nl, or_1228_nl, fsm_output[5]);
  assign nor_273_nl = ~((fsm_output[7]) | mux_1395_nl);
  assign or_1224_nl = (fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[8]);
  assign mux_1391_nl = MUX_s_1_2_2(or_1224_nl, or_tmp_1157, fsm_output[1]);
  assign or_1222_nl = (fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[6])
      | (~ (fsm_output[8]));
  assign mux_1392_nl = MUX_s_1_2_2(mux_1391_nl, or_1222_nl, fsm_output[2]);
  assign nor_276_nl = ~((~ (fsm_output[7])) | (fsm_output[5]) | mux_1392_nl);
  assign mux_1396_nl = MUX_s_1_2_2(nor_273_nl, nor_276_nl, fsm_output[3]);
  assign and_250_m1c = mux_1396_nl & (fsm_output[0]);
  assign and_98_nl = and_dcpl_82 & and_dcpl_79;
  assign nor_655_nl = ~((fsm_output[8]) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (fsm_output[5]));
  assign nor_656_nl = ~((~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[7]) |
      (fsm_output[5]));
  assign mux_459_nl = MUX_s_1_2_2(nor_655_nl, nor_656_nl, fsm_output[9]);
  assign nand_235_nl = ~((fsm_output[4:3]==2'b11) & mux_459_nl);
  assign or_1386_nl = (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[8]) | (~
      (fsm_output[2])) | (fsm_output[7]) | (fsm_output[5]);
  assign or_1387_nl = (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[2])
      | (fsm_output[7]) | (~ (fsm_output[5]));
  assign mux_458_nl = MUX_s_1_2_2(or_1386_nl, or_1387_nl, fsm_output[4]);
  assign mux_460_nl = MUX_s_1_2_2(nand_235_nl, mux_458_nl, fsm_output[6]);
  assign or_234_nl = (~ (fsm_output[8])) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[5]);
  assign or_233_nl = (~ (fsm_output[8])) | (fsm_output[2]) | (~ (fsm_output[7]))
      | (fsm_output[5]);
  assign mux_455_nl = MUX_s_1_2_2(or_234_nl, or_233_nl, fsm_output[9]);
  assign or_232_nl = (~ (fsm_output[9])) | (fsm_output[8]) | (~((fsm_output[2]) &
      (fsm_output[7]) & (fsm_output[5])));
  assign mux_456_nl = MUX_s_1_2_2(mux_455_nl, or_232_nl, fsm_output[3]);
  assign or_1388_nl = (fsm_output[4]) | mux_456_nl;
  assign or_1389_nl = (~ (fsm_output[4])) | (~ (fsm_output[3])) | (fsm_output[9])
      | (~ (fsm_output[8])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[5]);
  assign mux_457_nl = MUX_s_1_2_2(or_1388_nl, or_1389_nl, fsm_output[6]);
  assign mux_461_nl = MUX_s_1_2_2(mux_460_nl, mux_457_nl, fsm_output[1]);
  assign nor_740_nl = ~(mux_461_nl | (fsm_output[0]));
  assign nor_653_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[6])) | (~ (fsm_output[5]))
      | (fsm_output[2]) | (fsm_output[3]));
  assign nor_654_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[5]) | (~((fsm_output[3:2]==2'b11))));
  assign mux_462_nl = MUX_s_1_2_2(nor_653_nl, nor_654_nl, fsm_output[0]);
  assign and_103_nl = mux_462_nl & (fsm_output[4]) & (fsm_output[7]) & not_tmp_82;
  assign nor_651_nl = ~((fsm_output[1]) | (~((fsm_output[6]) & (fsm_output[3]) &
      (fsm_output[4]))));
  assign nor_652_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[3]) |
      (fsm_output[4]));
  assign mux_463_nl = MUX_s_1_2_2(nor_651_nl, nor_652_nl, fsm_output[0]);
  assign and_110_nl = mux_463_nl & (fsm_output[2]) & (~ (fsm_output[5])) & (~ (fsm_output[7]))
      & and_dcpl_91;
  assign nor_649_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[7])) | (fsm_output[5])
      | (~ (fsm_output[2])) | (fsm_output[4]));
  assign nor_650_nl = ~((fsm_output[1]) | (fsm_output[7]) | (~ (fsm_output[5])) |
      (fsm_output[2]) | (~ (fsm_output[4])));
  assign mux_464_nl = MUX_s_1_2_2(nor_649_nl, nor_650_nl, fsm_output[0]);
  assign and_116_nl = mux_464_nl & (~ (fsm_output[3])) & (fsm_output[6]) & and_dcpl_91;
  assign nor_647_nl = ~((~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[1]) |
      (fsm_output[7]) | (fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[3]));
  assign and_449_nl = (~ (fsm_output[9])) & (fsm_output[8]) & (fsm_output[1]) & (fsm_output[7])
      & (fsm_output[6]) & (~ (fsm_output[5])) & (fsm_output[3]);
  assign mux_465_nl = MUX_s_1_2_2(nor_647_nl, and_449_nl, fsm_output[0]);
  assign and_121_nl = mux_465_nl & (fsm_output[4]) & (~ (fsm_output[2]));
  assign nor_645_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[7])) | (fsm_output[6])
      | (fsm_output[2]) | (~ and_398_cse));
  assign nor_646_nl = ~((fsm_output[1]) | (fsm_output[7]) | (~ (fsm_output[6])) |
      (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[4]));
  assign mux_466_nl = MUX_s_1_2_2(nor_645_nl, nor_646_nl, fsm_output[0]);
  assign and_127_nl = mux_466_nl & (~ (fsm_output[5])) & (~ (fsm_output[8])) & (fsm_output[9]);
  assign nor_643_nl = ~((~ (fsm_output[8])) | (fsm_output[1]) | (fsm_output[7]) |
      (fsm_output[5]) | (fsm_output[3]));
  assign nor_644_nl = ~((fsm_output[8]) | (~((fsm_output[1]) & (fsm_output[7]) &
      (fsm_output[5]) & (fsm_output[3]))));
  assign mux_467_nl = MUX_s_1_2_2(nor_643_nl, nor_644_nl, fsm_output[0]);
  assign and_135_nl = mux_467_nl & (~ (fsm_output[4])) & (fsm_output[2]) & (~ (fsm_output[6]))
      & (fsm_output[9]);
  assign and_382_nl = (fsm_output[1]) & (fsm_output[6]) & (fsm_output[5]) & (fsm_output[2])
      & (~ (fsm_output[4]));
  assign nor_642_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[5]) | (fsm_output[2])
      | (~ (fsm_output[4])));
  assign mux_468_nl = MUX_s_1_2_2(and_382_nl, nor_642_nl, fsm_output[0]);
  assign and_145_nl = mux_468_nl & (fsm_output[3]) & (~ (fsm_output[7])) & (fsm_output[8])
      & (fsm_output[9]);
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_9_11_2(COMP_LOOP_acc_psp_sva_1, (z_out_6_12_1[11:3]),
      COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_12_1_1_sva[11:3]), (COMP_LOOP_acc_1_cse_2_sva[11:3]),
      (COMP_LOOP_acc_11_psp_sva[10:2]), (COMP_LOOP_acc_1_cse_4_sva[11:3]), (COMP_LOOP_acc_13_psp_sva[9:1]),
      (COMP_LOOP_acc_1_cse_6_sva[11:3]), (COMP_LOOP_acc_14_psp_sva[10:2]), (COMP_LOOP_acc_1_cse_sva[11:3]),
      {and_dcpl_71 , COMP_LOOP_or_3_cse , and_98_nl , nor_740_nl , and_103_nl , and_110_nl
      , and_116_nl , and_121_nl , and_127_nl , and_135_nl , and_145_nl});
  assign vec_rsc_0_0_i_da_d_pff = modulo_result_mux_1_cse;
  assign or_1375_nl = (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | mux_tmp_473;
  assign mux_484_nl = MUX_s_1_2_2(or_1375_nl, mux_483_cse, fsm_output[2]);
  assign or_1378_nl = (VEC_LOOP_j_sva_11_0[0]) | mux_tmp_472;
  assign mux_482_nl = MUX_s_1_2_2(nand_232_cse, or_1378_nl, fsm_output[2]);
  assign mux_485_nl = MUX_s_1_2_2(mux_484_nl, mux_482_nl, fsm_output[8]);
  assign nand_233_nl = ~((fsm_output[4]) & not_tmp_166);
  assign mux_479_nl = MUX_s_1_2_2(nand_233_nl, or_1379_cse, fsm_output[2]);
  assign mux_476_nl = MUX_s_1_2_2(or_277_cse, mux_tmp_469, fsm_output[6]);
  assign or_1382_nl = (fsm_output[4]) | mux_476_nl;
  assign mux_478_nl = MUX_s_1_2_2(mux_477_cse, or_1382_nl, fsm_output[2]);
  assign mux_480_nl = MUX_s_1_2_2(mux_479_nl, mux_478_nl, fsm_output[8]);
  assign mux_486_nl = MUX_s_1_2_2(mux_485_nl, mux_480_nl, fsm_output[1]);
  assign or_1383_nl = (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | mux_tmp_473;
  assign or_1384_nl = (~ (fsm_output[2])) | (VEC_LOOP_j_sva_11_0[0]) | mux_tmp_472;
  assign mux_474_nl = MUX_s_1_2_2(or_1383_nl, or_1384_nl, fsm_output[8]);
  assign nand_234_nl = ~(nor_265_cse & not_tmp_166);
  assign or_1385_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | mux_tmp_469;
  assign mux_471_nl = MUX_s_1_2_2(nand_234_nl, or_1385_nl, fsm_output[8]);
  assign mux_475_nl = MUX_s_1_2_2(mux_474_nl, mux_471_nl, fsm_output[1]);
  assign or_260_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000);
  assign mux_487_nl = MUX_s_1_2_2(mux_486_nl, mux_475_nl, or_260_nl);
  assign vec_rsc_0_0_i_wea_d_pff = ~(mux_487_nl | (fsm_output[0]));
  assign nor_612_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_6_12_1[2:0]!=3'b000) |
      (fsm_output[4]) | not_tmp_171);
  assign nor_613_nl = ~((z_out_6_12_1[2:0]!=3'b000) | (fsm_output[7:3]!=5'b01110));
  assign mux_499_nl = MUX_s_1_2_2(nor_612_nl, nor_613_nl, fsm_output[9]);
  assign nor_614_nl = ~((z_out_6_12_1[2:0]!=3'b000) | (~ (fsm_output[9])) | (~ (fsm_output[6]))
      | (fsm_output[5]) | not_tmp_170);
  assign mux_500_nl = MUX_s_1_2_2(mux_499_nl, nor_614_nl, fsm_output[1]);
  assign nor_615_nl = ~((z_out_6_12_1[2:0]!=3'b000) | (fsm_output[7:3]!=5'b01011));
  assign nor_616_nl = ~((z_out_6_12_1[2:0]!=3'b000) | (fsm_output[7:3]!=5'b00000));
  assign mux_498_nl = MUX_s_1_2_2(nor_615_nl, nor_616_nl, fsm_output[9]);
  assign and_377_nl = (fsm_output[1]) & mux_498_nl;
  assign mux_501_nl = MUX_s_1_2_2(mux_500_nl, and_377_nl, fsm_output[2]);
  assign nor_617_nl = ~((z_out_6_12_1[2:0]!=3'b000) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[3])
      | (fsm_output[7]));
  assign or_311_nl = (z_out_6_12_1[2:0]!=3'b000) | (fsm_output[6:5]!=2'b00) | not_tmp_170;
  assign or_309_nl = (z_out_6_12_1[2:0]!=3'b000) | (fsm_output[7:3]!=5'b01000);
  assign mux_496_nl = MUX_s_1_2_2(or_311_nl, or_309_nl, fsm_output[9]);
  assign nor_618_nl = ~((fsm_output[1]) | mux_496_nl);
  assign mux_497_nl = MUX_s_1_2_2(nor_617_nl, nor_618_nl, fsm_output[2]);
  assign mux_502_nl = MUX_s_1_2_2(mux_501_nl, mux_497_nl, fsm_output[8]);
  assign nor_619_nl = ~((VEC_LOOP_j_sva_11_0[2:1]!=2'b00) | (~ (fsm_output[1])) |
      (fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[7:3]!=5'b00110));
  assign nor_620_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b000) | (fsm_output[6:5]!=2'b00)
      | not_tmp_170);
  assign nor_621_nl = ~((COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b000) | (fsm_output[7:3]!=5'b01000));
  assign mux_492_nl = MUX_s_1_2_2(nor_620_nl, nor_621_nl, fsm_output[9]);
  assign nor_622_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00) | (~ (fsm_output[9]))
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[6:4]!=3'b010) | not_tmp_171);
  assign mux_493_nl = MUX_s_1_2_2(mux_492_nl, nor_622_nl, fsm_output[1]);
  assign and_378_nl = COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & mux_493_nl;
  assign mux_494_nl = MUX_s_1_2_2(nor_619_nl, and_378_nl, fsm_output[2]);
  assign nor_623_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | mux_tmp_488);
  assign mux_489_nl = MUX_s_1_2_2(nor_623_nl, nor_624_cse, fsm_output[1]);
  assign nor_625_nl = ~((fsm_output[1]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | mux_tmp_488);
  assign mux_490_nl = MUX_s_1_2_2(mux_489_nl, nor_625_nl, or_294_cse);
  assign nor_626_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00)
      | (~ (fsm_output[1])) | (fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[7:3]!=5'b00000));
  assign mux_491_nl = MUX_s_1_2_2(mux_490_nl, nor_626_nl, fsm_output[2]);
  assign mux_495_nl = MUX_s_1_2_2(mux_494_nl, mux_491_nl, fsm_output[8]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_502_nl,
      mux_495_nl, fsm_output[0]);
  assign or_1366_nl = (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | mux_tmp_473;
  assign mux_519_nl = MUX_s_1_2_2(or_1366_nl, mux_483_cse, fsm_output[2]);
  assign nand_228_nl = ~((VEC_LOOP_j_sva_11_0[0]) & not_tmp_178);
  assign mux_517_nl = MUX_s_1_2_2(nand_232_cse, nand_228_nl, fsm_output[2]);
  assign mux_520_nl = MUX_s_1_2_2(mux_519_nl, mux_517_nl, fsm_output[8]);
  assign nand_229_nl = ~((fsm_output[4]) & not_tmp_177);
  assign mux_514_nl = MUX_s_1_2_2(nand_229_nl, or_1379_cse, fsm_output[2]);
  assign mux_511_nl = MUX_s_1_2_2(or_277_cse, mux_tmp_504, fsm_output[6]);
  assign or_1372_nl = (fsm_output[4]) | mux_511_nl;
  assign mux_513_nl = MUX_s_1_2_2(mux_477_cse, or_1372_nl, fsm_output[2]);
  assign mux_515_nl = MUX_s_1_2_2(mux_514_nl, mux_513_nl, fsm_output[8]);
  assign mux_521_nl = MUX_s_1_2_2(mux_520_nl, mux_515_nl, fsm_output[1]);
  assign or_1373_nl = (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | mux_tmp_473;
  assign nand_230_nl = ~((fsm_output[2]) & (VEC_LOOP_j_sva_11_0[0]) & not_tmp_178);
  assign mux_509_nl = MUX_s_1_2_2(or_1373_nl, nand_230_nl, fsm_output[8]);
  assign nand_231_nl = ~(nor_265_cse & not_tmp_177);
  assign or_1374_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | mux_tmp_504;
  assign mux_506_nl = MUX_s_1_2_2(nand_231_nl, or_1374_nl, fsm_output[8]);
  assign mux_510_nl = MUX_s_1_2_2(mux_509_nl, mux_506_nl, fsm_output[1]);
  assign or_321_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001);
  assign mux_522_nl = MUX_s_1_2_2(mux_521_nl, mux_510_nl, or_321_nl);
  assign vec_rsc_0_1_i_wea_d_pff = ~(mux_522_nl | (fsm_output[0]));
  assign nor_582_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_6_12_1[2:0]!=3'b001) |
      (fsm_output[4]) | not_tmp_171);
  assign nor_583_nl = ~((z_out_6_12_1[2:0]!=3'b001) | (fsm_output[7:3]!=5'b01110));
  assign mux_534_nl = MUX_s_1_2_2(nor_582_nl, nor_583_nl, fsm_output[9]);
  assign nor_584_nl = ~((z_out_6_12_1[2:0]!=3'b001) | (~ (fsm_output[9])) | (~ (fsm_output[6]))
      | (fsm_output[5]) | not_tmp_170);
  assign mux_535_nl = MUX_s_1_2_2(mux_534_nl, nor_584_nl, fsm_output[1]);
  assign nor_585_nl = ~((z_out_6_12_1[2:0]!=3'b001) | (fsm_output[7:3]!=5'b01011));
  assign nor_586_nl = ~((z_out_6_12_1[2:0]!=3'b001) | (fsm_output[7:3]!=5'b00000));
  assign mux_533_nl = MUX_s_1_2_2(nor_585_nl, nor_586_nl, fsm_output[9]);
  assign and_370_nl = (fsm_output[1]) & mux_533_nl;
  assign mux_536_nl = MUX_s_1_2_2(mux_535_nl, and_370_nl, fsm_output[2]);
  assign nor_587_nl = ~((z_out_6_12_1[2:0]!=3'b001) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[3])
      | (fsm_output[7]));
  assign or_369_nl = (z_out_6_12_1[2:0]!=3'b001) | (fsm_output[6:5]!=2'b00) | not_tmp_170;
  assign or_367_nl = (z_out_6_12_1[2:0]!=3'b001) | (fsm_output[7:3]!=5'b01000);
  assign mux_531_nl = MUX_s_1_2_2(or_369_nl, or_367_nl, fsm_output[9]);
  assign nor_588_nl = ~((fsm_output[1]) | mux_531_nl);
  assign mux_532_nl = MUX_s_1_2_2(nor_587_nl, nor_588_nl, fsm_output[2]);
  assign mux_537_nl = MUX_s_1_2_2(mux_536_nl, mux_532_nl, fsm_output[8]);
  assign nor_589_nl = ~((VEC_LOOP_j_sva_11_0[2:1]!=2'b00) | (~ (fsm_output[1])) |
      (fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b00110));
  assign nor_590_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b001) | (fsm_output[6:5]!=2'b00)
      | not_tmp_170);
  assign nor_591_nl = ~((COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b001) | (fsm_output[7:3]!=5'b01000));
  assign mux_527_nl = MUX_s_1_2_2(nor_590_nl, nor_591_nl, fsm_output[9]);
  assign nor_592_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b00) | (~ (fsm_output[9]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[6:4]!=3'b010) | not_tmp_171);
  assign mux_528_nl = MUX_s_1_2_2(mux_527_nl, nor_592_nl, fsm_output[1]);
  assign and_371_nl = COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & mux_528_nl;
  assign mux_529_nl = MUX_s_1_2_2(nor_589_nl, and_371_nl, fsm_output[2]);
  assign nor_593_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | mux_tmp_523);
  assign mux_524_nl = MUX_s_1_2_2(nor_593_nl, nor_594_cse, fsm_output[1]);
  assign nor_595_nl = ~((fsm_output[1]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | mux_tmp_523);
  assign mux_525_nl = MUX_s_1_2_2(mux_524_nl, nor_595_nl, or_294_cse);
  assign nor_596_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b00)
      | (~ (fsm_output[1])) | (fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b00000));
  assign mux_526_nl = MUX_s_1_2_2(mux_525_nl, nor_596_nl, fsm_output[2]);
  assign mux_530_nl = MUX_s_1_2_2(mux_529_nl, mux_526_nl, fsm_output[8]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_537_nl,
      mux_530_nl, fsm_output[0]);
  assign nand_222_nl = ~(nor_114_cse & not_tmp_190);
  assign mux_554_nl = MUX_s_1_2_2(nand_222_nl, mux_483_cse, fsm_output[2]);
  assign or_1359_nl = (VEC_LOOP_j_sva_11_0[0]) | mux_tmp_542;
  assign mux_552_nl = MUX_s_1_2_2(nand_232_cse, or_1359_nl, fsm_output[2]);
  assign mux_555_nl = MUX_s_1_2_2(mux_554_nl, mux_552_nl, fsm_output[8]);
  assign nand_224_nl = ~((fsm_output[4]) & not_tmp_189);
  assign mux_549_nl = MUX_s_1_2_2(nand_224_nl, or_1379_cse, fsm_output[2]);
  assign mux_546_nl = MUX_s_1_2_2(or_277_cse, mux_tmp_539, fsm_output[6]);
  assign or_1363_nl = (fsm_output[4]) | mux_546_nl;
  assign mux_548_nl = MUX_s_1_2_2(mux_477_cse, or_1363_nl, fsm_output[2]);
  assign mux_550_nl = MUX_s_1_2_2(mux_549_nl, mux_548_nl, fsm_output[8]);
  assign mux_556_nl = MUX_s_1_2_2(mux_555_nl, mux_550_nl, fsm_output[1]);
  assign nand_225_nl = ~(nor_112_cse & not_tmp_190);
  assign or_1364_nl = (~ (fsm_output[2])) | (VEC_LOOP_j_sva_11_0[0]) | mux_tmp_542;
  assign mux_544_nl = MUX_s_1_2_2(nand_225_nl, or_1364_nl, fsm_output[8]);
  assign nand_226_nl = ~(nor_265_cse & not_tmp_189);
  assign or_1365_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | mux_tmp_539;
  assign mux_541_nl = MUX_s_1_2_2(nand_226_nl, or_1365_nl, fsm_output[8]);
  assign mux_545_nl = MUX_s_1_2_2(mux_544_nl, mux_541_nl, fsm_output[1]);
  assign or_379_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010);
  assign mux_557_nl = MUX_s_1_2_2(mux_556_nl, mux_545_nl, or_379_nl);
  assign vec_rsc_0_2_i_wea_d_pff = ~(mux_557_nl | (fsm_output[0]));
  assign nor_552_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_6_12_1[2:0]!=3'b010) |
      (fsm_output[4]) | not_tmp_171);
  assign nor_553_nl = ~((z_out_6_12_1[2:0]!=3'b010) | (fsm_output[7:3]!=5'b01110));
  assign mux_569_nl = MUX_s_1_2_2(nor_552_nl, nor_553_nl, fsm_output[9]);
  assign nor_554_nl = ~((z_out_6_12_1[2:0]!=3'b010) | (~ (fsm_output[9])) | (~ (fsm_output[6]))
      | (fsm_output[5]) | not_tmp_170);
  assign mux_570_nl = MUX_s_1_2_2(mux_569_nl, nor_554_nl, fsm_output[1]);
  assign nor_555_nl = ~((z_out_6_12_1[2:0]!=3'b010) | (fsm_output[7:3]!=5'b01011));
  assign nor_556_nl = ~((z_out_6_12_1[2:0]!=3'b010) | (fsm_output[7:3]!=5'b00000));
  assign mux_568_nl = MUX_s_1_2_2(nor_555_nl, nor_556_nl, fsm_output[9]);
  assign and_363_nl = (fsm_output[1]) & mux_568_nl;
  assign mux_571_nl = MUX_s_1_2_2(mux_570_nl, and_363_nl, fsm_output[2]);
  assign nor_557_nl = ~((z_out_6_12_1[2:0]!=3'b010) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[3])
      | (fsm_output[7]));
  assign or_425_nl = (z_out_6_12_1[2:0]!=3'b010) | (fsm_output[6:5]!=2'b00) | not_tmp_170;
  assign or_423_nl = (z_out_6_12_1[2:0]!=3'b010) | (fsm_output[7:3]!=5'b01000);
  assign mux_566_nl = MUX_s_1_2_2(or_425_nl, or_423_nl, fsm_output[9]);
  assign nor_558_nl = ~((fsm_output[1]) | mux_566_nl);
  assign mux_567_nl = MUX_s_1_2_2(nor_557_nl, nor_558_nl, fsm_output[2]);
  assign mux_572_nl = MUX_s_1_2_2(mux_571_nl, mux_567_nl, fsm_output[8]);
  assign nor_559_nl = ~((VEC_LOOP_j_sva_11_0[2:1]!=2'b01) | (~ (fsm_output[1])) |
      (fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[7:3]!=5'b00110));
  assign nor_560_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b010) | (fsm_output[6:5]!=2'b00)
      | not_tmp_170);
  assign nor_561_nl = ~((COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b010) | (fsm_output[7:3]!=5'b01000));
  assign mux_562_nl = MUX_s_1_2_2(nor_560_nl, nor_561_nl, fsm_output[9]);
  assign nor_562_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01) | (~ (fsm_output[9]))
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[6:4]!=3'b010) | not_tmp_171);
  assign mux_563_nl = MUX_s_1_2_2(mux_562_nl, nor_562_nl, fsm_output[1]);
  assign and_364_nl = COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & mux_563_nl;
  assign mux_564_nl = MUX_s_1_2_2(nor_559_nl, and_364_nl, fsm_output[2]);
  assign nor_563_nl = ~((fsm_output[1]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | mux_tmp_558);
  assign nor_564_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | mux_tmp_558);
  assign mux_559_nl = MUX_s_1_2_2(nor_564_nl, nor_624_cse, fsm_output[1]);
  assign mux_560_nl = MUX_s_1_2_2(nor_563_nl, mux_559_nl, nor_115_cse);
  assign nor_566_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01)
      | (~ (fsm_output[1])) | (fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[7:3]!=5'b00000));
  assign mux_561_nl = MUX_s_1_2_2(mux_560_nl, nor_566_nl, fsm_output[2]);
  assign mux_565_nl = MUX_s_1_2_2(mux_564_nl, mux_561_nl, fsm_output[8]);
  assign vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_572_nl,
      mux_565_nl, fsm_output[0]);
  assign nand_215_nl = ~((VEC_LOOP_j_sva_11_0[1:0]==2'b11) & not_tmp_190);
  assign mux_589_nl = MUX_s_1_2_2(nand_215_nl, mux_483_cse, fsm_output[2]);
  assign nand_217_nl = ~((VEC_LOOP_j_sva_11_0[0]) & not_tmp_202);
  assign mux_587_nl = MUX_s_1_2_2(nand_232_cse, nand_217_nl, fsm_output[2]);
  assign mux_590_nl = MUX_s_1_2_2(mux_589_nl, mux_587_nl, fsm_output[8]);
  assign nand_218_nl = ~((fsm_output[4]) & not_tmp_201);
  assign mux_584_nl = MUX_s_1_2_2(nand_218_nl, or_1379_cse, fsm_output[2]);
  assign mux_581_nl = MUX_s_1_2_2(or_277_cse, mux_tmp_574, fsm_output[6]);
  assign or_1355_nl = (fsm_output[4]) | mux_581_nl;
  assign mux_583_nl = MUX_s_1_2_2(mux_477_cse, or_1355_nl, fsm_output[2]);
  assign mux_585_nl = MUX_s_1_2_2(mux_584_nl, mux_583_nl, fsm_output[8]);
  assign mux_591_nl = MUX_s_1_2_2(mux_590_nl, mux_585_nl, fsm_output[1]);
  assign nand_219_nl = ~(nor_122_cse & not_tmp_190);
  assign nand_220_nl = ~((fsm_output[2]) & (VEC_LOOP_j_sva_11_0[0]) & not_tmp_202);
  assign mux_579_nl = MUX_s_1_2_2(nand_219_nl, nand_220_nl, fsm_output[8]);
  assign nand_221_nl = ~(nor_265_cse & not_tmp_201);
  assign or_1356_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | mux_tmp_574;
  assign mux_576_nl = MUX_s_1_2_2(nand_221_nl, or_1356_nl, fsm_output[8]);
  assign mux_580_nl = MUX_s_1_2_2(mux_579_nl, mux_576_nl, fsm_output[1]);
  assign or_435_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b011);
  assign mux_592_nl = MUX_s_1_2_2(mux_591_nl, mux_580_nl, or_435_nl);
  assign vec_rsc_0_3_i_wea_d_pff = ~(mux_592_nl | (fsm_output[0]));
  assign nor_522_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_6_12_1[2:0]!=3'b011) |
      (fsm_output[4]) | not_tmp_171);
  assign nor_523_nl = ~((z_out_6_12_1[2:0]!=3'b011) | (fsm_output[7:3]!=5'b01110));
  assign mux_604_nl = MUX_s_1_2_2(nor_522_nl, nor_523_nl, fsm_output[9]);
  assign nor_524_nl = ~((z_out_6_12_1[2:0]!=3'b011) | (~ (fsm_output[9])) | (~ (fsm_output[6]))
      | (fsm_output[5]) | not_tmp_170);
  assign mux_605_nl = MUX_s_1_2_2(mux_604_nl, nor_524_nl, fsm_output[1]);
  assign nor_525_nl = ~((z_out_6_12_1[2:0]!=3'b011) | (fsm_output[7:3]!=5'b01011));
  assign nor_526_nl = ~((z_out_6_12_1[2:0]!=3'b011) | (fsm_output[7:3]!=5'b00000));
  assign mux_603_nl = MUX_s_1_2_2(nor_525_nl, nor_526_nl, fsm_output[9]);
  assign and_354_nl = (fsm_output[1]) & mux_603_nl;
  assign mux_606_nl = MUX_s_1_2_2(mux_605_nl, and_354_nl, fsm_output[2]);
  assign nor_527_nl = ~((z_out_6_12_1[2:0]!=3'b011) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[3])
      | (fsm_output[7]));
  assign or_478_nl = (z_out_6_12_1[2:0]!=3'b011) | (fsm_output[6:5]!=2'b00) | not_tmp_170;
  assign or_476_nl = (z_out_6_12_1[2:0]!=3'b011) | (fsm_output[7:3]!=5'b01000);
  assign mux_601_nl = MUX_s_1_2_2(or_478_nl, or_476_nl, fsm_output[9]);
  assign nor_528_nl = ~((fsm_output[1]) | mux_601_nl);
  assign mux_602_nl = MUX_s_1_2_2(nor_527_nl, nor_528_nl, fsm_output[2]);
  assign mux_607_nl = MUX_s_1_2_2(mux_606_nl, mux_602_nl, fsm_output[8]);
  assign nor_529_nl = ~((VEC_LOOP_j_sva_11_0[2:1]!=2'b01) | (~ (fsm_output[1])) |
      (fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b00110));
  assign nor_530_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b011) | (fsm_output[6:5]!=2'b00)
      | not_tmp_170);
  assign nor_531_nl = ~((COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b011) | (fsm_output[7:3]!=5'b01000));
  assign mux_597_nl = MUX_s_1_2_2(nor_530_nl, nor_531_nl, fsm_output[9]);
  assign nor_532_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b01) | (~ (fsm_output[9]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[6:4]!=3'b010) | not_tmp_171);
  assign mux_598_nl = MUX_s_1_2_2(mux_597_nl, nor_532_nl, fsm_output[1]);
  assign and_355_nl = COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & mux_598_nl;
  assign mux_599_nl = MUX_s_1_2_2(nor_529_nl, and_355_nl, fsm_output[2]);
  assign nor_533_nl = ~((fsm_output[1]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | mux_tmp_593);
  assign nor_534_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | mux_tmp_593);
  assign mux_594_nl = MUX_s_1_2_2(nor_534_nl, nor_594_cse, fsm_output[1]);
  assign mux_595_nl = MUX_s_1_2_2(nor_533_nl, mux_594_nl, nor_115_cse);
  assign nor_536_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b01)
      | (~ (fsm_output[1])) | (fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b00000));
  assign mux_596_nl = MUX_s_1_2_2(mux_595_nl, nor_536_nl, fsm_output[2]);
  assign mux_600_nl = MUX_s_1_2_2(mux_599_nl, mux_596_nl, fsm_output[8]);
  assign vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_607_nl,
      mux_600_nl, fsm_output[0]);
  assign or_1339_nl = (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | mux_tmp_620;
  assign or_1340_nl = (~ (fsm_output[2])) | (VEC_LOOP_j_sva_11_0[0]) | mux_tmp_616;
  assign mux_625_nl = MUX_s_1_2_2(or_1339_nl, or_1340_nl, fsm_output[8]);
  assign nand_212_nl = ~(nor_265_cse & not_tmp_214);
  assign or_1341_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | mux_tmp_609;
  assign mux_624_nl = MUX_s_1_2_2(nand_212_nl, or_1341_nl, fsm_output[8]);
  assign mux_626_nl = MUX_s_1_2_2(mux_625_nl, mux_624_nl, fsm_output[1]);
  assign or_1342_nl = (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | mux_tmp_620;
  assign mux_621_nl = MUX_s_1_2_2(or_1342_nl, mux_483_cse, fsm_output[2]);
  assign or_1345_nl = (VEC_LOOP_j_sva_11_0[0]) | mux_tmp_616;
  assign mux_618_nl = MUX_s_1_2_2(nand_232_cse, or_1345_nl, fsm_output[2]);
  assign mux_622_nl = MUX_s_1_2_2(mux_621_nl, mux_618_nl, fsm_output[8]);
  assign nand_214_nl = ~((fsm_output[4]) & not_tmp_214);
  assign mux_614_nl = MUX_s_1_2_2(nand_214_nl, or_1379_cse, fsm_output[2]);
  assign mux_610_nl = MUX_s_1_2_2(or_277_cse, mux_tmp_609, fsm_output[6]);
  assign or_1349_nl = (fsm_output[4]) | mux_610_nl;
  assign mux_612_nl = MUX_s_1_2_2(mux_477_cse, or_1349_nl, fsm_output[2]);
  assign mux_615_nl = MUX_s_1_2_2(mux_614_nl, mux_612_nl, fsm_output[8]);
  assign mux_623_nl = MUX_s_1_2_2(mux_622_nl, mux_615_nl, fsm_output[1]);
  assign nor_128_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b100));
  assign mux_627_nl = MUX_s_1_2_2(mux_626_nl, mux_623_nl, nor_128_nl);
  assign vec_rsc_0_4_i_wea_d_pff = ~(mux_627_nl | (fsm_output[0]));
  assign nor_492_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_6_12_1[2:0]!=3'b100) |
      (fsm_output[4]) | not_tmp_171);
  assign nor_493_nl = ~((z_out_6_12_1[2:0]!=3'b100) | (fsm_output[7:3]!=5'b01110));
  assign mux_639_nl = MUX_s_1_2_2(nor_492_nl, nor_493_nl, fsm_output[9]);
  assign nor_494_nl = ~((z_out_6_12_1[2:0]!=3'b100) | (~ (fsm_output[9])) | (~ (fsm_output[6]))
      | (fsm_output[5]) | not_tmp_170);
  assign mux_640_nl = MUX_s_1_2_2(mux_639_nl, nor_494_nl, fsm_output[1]);
  assign nor_495_nl = ~((z_out_6_12_1[2:0]!=3'b100) | (fsm_output[7:3]!=5'b01011));
  assign nor_496_nl = ~((z_out_6_12_1[2:0]!=3'b100) | (fsm_output[7:3]!=5'b00000));
  assign mux_638_nl = MUX_s_1_2_2(nor_495_nl, nor_496_nl, fsm_output[9]);
  assign and_349_nl = (fsm_output[1]) & mux_638_nl;
  assign mux_641_nl = MUX_s_1_2_2(mux_640_nl, and_349_nl, fsm_output[2]);
  assign nor_497_nl = ~((z_out_6_12_1[2:0]!=3'b100) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[3])
      | (fsm_output[7]));
  assign or_538_nl = (z_out_6_12_1[2:0]!=3'b100) | (fsm_output[6:5]!=2'b00) | not_tmp_170;
  assign or_536_nl = (z_out_6_12_1[2:0]!=3'b100) | (fsm_output[7:3]!=5'b01000);
  assign mux_636_nl = MUX_s_1_2_2(or_538_nl, or_536_nl, fsm_output[9]);
  assign nor_498_nl = ~((fsm_output[1]) | mux_636_nl);
  assign mux_637_nl = MUX_s_1_2_2(nor_497_nl, nor_498_nl, fsm_output[2]);
  assign mux_642_nl = MUX_s_1_2_2(mux_641_nl, mux_637_nl, fsm_output[8]);
  assign nor_499_nl = ~((VEC_LOOP_j_sva_11_0[2:1]!=2'b10) | (~ (fsm_output[1])) |
      (fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[7:3]!=5'b00110));
  assign nor_500_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b100) | (fsm_output[6:5]!=2'b00)
      | not_tmp_170);
  assign nor_501_nl = ~((COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b100) | (fsm_output[7:3]!=5'b01000));
  assign mux_632_nl = MUX_s_1_2_2(nor_500_nl, nor_501_nl, fsm_output[9]);
  assign nor_502_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10) | (~ (fsm_output[9]))
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[6:4]!=3'b010) | not_tmp_171);
  assign mux_633_nl = MUX_s_1_2_2(mux_632_nl, nor_502_nl, fsm_output[1]);
  assign and_350_nl = COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & mux_633_nl;
  assign mux_634_nl = MUX_s_1_2_2(nor_499_nl, and_350_nl, fsm_output[2]);
  assign nor_503_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | mux_tmp_628);
  assign mux_629_nl = MUX_s_1_2_2(nor_503_nl, nor_624_cse, fsm_output[1]);
  assign nor_505_nl = ~((fsm_output[1]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | mux_tmp_628);
  assign mux_630_nl = MUX_s_1_2_2(mux_629_nl, nor_505_nl, or_521_cse);
  assign nor_506_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10)
      | (~ (fsm_output[1])) | (fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[7:3]!=5'b00000));
  assign mux_631_nl = MUX_s_1_2_2(mux_630_nl, nor_506_nl, fsm_output[2]);
  assign mux_635_nl = MUX_s_1_2_2(mux_634_nl, mux_631_nl, fsm_output[8]);
  assign vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_642_nl,
      mux_635_nl, fsm_output[0]);
  assign or_1330_nl = (fsm_output[2]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | mux_tmp_620;
  assign nand_207_nl = ~((fsm_output[2]) & (VEC_LOOP_j_sva_11_0[0]) & not_tmp_226);
  assign mux_660_nl = MUX_s_1_2_2(or_1330_nl, nand_207_nl, fsm_output[8]);
  assign nand_208_nl = ~(nor_265_cse & not_tmp_225);
  assign or_1331_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | mux_tmp_644;
  assign mux_659_nl = MUX_s_1_2_2(nand_208_nl, or_1331_nl, fsm_output[8]);
  assign mux_661_nl = MUX_s_1_2_2(mux_660_nl, mux_659_nl, fsm_output[1]);
  assign or_1332_nl = (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | mux_tmp_620;
  assign mux_656_nl = MUX_s_1_2_2(or_1332_nl, mux_483_cse, fsm_output[2]);
  assign nand_210_nl = ~((VEC_LOOP_j_sva_11_0[0]) & not_tmp_226);
  assign mux_653_nl = MUX_s_1_2_2(nand_232_cse, nand_210_nl, fsm_output[2]);
  assign mux_657_nl = MUX_s_1_2_2(mux_656_nl, mux_653_nl, fsm_output[8]);
  assign nand_211_nl = ~((fsm_output[4]) & not_tmp_225);
  assign mux_649_nl = MUX_s_1_2_2(nand_211_nl, or_1379_cse, fsm_output[2]);
  assign mux_645_nl = MUX_s_1_2_2(or_277_cse, mux_tmp_644, fsm_output[6]);
  assign or_1338_nl = (fsm_output[4]) | mux_645_nl;
  assign mux_647_nl = MUX_s_1_2_2(mux_477_cse, or_1338_nl, fsm_output[2]);
  assign mux_650_nl = MUX_s_1_2_2(mux_649_nl, mux_647_nl, fsm_output[8]);
  assign mux_658_nl = MUX_s_1_2_2(mux_657_nl, mux_650_nl, fsm_output[1]);
  assign nor_135_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b101));
  assign mux_662_nl = MUX_s_1_2_2(mux_661_nl, mux_658_nl, nor_135_nl);
  assign vec_rsc_0_5_i_wea_d_pff = ~(mux_662_nl | (fsm_output[0]));
  assign nor_462_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_6_12_1[2:0]!=3'b101) |
      (fsm_output[4]) | not_tmp_171);
  assign nor_463_nl = ~((z_out_6_12_1[2:0]!=3'b101) | (fsm_output[7:3]!=5'b01110));
  assign mux_674_nl = MUX_s_1_2_2(nor_462_nl, nor_463_nl, fsm_output[9]);
  assign nor_464_nl = ~((z_out_6_12_1[2:0]!=3'b101) | (~ (fsm_output[9])) | (~ (fsm_output[6]))
      | (fsm_output[5]) | not_tmp_170);
  assign mux_675_nl = MUX_s_1_2_2(mux_674_nl, nor_464_nl, fsm_output[1]);
  assign nor_465_nl = ~((z_out_6_12_1[2:0]!=3'b101) | (fsm_output[7:3]!=5'b01011));
  assign nor_466_nl = ~((z_out_6_12_1[2:0]!=3'b101) | (fsm_output[7:3]!=5'b00000));
  assign mux_673_nl = MUX_s_1_2_2(nor_465_nl, nor_466_nl, fsm_output[9]);
  assign and_342_nl = (fsm_output[1]) & mux_673_nl;
  assign mux_676_nl = MUX_s_1_2_2(mux_675_nl, and_342_nl, fsm_output[2]);
  assign nor_467_nl = ~((z_out_6_12_1[2:0]!=3'b101) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[3])
      | (fsm_output[7]));
  assign or_595_nl = (z_out_6_12_1[2:0]!=3'b101) | (fsm_output[6:5]!=2'b00) | not_tmp_170;
  assign or_593_nl = (z_out_6_12_1[2:0]!=3'b101) | (fsm_output[7:3]!=5'b01000);
  assign mux_671_nl = MUX_s_1_2_2(or_595_nl, or_593_nl, fsm_output[9]);
  assign nor_468_nl = ~((fsm_output[1]) | mux_671_nl);
  assign mux_672_nl = MUX_s_1_2_2(nor_467_nl, nor_468_nl, fsm_output[2]);
  assign mux_677_nl = MUX_s_1_2_2(mux_676_nl, mux_672_nl, fsm_output[8]);
  assign nor_469_nl = ~((VEC_LOOP_j_sva_11_0[2:1]!=2'b10) | (~ (fsm_output[1])) |
      (fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b00110));
  assign nor_470_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b101) | (fsm_output[6:5]!=2'b00)
      | not_tmp_170);
  assign nor_471_nl = ~((COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b101) | (fsm_output[7:3]!=5'b01000));
  assign mux_667_nl = MUX_s_1_2_2(nor_470_nl, nor_471_nl, fsm_output[9]);
  assign nor_472_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b10) | (~ (fsm_output[9]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[6:4]!=3'b010) | not_tmp_171);
  assign mux_668_nl = MUX_s_1_2_2(mux_667_nl, nor_472_nl, fsm_output[1]);
  assign and_343_nl = COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & mux_668_nl;
  assign mux_669_nl = MUX_s_1_2_2(nor_469_nl, and_343_nl, fsm_output[2]);
  assign nor_473_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | mux_tmp_663);
  assign mux_664_nl = MUX_s_1_2_2(nor_473_nl, nor_594_cse, fsm_output[1]);
  assign nor_475_nl = ~((fsm_output[1]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | mux_tmp_663);
  assign mux_665_nl = MUX_s_1_2_2(mux_664_nl, nor_475_nl, or_521_cse);
  assign nor_476_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b10)
      | (~ (fsm_output[1])) | (fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b00000));
  assign mux_666_nl = MUX_s_1_2_2(mux_665_nl, nor_476_nl, fsm_output[2]);
  assign mux_670_nl = MUX_s_1_2_2(mux_669_nl, mux_666_nl, fsm_output[8]);
  assign vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_677_nl,
      mux_670_nl, fsm_output[0]);
  assign nand_202_nl = ~(nor_112_cse & not_tmp_239);
  assign or_1321_nl = (~ (fsm_output[2])) | (VEC_LOOP_j_sva_11_0[0]) | mux_tmp_686;
  assign mux_695_nl = MUX_s_1_2_2(nand_202_nl, or_1321_nl, fsm_output[8]);
  assign nand_203_nl = ~(nor_265_cse & not_tmp_237);
  assign or_1322_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | mux_tmp_679;
  assign mux_694_nl = MUX_s_1_2_2(nand_203_nl, or_1322_nl, fsm_output[8]);
  assign mux_696_nl = MUX_s_1_2_2(mux_695_nl, mux_694_nl, fsm_output[1]);
  assign nand_204_nl = ~(nor_114_cse & not_tmp_239);
  assign mux_691_nl = MUX_s_1_2_2(nand_204_nl, mux_483_cse, fsm_output[2]);
  assign or_1325_nl = (VEC_LOOP_j_sva_11_0[0]) | mux_tmp_686;
  assign mux_688_nl = MUX_s_1_2_2(nand_232_cse, or_1325_nl, fsm_output[2]);
  assign mux_692_nl = MUX_s_1_2_2(mux_691_nl, mux_688_nl, fsm_output[8]);
  assign nand_206_nl = ~((fsm_output[4]) & not_tmp_237);
  assign mux_684_nl = MUX_s_1_2_2(nand_206_nl, or_1379_cse, fsm_output[2]);
  assign mux_680_nl = MUX_s_1_2_2(or_277_cse, mux_tmp_679, fsm_output[6]);
  assign or_1329_nl = (fsm_output[4]) | mux_680_nl;
  assign mux_682_nl = MUX_s_1_2_2(mux_477_cse, or_1329_nl, fsm_output[2]);
  assign mux_685_nl = MUX_s_1_2_2(mux_684_nl, mux_682_nl, fsm_output[8]);
  assign mux_693_nl = MUX_s_1_2_2(mux_692_nl, mux_685_nl, fsm_output[1]);
  assign nor_143_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b110));
  assign mux_697_nl = MUX_s_1_2_2(mux_696_nl, mux_693_nl, nor_143_nl);
  assign vec_rsc_0_6_i_wea_d_pff = ~(mux_697_nl | (fsm_output[0]));
  assign nor_432_nl = ~((fsm_output[6:5]!=2'b10) | (z_out_6_12_1[2:0]!=3'b110) |
      (fsm_output[4]) | not_tmp_171);
  assign nor_433_nl = ~((z_out_6_12_1[2:0]!=3'b110) | (fsm_output[7:3]!=5'b01110));
  assign mux_709_nl = MUX_s_1_2_2(nor_432_nl, nor_433_nl, fsm_output[9]);
  assign nor_434_nl = ~((z_out_6_12_1[2:0]!=3'b110) | (~ (fsm_output[9])) | (~ (fsm_output[6]))
      | (fsm_output[5]) | not_tmp_170);
  assign mux_710_nl = MUX_s_1_2_2(mux_709_nl, nor_434_nl, fsm_output[1]);
  assign nor_435_nl = ~((z_out_6_12_1[2:0]!=3'b110) | (fsm_output[7:3]!=5'b01011));
  assign nor_436_nl = ~((z_out_6_12_1[2:0]!=3'b110) | (fsm_output[7:3]!=5'b00000));
  assign mux_708_nl = MUX_s_1_2_2(nor_435_nl, nor_436_nl, fsm_output[9]);
  assign and_334_nl = (fsm_output[1]) & mux_708_nl;
  assign mux_711_nl = MUX_s_1_2_2(mux_710_nl, and_334_nl, fsm_output[2]);
  assign nor_437_nl = ~((z_out_6_12_1[2:0]!=3'b110) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[5])) | (~ (fsm_output[4])) | (fsm_output[3])
      | (fsm_output[7]));
  assign or_650_nl = (z_out_6_12_1[2:0]!=3'b110) | (fsm_output[6:5]!=2'b00) | not_tmp_170;
  assign or_648_nl = (z_out_6_12_1[2:0]!=3'b110) | (fsm_output[7:3]!=5'b01000);
  assign mux_706_nl = MUX_s_1_2_2(or_650_nl, or_648_nl, fsm_output[9]);
  assign nor_438_nl = ~((fsm_output[1]) | mux_706_nl);
  assign mux_707_nl = MUX_s_1_2_2(nor_437_nl, nor_438_nl, fsm_output[2]);
  assign mux_712_nl = MUX_s_1_2_2(mux_711_nl, mux_707_nl, fsm_output[8]);
  assign nor_439_nl = ~((VEC_LOOP_j_sva_11_0[2:1]!=2'b11) | (~ (fsm_output[1])) |
      (fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[7:3]!=5'b00110));
  assign nor_440_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b110) | (fsm_output[6:5]!=2'b00)
      | not_tmp_170);
  assign nor_441_nl = ~((COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b110) | (fsm_output[7:3]!=5'b01000));
  assign mux_702_nl = MUX_s_1_2_2(nor_440_nl, nor_441_nl, fsm_output[9]);
  assign nor_442_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b11) | (~ (fsm_output[9]))
      | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[6:4]!=3'b010) | not_tmp_171);
  assign mux_703_nl = MUX_s_1_2_2(mux_702_nl, nor_442_nl, fsm_output[1]);
  assign and_335_nl = COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & mux_703_nl;
  assign mux_704_nl = MUX_s_1_2_2(nor_439_nl, and_335_nl, fsm_output[2]);
  assign nor_443_nl = ~((fsm_output[1]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | mux_tmp_698);
  assign nor_444_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | mux_tmp_698);
  assign mux_699_nl = MUX_s_1_2_2(nor_444_nl, nor_624_cse, fsm_output[1]);
  assign mux_700_nl = MUX_s_1_2_2(nor_443_nl, mux_699_nl, and_336_cse);
  assign nor_446_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b11)
      | (~ (fsm_output[1])) | (fsm_output[9]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[7:3]!=5'b00000));
  assign mux_701_nl = MUX_s_1_2_2(mux_700_nl, nor_446_nl, fsm_output[2]);
  assign mux_705_nl = MUX_s_1_2_2(mux_704_nl, mux_701_nl, fsm_output[8]);
  assign vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_712_nl,
      mux_705_nl, fsm_output[0]);
  assign nand_195_nl = ~(nor_122_cse & not_tmp_239);
  assign nand_196_nl = ~((fsm_output[2]) & (VEC_LOOP_j_sva_11_0[0]) & not_tmp_250);
  assign mux_730_nl = MUX_s_1_2_2(nand_195_nl, nand_196_nl, fsm_output[8]);
  assign nand_197_nl = ~(nor_265_cse & not_tmp_249);
  assign or_1314_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | mux_tmp_714;
  assign mux_729_nl = MUX_s_1_2_2(nand_197_nl, or_1314_nl, fsm_output[8]);
  assign mux_731_nl = MUX_s_1_2_2(mux_730_nl, mux_729_nl, fsm_output[1]);
  assign nand_198_nl = ~((VEC_LOOP_j_sva_11_0[1:0]==2'b11) & not_tmp_239);
  assign mux_726_nl = MUX_s_1_2_2(nand_198_nl, mux_483_cse, fsm_output[2]);
  assign nand_200_nl = ~((VEC_LOOP_j_sva_11_0[0]) & not_tmp_250);
  assign mux_723_nl = MUX_s_1_2_2(nand_232_cse, nand_200_nl, fsm_output[2]);
  assign mux_727_nl = MUX_s_1_2_2(mux_726_nl, mux_723_nl, fsm_output[8]);
  assign nand_201_nl = ~((fsm_output[4]) & not_tmp_249);
  assign mux_719_nl = MUX_s_1_2_2(nand_201_nl, or_1379_cse, fsm_output[2]);
  assign mux_715_nl = MUX_s_1_2_2(or_277_cse, mux_tmp_714, fsm_output[6]);
  assign or_1320_nl = (fsm_output[4]) | mux_715_nl;
  assign mux_717_nl = MUX_s_1_2_2(mux_477_cse, or_1320_nl, fsm_output[2]);
  assign mux_720_nl = MUX_s_1_2_2(mux_719_nl, mux_717_nl, fsm_output[8]);
  assign mux_728_nl = MUX_s_1_2_2(mux_727_nl, mux_720_nl, fsm_output[1]);
  assign and_333_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b111);
  assign mux_732_nl = MUX_s_1_2_2(mux_731_nl, mux_728_nl, and_333_nl);
  assign vec_rsc_0_7_i_wea_d_pff = ~(mux_732_nl | (fsm_output[0]));
  assign nor_404_nl = ~((z_out_6_12_1[2:0]!=3'b111) | (fsm_output[6:4]!=3'b100) |
      not_tmp_171);
  assign and_321_nl = (z_out_6_12_1[2:0]==3'b111) & (fsm_output[7:3]==5'b01110);
  assign mux_744_nl = MUX_s_1_2_2(nor_404_nl, and_321_nl, fsm_output[9]);
  assign nor_405_nl = ~((~((z_out_6_12_1[2:0]==3'b111) & (fsm_output[9]) & (fsm_output[6])
      & (fsm_output[4]) & (~ (fsm_output[5])))) | not_tmp_171);
  assign mux_745_nl = MUX_s_1_2_2(mux_744_nl, nor_405_nl, fsm_output[1]);
  assign and_323_nl = (z_out_6_12_1[2:0]==3'b111) & (fsm_output[7:3]==5'b01011);
  assign nor_406_nl = ~((z_out_6_12_1[2:0]!=3'b111) | (fsm_output[7:3]!=5'b00000));
  assign mux_743_nl = MUX_s_1_2_2(and_323_nl, nor_406_nl, fsm_output[9]);
  assign and_322_nl = (fsm_output[1]) & mux_743_nl;
  assign mux_746_nl = MUX_s_1_2_2(mux_745_nl, and_322_nl, fsm_output[2]);
  assign nor_407_nl = ~((z_out_6_12_1[2:0]!=3'b111) | (~ (fsm_output[1])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[4])) | (~ (fsm_output[5])) | (fsm_output[3])
      | (fsm_output[7]));
  assign or_702_nl = (z_out_6_12_1[2:0]!=3'b111) | (fsm_output[6:4]!=3'b001) | not_tmp_171;
  assign or_700_nl = (z_out_6_12_1[2:0]!=3'b111) | (fsm_output[7:3]!=5'b01000);
  assign mux_741_nl = MUX_s_1_2_2(or_702_nl, or_700_nl, fsm_output[9]);
  assign nor_408_nl = ~((fsm_output[1]) | mux_741_nl);
  assign mux_742_nl = MUX_s_1_2_2(nor_407_nl, nor_408_nl, fsm_output[2]);
  assign mux_747_nl = MUX_s_1_2_2(mux_746_nl, mux_742_nl, fsm_output[8]);
  assign nor_409_nl = ~((VEC_LOOP_j_sva_11_0[2:1]!=2'b11) | (~ (fsm_output[1])) |
      (fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b00110));
  assign nor_410_nl = ~((COMP_LOOP_acc_1_cse_2_sva[2:0]!=3'b111) | (fsm_output[6:4]!=3'b001)
      | not_tmp_171);
  assign nor_411_nl = ~((COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b111) | (fsm_output[7:3]!=5'b01000));
  assign mux_737_nl = MUX_s_1_2_2(nor_410_nl, nor_411_nl, fsm_output[9]);
  assign nor_412_nl = ~((COMP_LOOP_acc_14_psp_sva[1:0]!=2'b11) | (~ (fsm_output[9]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b10101));
  assign mux_738_nl = MUX_s_1_2_2(mux_737_nl, nor_412_nl, fsm_output[1]);
  assign and_324_nl = COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & mux_738_nl;
  assign mux_739_nl = MUX_s_1_2_2(nor_409_nl, and_324_nl, fsm_output[2]);
  assign nor_413_nl = ~((fsm_output[1]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | mux_tmp_733);
  assign nor_414_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | mux_tmp_733);
  assign nor_415_nl = ~((fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[6:4]!=3'b101)
      | not_tmp_171);
  assign mux_734_nl = MUX_s_1_2_2(nor_414_nl, nor_415_nl, fsm_output[1]);
  assign mux_735_nl = MUX_s_1_2_2(nor_413_nl, mux_734_nl, and_336_cse);
  assign nor_416_nl = ~((~ COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_sva[1:0]!=2'b11)
      | (~ (fsm_output[1])) | (fsm_output[9]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[7:3]!=5'b00000));
  assign mux_736_nl = MUX_s_1_2_2(mux_735_nl, nor_416_nl, fsm_output[2]);
  assign mux_740_nl = MUX_s_1_2_2(mux_739_nl, mux_736_nl, fsm_output[8]);
  assign vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_747_nl,
      mux_740_nl, fsm_output[0]);
  assign and_dcpl_218 = (fsm_output[3]) & (~ (fsm_output[5])) & (~ (fsm_output[2]));
  assign and_dcpl_223 = nor_692_cse & (fsm_output[1]) & (~ (fsm_output[6]));
  assign or_1409_nl = (~((fsm_output[9]) & (fsm_output[1]) & (fsm_output[2]) & (~
      (fsm_output[8])))) | nand_240_cse;
  assign or_1407_nl = (fsm_output[9]) | (fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[8]))
      | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_1417_nl = MUX_s_1_2_2(or_1409_nl, or_1407_nl, fsm_output[3]);
  assign nor_789_nl = ~((fsm_output[5]) | mux_1417_nl);
  assign and_709_nl = (fsm_output[3]) & (fsm_output[9]) & (fsm_output[1]) & (~ (fsm_output[2]))
      & (fsm_output[8]) & (fsm_output[0]) & (~ (fsm_output[6]));
  assign and_711_nl = (fsm_output[8]) & (fsm_output[0]) & (fsm_output[6]);
  assign nor_790_nl = ~((fsm_output[8]) | (fsm_output[0]) | (fsm_output[6]));
  assign mux_1415_nl = MUX_s_1_2_2(and_711_nl, nor_790_nl, fsm_output[2]);
  assign and_710_nl = (~((fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[1]))))
      & mux_1415_nl;
  assign mux_1416_nl = MUX_s_1_2_2(and_709_nl, and_710_nl, fsm_output[5]);
  assign mux_1418_nl = MUX_s_1_2_2(nor_789_nl, mux_1416_nl, fsm_output[4]);
  assign nand_259_nl = ~((fsm_output[2]) & (fsm_output[8]) & (fsm_output[0]) & (fsm_output[6]));
  assign or_1403_nl = (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | (fsm_output[6]);
  assign mux_1444_nl = MUX_s_1_2_2(nand_259_nl, or_1403_nl, fsm_output[1]);
  assign nor_791_nl = ~((~ (fsm_output[3])) | (fsm_output[9]) | mux_1444_nl);
  assign nor_792_nl = ~((fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[1]) |
      (fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[0])) | (fsm_output[6]));
  assign mux_1414_nl = MUX_s_1_2_2(nor_791_nl, nor_792_nl, fsm_output[5]);
  assign and_712_nl = (fsm_output[4]) & mux_1414_nl;
  assign not_tmp_519 = MUX_s_1_2_2(mux_1418_nl, and_712_nl, fsm_output[7]);
  assign mux_tmp_1422 = MUX_s_1_2_2(or_718_cse, or_tmp_677, fsm_output[6]);
  assign mux_tmp_1425 = MUX_s_1_2_2(or_tmp_682, or_718_cse, fsm_output[6]);
  assign nor_784_nl = ~((~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[9]))
      | (~ (fsm_output[1])) | (~ (fsm_output[6])) | (~ (fsm_output[8])) | (fsm_output[0])
      | (fsm_output[7]));
  assign nand_249_nl = ~((fsm_output[1]) & (~ mux_tmp_1425));
  assign or_1425_nl = (fsm_output[1]) | (fsm_output[8]) | (fsm_output[0]) | (fsm_output[7]);
  assign mux_1427_nl = MUX_s_1_2_2(nand_249_nl, or_1425_nl, fsm_output[9]);
  assign nor_785_nl = ~((fsm_output[4]) | mux_1427_nl);
  assign and_713_nl = (fsm_output[1]) & (fsm_output[8]) & (~ (fsm_output[0])) & (fsm_output[7]);
  assign nor_787_nl = ~((fsm_output[1]) | mux_tmp_1425);
  assign mux_1426_nl = MUX_s_1_2_2(and_713_nl, nor_787_nl, fsm_output[9]);
  assign and_708_nl = (fsm_output[4]) & mux_1426_nl;
  assign mux_1428_nl = MUX_s_1_2_2(nor_785_nl, and_708_nl, fsm_output[2]);
  assign mux_1429_nl = MUX_s_1_2_2(nor_784_nl, mux_1428_nl, fsm_output[3]);
  assign or_1420_nl = (fsm_output[9]) | (fsm_output[1]) | mux_tmp_1422;
  assign nand_247_nl = ~((fsm_output[9]) & (fsm_output[1]) & (~ mux_tmp_1422));
  assign mux_1423_nl = MUX_s_1_2_2(or_1420_nl, nand_247_nl, fsm_output[4]);
  assign mux_1420_nl = MUX_s_1_2_2(or_tmp_9, or_730_cse, fsm_output[8]);
  assign mux_1421_nl = MUX_s_1_2_2(mux_1420_nl, or_tmp_682, fsm_output[6]);
  assign or_1415_nl = (~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[1]) | mux_1421_nl;
  assign mux_1424_nl = MUX_s_1_2_2(mux_1423_nl, or_1415_nl, fsm_output[2]);
  assign nor_788_nl = ~((fsm_output[3]) | mux_1424_nl);
  assign not_tmp_524 = MUX_s_1_2_2(mux_1429_nl, nor_788_nl, fsm_output[5]);
  assign or_1456_nl = (~ (fsm_output[9])) | (fsm_output[6]) | (fsm_output[8]) | (~
      (fsm_output[2]));
  assign nand_nl = ~((fsm_output[9]) & (fsm_output[6]) & (fsm_output[8]) & (~ (fsm_output[2])));
  assign mux_1433_nl = MUX_s_1_2_2(or_1456_nl, nand_nl, fsm_output[1]);
  assign or_1457_nl = (~ (fsm_output[1])) | (fsm_output[9]) | (~ (fsm_output[6]))
      | (fsm_output[8]) | (~ (fsm_output[2]));
  assign mux_1434_nl = MUX_s_1_2_2(mux_1433_nl, or_1457_nl, fsm_output[7]);
  assign mux_1435_nl = MUX_s_1_2_2(or_798_cse, mux_1434_nl, fsm_output[4]);
  assign mux_1436_nl = MUX_s_1_2_2(or_1312_cse, mux_1435_nl, fsm_output[3]);
  assign nor_775_nl = ~((fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[6])) |
      (fsm_output[8]) | (~ (fsm_output[2])));
  assign nor_776_nl = ~((~ (fsm_output[9])) | (~ (fsm_output[6])) | (fsm_output[8])
      | (fsm_output[2]));
  assign nor_777_nl = ~((fsm_output[9]) | (fsm_output[6]) | (~ (fsm_output[8])) |
      (fsm_output[2]));
  assign mux_1431_nl = MUX_s_1_2_2(nor_776_nl, nor_777_nl, fsm_output[1]);
  assign mux_1432_nl = MUX_s_1_2_2(nor_775_nl, mux_1431_nl, fsm_output[7]);
  assign nand_256_nl = ~((~((fsm_output[4:3]!=2'b10))) & mux_1432_nl);
  assign mux_1437_nl = MUX_s_1_2_2(mux_1436_nl, nand_256_nl, fsm_output[5]);
  assign and_dcpl_246 = ~(mux_1437_nl | (fsm_output[0]));
  assign nor_tmp_272 = (fsm_output[1]) & (fsm_output[4]);
  assign nor_780_nl = ~((fsm_output[1]) | (fsm_output[4]));
  assign mux_1440_nl = MUX_s_1_2_2(nor_780_nl, nor_tmp_272, fsm_output[9]);
  assign nor_779_nl = ~((fsm_output[7:6]!=2'b00) | (~((fsm_output[8]) & mux_1440_nl)));
  assign nor_781_nl = ~((fsm_output[9:8]!=2'b00) | (~ nor_tmp_272));
  assign nor_782_nl = ~((~ (fsm_output[8])) | (fsm_output[9]) | (fsm_output[1]) |
      (~ (fsm_output[4])));
  assign mux_1439_nl = MUX_s_1_2_2(nor_781_nl, nor_782_nl, fsm_output[6]);
  assign and_nl = (fsm_output[7]) & mux_1439_nl;
  assign mux_1441_nl = MUX_s_1_2_2(nor_779_nl, and_nl, fsm_output[2]);
  assign mux_1442_nl = MUX_s_1_2_2(nor_365_cse, mux_1441_nl, fsm_output[3]);
  assign nand_262_nl = ~((fsm_output[6]) & (fsm_output[8]) & (~ (fsm_output[9]))
      & nor_tmp_272);
  assign or_1442_nl = (fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[9])) | (fsm_output[1])
      | (~ (fsm_output[4]));
  assign mux_1438_nl = MUX_s_1_2_2(nand_262_nl, or_1442_nl, fsm_output[7]);
  assign nor_783_nl = ~((fsm_output[3:2]!=2'b00) | mux_1438_nl);
  assign mux_1443_nl = MUX_s_1_2_2(mux_1442_nl, nor_783_nl, fsm_output[5]);
  assign and_dcpl_247 = mux_1443_nl & (fsm_output[0]);
  assign and_dcpl_248 = (~ (fsm_output[6])) & (fsm_output[0]);
  assign and_dcpl_256 = nor_692_cse & (fsm_output[5:1]==5'b00000) & and_dcpl_248;
  assign and_dcpl_262 = nor_692_cse & (fsm_output[5:1]==5'b11010) & and_dcpl_248;
  assign and_dcpl_265 = (~ (fsm_output[2])) & (fsm_output[4]) & (fsm_output[1]);
  assign and_dcpl_267 = (~ (fsm_output[3])) & (fsm_output[5]);
  assign and_dcpl_271 = nor_692_cse & and_dcpl_267 & and_dcpl_265 & (~ (fsm_output[6]))
      & (fsm_output[0]);
  assign and_dcpl_277 = (fsm_output[9:7]==3'b010) & and_dcpl_267 & and_dcpl_265 &
      (~ (fsm_output[6])) & (~ (fsm_output[0]));
  assign and_dcpl_278 = (fsm_output[6]) & (~ (fsm_output[0]));
  assign and_dcpl_280 = (fsm_output[3]) & (~ (fsm_output[5]));
  assign and_dcpl_284 = (fsm_output[9:7]==3'b101) & and_dcpl_280 & and_dcpl_265 &
      and_dcpl_278;
  assign and_dcpl_289 = nor_692_cse & and_dcpl_280 & (fsm_output[2]) & (fsm_output[4])
      & (fsm_output[1]) & and_dcpl_278;
  assign and_dcpl_291 = (~ (fsm_output[2])) & (fsm_output[4]);
  assign and_dcpl_298 = nor_692_cse & and_dcpl_267 & and_dcpl_291 & (fsm_output[1])
      & (~ (fsm_output[6])) & (fsm_output[0]);
  assign and_dcpl_300 = (fsm_output[2]) & (fsm_output[4]);
  assign and_dcpl_305 = nor_692_cse & and_dcpl_280 & and_dcpl_300 & (fsm_output[1])
      & and_dcpl_278;
  assign and_dcpl_309 = (fsm_output[7]) & (~ (fsm_output[9]));
  assign and_dcpl_312 = and_dcpl_309 & (~ (fsm_output[8])) & and_dcpl_280 & (~ (fsm_output[2]))
      & (~ (fsm_output[4])) & (~ (fsm_output[1])) & and_dcpl_278;
  assign and_dcpl_313 = ~((fsm_output[6]) | (fsm_output[0]));
  assign and_dcpl_318 = and_dcpl_309 & (fsm_output[8]) & and_dcpl_280 & and_dcpl_300
      & (~ (fsm_output[1])) & and_dcpl_313;
  assign and_dcpl_324 = (fsm_output[9:7]==3'b100);
  assign and_dcpl_326 = and_dcpl_324 & (fsm_output[5:1]==5'b00011) & and_dcpl_313;
  assign and_dcpl_330 = and_dcpl_324 & and_dcpl_267 & and_dcpl_291 & (~ (fsm_output[1]))
      & and_dcpl_278;
  assign and_dcpl_342 = and_dcpl_291 & (fsm_output[1]);
  assign and_dcpl_355 = (fsm_output[2]) & (~ (fsm_output[4]));
  assign nor_797_cse = ~((fsm_output[3]) | (fsm_output[5]));
  assign and_dcpl_359 = (fsm_output[9:8]==2'b10);
  assign and_dcpl_360 = and_dcpl_359 & (~ (fsm_output[7]));
  assign and_dcpl_410 = (~ (fsm_output[7])) & (fsm_output[9]);
  assign and_dcpl_411 = and_dcpl_410 & (~ (fsm_output[8]));
  assign and_dcpl_442 = ~((fsm_output!=10'b0000001001));
  assign and_dcpl_451 = nor_692_cse & (fsm_output[6:0]==7'b0110011);
  assign and_dcpl_460 = (fsm_output==10'b1101000100);
  assign and_dcpl_467 = nor_692_cse & (fsm_output[6:0]==7'b0001010);
  assign and_243_m1c = and_dcpl_76 & and_dcpl_157;
  assign nor_tmp_273 = ((~ (fsm_output[1])) | (fsm_output[9])) & (fsm_output[7]);
  assign mux_tmp_1456 = MUX_s_1_2_2(mux_tmp_898, or_tmp_72, and_303_cse);
  assign or_tmp_1262 = (fsm_output[0]) | (fsm_output[9]);
  assign or_tmp_1267 = (fsm_output[8]) | (fsm_output[0]) | (~ (fsm_output[9]));
  assign or_tmp_1269 = nor_820_cse | (fsm_output[0]) | (fsm_output[9]);
  assign or_tmp_1273 = (~ (fsm_output[6])) | (~ (fsm_output[8])) | (fsm_output[0])
      | (fsm_output[9]);
  assign or_tmp_1274 = (fsm_output[6]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (~ (fsm_output[8])) | (~ (fsm_output[0])) | (fsm_output[9]);
  assign not_tmp_621 = ~((fsm_output[0]) & (fsm_output[9]));
  assign COMP_LOOP_or_39_itm = and_dcpl_247 | and_dcpl_262;
  assign operator_64_false_1_nor_1_itm = ~(and_dcpl_271 | and_dcpl_284 | and_dcpl_289);
  assign COMP_LOOP_or_43_itm = and_dcpl_305 | and_dcpl_312 | and_dcpl_318 | and_dcpl_326
      | and_dcpl_330;
  always @(posedge clk) begin
    if ( mux_453_itm ) begin
      p_sva <= p_rsci_idat;
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_53 & and_dcpl_33 & and_dcpl_50) | STAGE_LOOP_i_3_0_sva_mx0c1 )
        begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, STAGE_LOOP_i_3_0_sva_2, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_7_obj_ld_cse <= 1'b0;
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= 1'b0;
      modExp_exp_1_0_1_sva_1 <= 1'b0;
      modExp_exp_1_7_1_sva <= 1'b0;
      modExp_exp_1_2_1_sva <= 1'b0;
      modExp_exp_1_1_1_sva <= 1'b0;
      COMP_LOOP_COMP_LOOP_nor_1_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_124_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_125_itm <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_7_obj_ld_cse <= and_dcpl_23 & and_dcpl_33 & (fsm_output[7])
          & (~ (fsm_output[1])) & (fsm_output[8]) & (fsm_output[9]) & (fsm_output[0])
          & (~ STAGE_LOOP_acc_itm_2_1);
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= (operator_64_false_1_mux1h_nl & (mux_1171_nl
          | (fsm_output[1:0]!=2'b00))) | (mux_1215_nl & (fsm_output[1:0]==2'b10));
      modExp_exp_1_0_1_sva_1 <= (COMP_LOOP_mux_42_nl & (~(mux_1218_nl & (fsm_output[2])
          & (~ (fsm_output[0]))))) | (~(mux_1266_nl | (fsm_output[2]) | (fsm_output[0])));
      modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_32_nl & (~(mux_1295_nl & (fsm_output[0])));
      modExp_exp_1_2_1_sva <= COMP_LOOP_mux1h_46_nl & (~ and_dcpl_191);
      modExp_exp_1_1_1_sva <= (COMP_LOOP_mux1h_48_nl & (mux_1311_nl | (fsm_output[9])))
          | (~(mux_1314_nl | (fsm_output[0])));
      COMP_LOOP_COMP_LOOP_nor_1_itm <= ~((z_out_6_12_1[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_12_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_12_cse,
          COMP_LOOP_COMP_LOOP_and_11_cse, modExp_while_or_1_cse);
      COMP_LOOP_COMP_LOOP_and_124_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_13_cse,
          COMP_LOOP_COMP_LOOP_and_12_cse, modExp_while_or_1_cse);
      COMP_LOOP_COMP_LOOP_and_125_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_37_cse,
          COMP_LOOP_COMP_LOOP_and_13_cse, modExp_while_or_1_cse);
    end
  end
  always @(posedge clk) begin
    modulo_result_rem_cmp_a <= MUX1HOT_v_64_5_2(z_out, operator_64_false_acc_mut_63_0,
        COMP_LOOP_1_acc_8_itm, COMP_LOOP_1_mul_mut, COMP_LOOP_1_acc_5_mut_mx0w5,
        {modulo_result_or_nl , (~ mux_802_nl) , (~ mux_848_nl) , mux_880_nl , and_dcpl_151});
    modulo_result_rem_cmp_b <= p_sva;
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_2, ({operator_64_false_acc_mut_64
        , operator_64_false_acc_mut_63_0}), and_dcpl_156);
    operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_156);
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_446_cse, mux_444_nl, fsm_output[0]) ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_1493_nl ) begin
      operator_64_false_acc_mut_64 <= operator_64_false_operator_64_false_mux_rgt[64];
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_1519_nl, mux_1503_nl, fsm_output[5]) ) begin
      operator_64_false_acc_mut_63_0 <= operator_64_false_operator_64_false_mux_rgt[63:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_sva_11_0 <= 12'b000000000000;
    end
    else if ( (~(mux_tmp_1013 | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[7])
        | (~ not_tmp_82))) | VEC_LOOP_j_sva_11_0_mx0c1 ) begin
      VEC_LOOP_j_sva_11_0 <= MUX_v_12_2_2(12'b000000000000, (z_out_1[11:0]), VEC_LOOP_j_sva_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_k_9_3_sva_5_0 <= 6'b000000;
    end
    else if ( MUX_s_1_2_2(mux_1522_nl, nor_827_nl, fsm_output[6]) ) begin
      COMP_LOOP_k_9_3_sva_5_0 <= MUX_v_6_2_2(6'b000000, (z_out_8[5:0]), or_1460_nl);
    end
  end
  always @(posedge clk) begin
    if ( (operator_64_false_slc_modExp_exp_0_1_itm | modExp_result_sva_mx0c0 | (~
        mux_1035_nl)) & (modExp_result_sva_mx0c0 | modExp_result_and_rgt | modExp_result_and_1_rgt)
        ) begin
      modExp_result_sva <= MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modulo_result_rem_cmp_z, modulo_qr_sva_1_mx1w1, {modExp_result_sva_mx0c0
          , modExp_result_and_rgt , modExp_result_and_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_82 & and_dcpl_157) | modExp_base_sva_mx0c1 ) begin
      modExp_base_sva <= MUX_v_64_2_2(r_sva, modulo_result_mux_1_cse, modExp_base_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_64_false_slc_modExp_exp_0_1_itm <= 1'b0;
    end
    else if ( (~(mux_tmp_1013 | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[7])
        | (fsm_output[8]) | (fsm_output[9]))) & or_dcpl_3 ) begin
      operator_64_false_slc_modExp_exp_0_1_itm <= MUX_s_1_2_2((operator_66_true_div_cmp_z[0]),
          (modExp_exp_sva_rsp_1[0]), or_dcpl_56);
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_3 ) begin
      operator_64_false_slc_modExp_exp_63_1_itm <= operator_64_false_slc_modExp_exp_63_1_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_11_itm <= 1'b0;
    end
    else if ( and_dcpl_150 | and_dcpl_177 | and_dcpl_77 | and_dcpl_90 | and_dcpl_98
        | and_dcpl_104 | and_dcpl_109 | and_dcpl_116 | and_dcpl_126 | and_dcpl_134
        ) begin
      COMP_LOOP_COMP_LOOP_and_11_itm <= MUX1HOT_s_1_4_2((~ (z_out_8[63])), (~ (z_out_2[8])),
          COMP_LOOP_COMP_LOOP_and_11_cse, COMP_LOOP_COMP_LOOP_and_37_cse, {and_dcpl_150
          , and_dcpl_177 , and_dcpl_77 , modExp_while_or_1_cse});
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_82 & and_dcpl_66) | mux_1134_nl | and_dcpl_151 ) begin
      COMP_LOOP_1_acc_8_itm <= MUX_v_64_2_2(z_out, (z_out_2[63:0]), and_dcpl_151);
    end
  end
  always @(posedge clk) begin
    if ( ~(or_dcpl_62 | (~ (fsm_output[5])) | (fsm_output[6]) | (fsm_output[7]) |
        (~ (fsm_output[1])) | (fsm_output[8]) | or_1275_cse) ) begin
      COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_58_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_30_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_32_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_4_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_5_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_6_itm <= 1'b0;
    end
    else if ( mux_1151_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= ~((VEC_LOOP_j_sva_11_0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_58_itm <= (z_out_8[0]) & (VEC_LOOP_j_sva_11_0[0]) &
          (~ (z_out_8[1]));
      COMP_LOOP_COMP_LOOP_and_30_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[2:0]==3'b011);
      COMP_LOOP_COMP_LOOP_and_32_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[2:0]==3'b101);
      COMP_LOOP_COMP_LOOP_and_4_itm <= (VEC_LOOP_j_sva_11_0[2:0]==3'b101);
      COMP_LOOP_COMP_LOOP_and_5_itm <= (VEC_LOOP_j_sva_11_0[2:0]==3'b110);
      COMP_LOOP_COMP_LOOP_and_6_itm <= (VEC_LOOP_j_sva_11_0[2:0]==3'b111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_2_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(nor_808_nl, and_714_nl, fsm_output[8]) ) begin
      COMP_LOOP_COMP_LOOP_and_2_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_2_nl,
          (~ (readslicef_10_1_9(COMP_LOOP_1_acc_nl))), and_dcpl_134);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 11'b00000000000;
    end
    else if ( mux_1157_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_11_psp_sva <= z_out_8[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 12'b000000000000;
    end
    else if ( ~(mux_1160_nl & not_tmp_82) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_4_sva <= 12'b000000000000;
    end
    else if ( mux_1162_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_4_sva <= z_out_1[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_384, or_1038_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_13_psp_sva <= z_out_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_6_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_384, or_1043_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_6_sva <= nl_COMP_LOOP_acc_1_cse_6_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_14_psp_sva <= 11'b00000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_384, and_212_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_14_psp_sva <= z_out_7[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_384, and_214_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_sva <= nl_COMP_LOOP_acc_1_cse_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_6_1_sva <= 1'b0;
      modExp_exp_1_5_1_sva <= 1'b0;
      modExp_exp_1_4_1_sva <= 1'b0;
      modExp_exp_1_3_1_sva <= 1'b0;
    end
    else if ( mux_1289_itm ) begin
      modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[3]), modExp_exp_1_7_1_sva,
          (COMP_LOOP_k_9_3_sva_5_0[4]), {and_dcpl_191 , and_dcpl_194 , and_dcpl_192});
      modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[2]), modExp_exp_1_6_1_sva,
          (COMP_LOOP_k_9_3_sva_5_0[3]), {and_dcpl_191 , and_dcpl_194 , and_dcpl_192});
      modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[1]), modExp_exp_1_5_1_sva,
          (COMP_LOOP_k_9_3_sva_5_0[2]), {and_dcpl_191 , and_dcpl_194 , and_dcpl_192});
      modExp_exp_1_3_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[0]), modExp_exp_1_4_1_sva,
          (COMP_LOOP_k_9_3_sva_5_0[1]), {and_dcpl_191 , and_dcpl_194 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_191 | tmp_10_lpi_4_dfm_mx0c1 | tmp_10_lpi_4_dfm_mx0c2 | tmp_10_lpi_4_dfm_mx0c3
        | tmp_10_lpi_4_dfm_mx0c4 | tmp_10_lpi_4_dfm_mx0c5 | tmp_10_lpi_4_dfm_mx0c6
        | tmp_10_lpi_4_dfm_mx0c7 ) begin
      tmp_10_lpi_4_dfm <= MUX1HOT_v_64_8_2(vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d,
          vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d,
          vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d, {COMP_LOOP_or_15_nl , COMP_LOOP_or_16_nl
          , COMP_LOOP_or_17_nl , COMP_LOOP_or_18_nl , COMP_LOOP_or_19_nl , COMP_LOOP_or_20_nl
          , COMP_LOOP_or_21_nl , COMP_LOOP_or_22_nl});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_1383_nl, mux_1360_nl, fsm_output[2]) ) begin
      COMP_LOOP_1_mul_mut <= MUX1HOT_v_64_12_2(modExp_result_sva, modulo_result_rem_cmp_z,
          modulo_qr_sva_1_mx1w1, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d,
          vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d,
          vec_rsc_0_7_i_qa_d, z_out, {COMP_LOOP_nor_97_cse , COMP_LOOP_or_26_nl ,
          COMP_LOOP_or_27_nl , COMP_LOOP_or_7_nl , COMP_LOOP_or_8_nl , COMP_LOOP_or_9_nl
          , COMP_LOOP_or_10_nl , COMP_LOOP_or_11_nl , COMP_LOOP_or_12_nl , COMP_LOOP_or_13_nl
          , COMP_LOOP_or_14_nl , nor_746_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= 12'b000000000000;
    end
    else if ( COMP_LOOP_or_3_cse ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_6_12_1;
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_77 | and_dcpl_152 | and_dcpl_90 | and_dcpl_104 | and_dcpl_109 |
        and_dcpl_116 ) begin
      COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((z_out_4[9]), (z_out_2[8]),
          and_dcpl_152);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_sva_rsp_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_1038_nl | (fsm_output[7:6]!=2'b00) | (~ not_tmp_82) ) begin
      modExp_exp_sva_rsp_1 <= operator_64_false_slc_modExp_exp_63_1_3;
    end
  end
  assign or_767_nl = (~ (fsm_output[9])) | (fsm_output[1]) | (~ (fsm_output[3]))
      | (fsm_output[5]);
  assign or_766_nl = (fsm_output[9]) | (fsm_output[1]) | (fsm_output[3]) | (~ (fsm_output[5]));
  assign mux_852_nl = MUX_s_1_2_2(or_767_nl, or_766_nl, fsm_output[6]);
  assign or_764_nl = (~ (fsm_output[6])) | (fsm_output[9]) | (~ (fsm_output[1]))
      | (~ (fsm_output[3])) | (fsm_output[5]);
  assign mux_853_nl = MUX_s_1_2_2(mux_852_nl, or_764_nl, fsm_output[7]);
  assign nor_392_nl = ~((fsm_output[8]) | mux_853_nl);
  assign nor_393_nl = ~((~ (fsm_output[8])) | (fsm_output[7]) | (~ (fsm_output[6]))
      | (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[5]));
  assign mux_854_nl = MUX_s_1_2_2(nor_392_nl, nor_393_nl, fsm_output[2]);
  assign nor_394_nl = ~((fsm_output[8]) | (fsm_output[7]) | (~ (fsm_output[6])) |
      (~ (fsm_output[9])) | (~ (fsm_output[1])) | (fsm_output[3]) | (~ (fsm_output[5])));
  assign nor_395_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[6])) | (~ (fsm_output[9]))
      | (fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[5]));
  assign nor_396_nl = ~((fsm_output[6]) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[3])
      | (~ (fsm_output[5])));
  assign mux_849_nl = MUX_s_1_2_2(nor_396_nl, nor_397_cse, fsm_output[7]);
  assign mux_850_nl = MUX_s_1_2_2(nor_395_nl, mux_849_nl, fsm_output[8]);
  assign mux_851_nl = MUX_s_1_2_2(nor_394_nl, mux_850_nl, fsm_output[2]);
  assign mux_855_nl = MUX_s_1_2_2(mux_854_nl, mux_851_nl, fsm_output[4]);
  assign mux_856_nl = MUX_s_1_2_2(mux_855_nl, nor_398_cse, fsm_output[0]);
  assign modulo_result_or_nl = and_dcpl_150 | and_dcpl_152 | mux_856_nl;
  assign mux_797_nl = MUX_s_1_2_2(or_91_cse, (~ or_90_cse), fsm_output[6]);
  assign or_733_nl = (fsm_output[8]) | nor_tmp_166;
  assign mux_796_nl = MUX_s_1_2_2((~ nor_tmp_168), or_733_nl, fsm_output[6]);
  assign mux_798_nl = MUX_s_1_2_2(mux_797_nl, mux_796_nl, and_316_cse);
  assign mux_799_nl = MUX_s_1_2_2(mux_798_nl, mux_tmp_164, fsm_output[5]);
  assign mux_792_nl = MUX_s_1_2_2((~ or_tmp_682), nor_tmp_168, fsm_output[6]);
  assign mux_791_nl = MUX_s_1_2_2(nor_tmp_166, nor_tmp_13, fsm_output[6]);
  assign mux_793_nl = MUX_s_1_2_2(mux_792_nl, mux_791_nl, fsm_output[1]);
  assign mux_789_nl = MUX_s_1_2_2((~ or_tmp_9), (fsm_output[7]), or_731_cse);
  assign mux_790_nl = MUX_s_1_2_2(mux_789_nl, mux_tmp_773, fsm_output[1]);
  assign mux_794_nl = MUX_s_1_2_2(mux_793_nl, mux_790_nl, fsm_output[2]);
  assign mux_795_nl = MUX_s_1_2_2(mux_tmp_777, (~ mux_794_nl), fsm_output[5]);
  assign mux_800_nl = MUX_s_1_2_2(mux_799_nl, mux_795_nl, fsm_output[4]);
  assign mux_783_nl = MUX_s_1_2_2(or_730_cse, or_tmp_9, fsm_output[8]);
  assign mux_784_nl = MUX_s_1_2_2((~ nor_tmp_13), mux_783_nl, fsm_output[6]);
  assign mux_781_nl = MUX_s_1_2_2(or_tmp_9, (~ (fsm_output[7])), fsm_output[8]);
  assign mux_782_nl = MUX_s_1_2_2(mux_781_nl, or_90_cse, fsm_output[6]);
  assign mux_785_nl = MUX_s_1_2_2(mux_784_nl, mux_782_nl, fsm_output[1]);
  assign mux_786_nl = MUX_s_1_2_2(mux_785_nl, mux_tmp_777, fsm_output[2]);
  assign mux_787_nl = MUX_s_1_2_2(mux_786_nl, mux_tmp_164, fsm_output[5]);
  assign or_728_nl = (fsm_output[0]) | (~ (fsm_output[7]));
  assign mux_775_nl = MUX_s_1_2_2((fsm_output[7]), or_728_nl, fsm_output[8]);
  assign mux_776_nl = MUX_s_1_2_2(mux_775_nl, or_90_cse, fsm_output[6]);
  assign mux_778_nl = MUX_s_1_2_2(mux_tmp_777, mux_776_nl, fsm_output[1]);
  assign or_727_nl = (fsm_output[6]) | or_tmp_679;
  assign mux_774_nl = MUX_s_1_2_2(or_727_nl, mux_tmp_760, fsm_output[1]);
  assign mux_779_nl = MUX_s_1_2_2(mux_778_nl, mux_774_nl, fsm_output[2]);
  assign mux_780_nl = MUX_s_1_2_2(mux_779_nl, (~ mux_tmp_773), fsm_output[5]);
  assign mux_788_nl = MUX_s_1_2_2(mux_787_nl, mux_780_nl, fsm_output[4]);
  assign mux_801_nl = MUX_s_1_2_2(mux_800_nl, mux_788_nl, fsm_output[3]);
  assign or_726_nl = (~((~ (fsm_output[6])) | (fsm_output[8]))) | (fsm_output[7]);
  assign mux_766_nl = MUX_s_1_2_2((fsm_output[7]), or_tmp_682, fsm_output[6]);
  assign mux_767_nl = MUX_s_1_2_2(or_726_nl, mux_766_nl, fsm_output[1]);
  assign mux_764_nl = MUX_s_1_2_2(or_tmp_677, or_tmp_681, fsm_output[6]);
  assign mux_763_nl = MUX_s_1_2_2(or_tmp_681, or_91_cse, fsm_output[6]);
  assign mux_765_nl = MUX_s_1_2_2(mux_764_nl, mux_763_nl, fsm_output[1]);
  assign mux_768_nl = MUX_s_1_2_2(mux_767_nl, mux_765_nl, fsm_output[2]);
  assign mux_769_nl = MUX_s_1_2_2(mux_768_nl, or_tmp_672, fsm_output[5]);
  assign mux_761_nl = MUX_s_1_2_2(mux_tmp_760, mux_tmp_164, or_722_cse);
  assign mux_762_nl = MUX_s_1_2_2(or_91_cse, mux_761_nl, fsm_output[5]);
  assign mux_770_nl = MUX_s_1_2_2(mux_769_nl, mux_762_nl, fsm_output[4]);
  assign mux_756_nl = MUX_s_1_2_2(or_tmp_679, or_tmp_677, fsm_output[6]);
  assign mux_757_nl = MUX_s_1_2_2(or_tmp_672, mux_756_nl, and_316_cse);
  assign mux_758_nl = MUX_s_1_2_2(or_91_cse, mux_757_nl, fsm_output[5]);
  assign mux_752_nl = MUX_s_1_2_2(or_91_cse, or_718_cse, fsm_output[6]);
  assign or_716_nl = (~ (fsm_output[6])) | (~ (fsm_output[0])) | (fsm_output[7]);
  assign mux_753_nl = MUX_s_1_2_2(mux_752_nl, or_716_nl, fsm_output[1]);
  assign or_715_nl = (fsm_output[8]) | (~ (fsm_output[0])) | (fsm_output[7]);
  assign mux_750_nl = MUX_s_1_2_2(or_715_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_751_nl = MUX_s_1_2_2(mux_750_nl, or_tmp_672, fsm_output[1]);
  assign mux_754_nl = MUX_s_1_2_2(mux_753_nl, mux_751_nl, fsm_output[2]);
  assign mux_755_nl = MUX_s_1_2_2(mux_754_nl, mux_tmp_164, fsm_output[5]);
  assign mux_759_nl = MUX_s_1_2_2(mux_758_nl, mux_755_nl, fsm_output[4]);
  assign mux_771_nl = MUX_s_1_2_2(mux_770_nl, mux_759_nl, fsm_output[3]);
  assign mux_802_nl = MUX_s_1_2_2(mux_801_nl, mux_771_nl, fsm_output[9]);
  assign mux_842_nl = MUX_s_1_2_2(or_831_cse, (~ (fsm_output[8])), fsm_output[7]);
  assign mux_843_nl = MUX_s_1_2_2(mux_842_nl, or_tmp_73, fsm_output[6]);
  assign mux_841_nl = MUX_s_1_2_2(or_831_cse, or_tmp_73, fsm_output[6]);
  assign mux_844_nl = MUX_s_1_2_2(mux_843_nl, mux_841_nl, fsm_output[1]);
  assign or_754_nl = (~ (fsm_output[7])) | (fsm_output[0]) | (~ (fsm_output[9]))
      | (fsm_output[8]);
  assign mux_839_nl = MUX_s_1_2_2(nand_244_cse, or_754_nl, fsm_output[6]);
  assign or_753_nl = (fsm_output[9:7]!=3'b011);
  assign mux_838_nl = MUX_s_1_2_2(mux_tmp_833, or_753_nl, fsm_output[6]);
  assign mux_840_nl = MUX_s_1_2_2(mux_839_nl, mux_838_nl, fsm_output[1]);
  assign mux_845_nl = MUX_s_1_2_2(mux_844_nl, mux_840_nl, fsm_output[2]);
  assign mux_846_nl = MUX_s_1_2_2(mux_845_nl, mux_tmp_823, fsm_output[5]);
  assign or_751_nl = and_312_cse | (fsm_output[8]);
  assign mux_834_nl = MUX_s_1_2_2(or_751_nl, mux_tmp_833, fsm_output[6]);
  assign or_748_nl = (~(nor_400_cse | (fsm_output[9]))) | (fsm_output[8]);
  assign mux_832_nl = MUX_s_1_2_2(or_748_nl, mux_417_cse, fsm_output[6]);
  assign mux_835_nl = MUX_s_1_2_2(mux_834_nl, mux_832_nl, fsm_output[1]);
  assign mux_836_nl = MUX_s_1_2_2(mux_835_nl, mux_438_cse, fsm_output[2]);
  assign mux_837_nl = MUX_s_1_2_2(mux_tmp_825, mux_836_nl, fsm_output[5]);
  assign mux_847_nl = MUX_s_1_2_2(mux_846_nl, mux_837_nl, fsm_output[4]);
  assign or_745_nl = nor_401_cse | (fsm_output[8]);
  assign mux_826_nl = MUX_s_1_2_2(or_745_nl, or_831_cse, fsm_output[7]);
  assign mux_828_nl = MUX_s_1_2_2(mux_417_cse, mux_826_nl, fsm_output[6]);
  assign mux_829_nl = MUX_s_1_2_2(mux_828_nl, mux_tmp_825, or_722_cse);
  assign mux_820_nl = MUX_s_1_2_2(not_tmp_276, or_1483_cse, or_730_cse);
  assign mux_821_nl = MUX_s_1_2_2(mux_820_nl, nand_244_cse, fsm_output[6]);
  assign mux_824_nl = MUX_s_1_2_2(mux_tmp_823, mux_821_nl, and_316_cse);
  assign mux_830_nl = MUX_s_1_2_2(mux_829_nl, mux_824_nl, fsm_output[5]);
  assign mux_815_nl = MUX_s_1_2_2(or_831_cse, or_1483_cse, fsm_output[7]);
  assign mux_816_nl = MUX_s_1_2_2(mux_815_nl, mux_tmp_814, fsm_output[6]);
  assign mux_812_nl = MUX_s_1_2_2(or_831_cse, (fsm_output[8]), fsm_output[7]);
  assign or_740_nl = (fsm_output[7]) | ((fsm_output[0]) & (fsm_output[9])) | (fsm_output[8]);
  assign mux_813_nl = MUX_s_1_2_2(mux_812_nl, or_740_nl, fsm_output[6]);
  assign mux_817_nl = MUX_s_1_2_2(mux_816_nl, mux_813_nl, fsm_output[1]);
  assign nand_127_nl = ~(or_1275_cse & (fsm_output[8]));
  assign mux_809_nl = MUX_s_1_2_2(nand_127_nl, or_tmp_73, fsm_output[7]);
  assign mux_808_nl = MUX_s_1_2_2((fsm_output[9]), or_831_cse, fsm_output[0]);
  assign or_737_nl = (fsm_output[7]) | mux_808_nl;
  assign mux_810_nl = MUX_s_1_2_2(mux_809_nl, or_737_nl, fsm_output[6]);
  assign mux_806_nl = MUX_s_1_2_2(not_tmp_276, or_tmp_73, fsm_output[7]);
  assign mux_807_nl = MUX_s_1_2_2(mux_806_nl, or_831_cse, fsm_output[6]);
  assign mux_811_nl = MUX_s_1_2_2(mux_810_nl, mux_807_nl, fsm_output[1]);
  assign mux_818_nl = MUX_s_1_2_2(mux_817_nl, mux_811_nl, fsm_output[2]);
  assign mux_819_nl = MUX_s_1_2_2(mux_818_nl, mux_438_cse, fsm_output[5]);
  assign mux_831_nl = MUX_s_1_2_2(mux_830_nl, mux_819_nl, fsm_output[4]);
  assign mux_848_nl = MUX_s_1_2_2(mux_847_nl, mux_831_nl, fsm_output[3]);
  assign nor_377_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[6]));
  assign nor_378_nl = ~(nor_379_cse | (fsm_output[9]) | (~ (fsm_output[6])));
  assign mux_875_nl = MUX_s_1_2_2(nor_378_nl, mux_tmp_865, fsm_output[1]);
  assign mux_876_nl = MUX_s_1_2_2(mux_875_nl, mux_tmp_860, fsm_output[2]);
  assign mux_877_nl = MUX_s_1_2_2(nor_377_nl, mux_876_nl, fsm_output[5]);
  assign or_789_nl = (~ (fsm_output[9])) | (fsm_output[6]);
  assign mux_872_nl = MUX_s_1_2_2(or_789_nl, or_tmp_737, fsm_output[4]);
  assign or_788_nl = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[6]));
  assign mux_873_nl = MUX_s_1_2_2(mux_872_nl, or_788_nl, and_316_cse);
  assign mux_874_nl = MUX_s_1_2_2(mux_873_nl, or_tmp_738, fsm_output[5]);
  assign mux_878_nl = MUX_s_1_2_2(mux_877_nl, (~ mux_874_nl), fsm_output[7]);
  assign nor_380_nl = ~((~((fsm_output[1]) | (fsm_output[0]) | (fsm_output[4])))
      | (~ (fsm_output[9])) | (fsm_output[6]));
  assign nor_382_nl = ~((fsm_output[4]) | (~ (fsm_output[9])) | (fsm_output[6]));
  assign mux_869_nl = MUX_s_1_2_2(nor_380_nl, nor_382_nl, fsm_output[2]);
  assign mux_870_nl = MUX_s_1_2_2(mux_869_nl, mux_tmp_860, fsm_output[5]);
  assign nor_383_nl = ~((~(and_303_cse | (fsm_output[4]))) | (fsm_output[9]) | (~
      (fsm_output[6])));
  assign mux_866_nl = MUX_s_1_2_2(mux_tmp_865, mux_tmp_860, fsm_output[1]);
  assign mux_867_nl = MUX_s_1_2_2(nor_383_nl, mux_866_nl, fsm_output[2]);
  assign mux_868_nl = MUX_s_1_2_2(mux_867_nl, (~ or_tmp_738), fsm_output[5]);
  assign mux_871_nl = MUX_s_1_2_2(mux_870_nl, mux_868_nl, fsm_output[7]);
  assign mux_879_nl = MUX_s_1_2_2(mux_878_nl, mux_871_nl, fsm_output[3]);
  assign and_304_nl = ((~ (fsm_output[4])) | (fsm_output[9])) & (fsm_output[6]);
  assign and_305_nl = (fsm_output[2:0]==3'b111);
  assign mux_861_nl = MUX_s_1_2_2(mux_tmp_860, and_304_nl, and_305_nl);
  assign and_306_nl = (fsm_output[2]) & (~((~((fsm_output[1:0]!=2'b00))) | (~ (fsm_output[4]))
      | (fsm_output[9]) | (fsm_output[6])));
  assign mux_862_nl = MUX_s_1_2_2(mux_861_nl, and_306_nl, fsm_output[5]);
  assign and_307_nl = (fsm_output[5]) & (~((or_722_cse & (fsm_output[4])) | (fsm_output[9])
      | (fsm_output[6])));
  assign mux_863_nl = MUX_s_1_2_2(mux_862_nl, and_307_nl, fsm_output[7]);
  assign and_446_nl = (~(or_722_cse & (fsm_output[4]))) & and_434_cse;
  assign nor_389_nl = ~((~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[6]));
  assign mux_858_nl = MUX_s_1_2_2(and_446_nl, nor_389_nl, fsm_output[5]);
  assign nor_390_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[1])) | (~ (fsm_output[0]))
      | (~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[6]));
  assign nor_391_nl = ~((fsm_output[4]) | (fsm_output[9]) | (fsm_output[6]));
  assign mux_857_nl = MUX_s_1_2_2(nor_390_nl, nor_391_nl, fsm_output[5]);
  assign mux_859_nl = MUX_s_1_2_2(mux_858_nl, mux_857_nl, fsm_output[7]);
  assign mux_864_nl = MUX_s_1_2_2(mux_863_nl, mux_859_nl, fsm_output[3]);
  assign mux_880_nl = MUX_s_1_2_2(mux_879_nl, mux_864_nl, fsm_output[8]);
  assign operator_64_false_1_or_2_nl = and_dcpl_71 | and_dcpl_126;
  assign or_1066_nl = (fsm_output[6:5]!=2'b00) | or_tmp_63;
  assign mux_1204_nl = MUX_s_1_2_2(or_1066_nl, mux_tmp_1203, fsm_output[7]);
  assign mux_1205_nl = MUX_s_1_2_2(mux_1204_nl, mux_tmp_1187, fsm_output[1]);
  assign mux_1210_nl = MUX_s_1_2_2(mux_1209_itm, (~ mux_1205_nl), fsm_output[8]);
  assign mux_1200_nl = MUX_s_1_2_2((~ mux_tmp_1199), or_tmp_970, fsm_output[7]);
  assign mux_1201_nl = MUX_s_1_2_2(mux_1200_nl, mux_tmp_1179, fsm_output[1]);
  assign or_1064_nl = (fsm_output[7]) | ((fsm_output[6]) & or_tmp_60);
  assign mux_1198_nl = MUX_s_1_2_2(or_1064_nl, or_tmp_993, fsm_output[1]);
  assign mux_1202_nl = MUX_s_1_2_2((~ mux_1201_nl), mux_1198_nl, fsm_output[8]);
  assign mux_1211_nl = MUX_s_1_2_2(mux_1210_nl, mux_1202_nl, fsm_output[9]);
  assign or_1063_nl = (fsm_output[5]) | and_dcpl_81;
  assign mux_1193_nl = MUX_s_1_2_2((~ and_tmp_2), or_1063_nl, fsm_output[6]);
  assign mux_1194_nl = MUX_s_1_2_2(mux_1193_nl, mux_tmp_1192, fsm_output[7]);
  assign mux_1195_nl = MUX_s_1_2_2(mux_1194_nl, mux_tmp_1191, fsm_output[1]);
  assign mux_1183_nl = MUX_s_1_2_2(or_217_cse, mux_tmp_1182, fsm_output[7]);
  assign mux_1188_nl = MUX_s_1_2_2(mux_tmp_1187, mux_1183_nl, fsm_output[1]);
  assign mux_1196_nl = MUX_s_1_2_2(mux_1195_nl, (~ mux_1188_nl), fsm_output[8]);
  assign nor_318_nl = ~((fsm_output[6]) | and_292_cse);
  assign mux_1176_nl = MUX_s_1_2_2(mux_tmp_1175, nor_318_nl, fsm_output[7]);
  assign mux_1180_nl = MUX_s_1_2_2((~ mux_tmp_1179), mux_1176_nl, fsm_output[1]);
  assign mux_1173_nl = MUX_s_1_2_2(or_tmp_993, or_857_cse, fsm_output[1]);
  assign mux_1181_nl = MUX_s_1_2_2(mux_1180_nl, mux_1173_nl, fsm_output[8]);
  assign mux_1197_nl = MUX_s_1_2_2(mux_1196_nl, mux_1181_nl, fsm_output[9]);
  assign mux_1212_nl = MUX_s_1_2_2(mux_1211_nl, mux_1197_nl, fsm_output[0]);
  assign operator_64_false_1_mux1h_nl = MUX1HOT_s_1_4_2((z_out_3[6]), modExp_exp_1_0_1_sva_1,
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm, (z_out_3[7]), {operator_64_false_1_or_2_nl
      , and_dcpl_174 , (~ mux_1212_nl) , and_dcpl_98});
  assign or_964_nl = (fsm_output[9]) | not_tmp_375;
  assign or_1052_nl = (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[4]));
  assign mux_1170_nl = MUX_s_1_2_2(or_964_nl, or_1052_nl, fsm_output[7]);
  assign or_1401_nl = (~ (fsm_output[5])) | (fsm_output[8]) | (fsm_output[6]) | mux_1170_nl;
  assign nor_320_nl = ~((fsm_output[7]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[4]));
  assign nor_321_nl = ~((~ (fsm_output[7])) | (fsm_output[9]) | not_tmp_375);
  assign mux_1169_nl = MUX_s_1_2_2(nor_320_nl, nor_321_nl, fsm_output[6]);
  assign nand_243_nl = ~((~((fsm_output[5]) | (~ (fsm_output[8])))) & mux_1169_nl);
  assign mux_1171_nl = MUX_s_1_2_2(or_1401_nl, nand_243_nl, fsm_output[3]);
  assign nor_314_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[9]))
      | (fsm_output[7]) | (fsm_output[5]));
  assign nor_315_nl = ~((fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[9]) |
      (fsm_output[7]) | (~ (fsm_output[5])));
  assign mux_1214_nl = MUX_s_1_2_2(nor_314_nl, nor_315_nl, fsm_output[4]);
  assign and_267_nl = (fsm_output[6]) & mux_1214_nl;
  assign nor_316_nl = ~((~ (fsm_output[8])) | (~ (fsm_output[9])) | (fsm_output[7])
      | (fsm_output[5]));
  assign nor_317_nl = ~((fsm_output[8]) | (fsm_output[9]) | (~ (fsm_output[7])) |
      (fsm_output[5]));
  assign mux_1213_nl = MUX_s_1_2_2(nor_316_nl, nor_317_nl, fsm_output[2]);
  assign and_268_nl = (~((fsm_output[6]) | (~ (fsm_output[4])))) & mux_1213_nl;
  assign mux_1215_nl = MUX_s_1_2_2(and_267_nl, and_268_nl, fsm_output[3]);
  assign nand_109_nl = ~((~ (fsm_output[1])) & (fsm_output[6]) & (fsm_output[9])
      & (fsm_output[4]) & (fsm_output[3]) & (fsm_output[7]) & (~ (fsm_output[5])));
  assign or_1103_nl = (fsm_output[6]) | (fsm_output[9]) | (~ (fsm_output[4])) | (fsm_output[3])
      | (fsm_output[7]) | (~ (fsm_output[5]));
  assign or_1101_nl = (fsm_output[9]) | (~ (fsm_output[4])) | (~ (fsm_output[3]))
      | (~ (fsm_output[7])) | (fsm_output[5]);
  assign mux_1260_nl = MUX_s_1_2_2(or_1101_nl, or_tmp_1034, fsm_output[6]);
  assign mux_1261_nl = MUX_s_1_2_2(or_1103_nl, mux_1260_nl, fsm_output[1]);
  assign mux_1262_nl = MUX_s_1_2_2(nand_109_nl, mux_1261_nl, fsm_output[8]);
  assign or_1098_nl = (fsm_output[9]) | (~ (fsm_output[4])) | (~ (fsm_output[3]))
      | (fsm_output[7]) | (fsm_output[5]);
  assign mux_1258_nl = MUX_s_1_2_2(or_tmp_1034, or_1098_nl, fsm_output[6]);
  assign mux_1259_nl = MUX_s_1_2_2(mux_1258_nl, nand_82_cse, fsm_output[1]);
  assign or_1100_nl = (fsm_output[8]) | mux_1259_nl;
  assign mux_1263_nl = MUX_s_1_2_2(mux_1262_nl, or_1100_nl, fsm_output[2]);
  assign and_222_nl = (~ mux_1263_nl) & (fsm_output[0]);
  assign COMP_LOOP_mux_42_nl = MUX_s_1_2_2(modExp_exp_1_0_1_sva_1, modExp_exp_1_1_1_sva,
      and_222_nl);
  assign or_1078_nl = (~ (fsm_output[9])) | (~ (fsm_output[6])) | (~ (fsm_output[1]))
      | (fsm_output[8]) | (fsm_output[5]);
  assign or_1077_nl = (fsm_output[9]) | (fsm_output[6]) | (fsm_output[1]) | (fsm_output[8])
      | (~ (fsm_output[5]));
  assign mux_1217_nl = MUX_s_1_2_2(or_1078_nl, or_1077_nl, fsm_output[4]);
  assign nor_312_nl = ~((fsm_output[7]) | mux_1217_nl);
  assign or_1074_nl = (~ (fsm_output[1])) | (fsm_output[8]) | (fsm_output[5]);
  assign or_1073_nl = (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[5]);
  assign mux_1216_nl = MUX_s_1_2_2(or_1074_nl, or_1073_nl, fsm_output[6]);
  assign nor_313_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[4])) | (fsm_output[9])
      | mux_1216_nl);
  assign mux_1218_nl = MUX_s_1_2_2(nor_312_nl, nor_313_nl, fsm_output[3]);
  assign nor_305_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[1])) | (fsm_output[9])
      | (~((fsm_output[6]) & (fsm_output[4]))));
  assign or_1109_nl = (fsm_output[9]) | (fsm_output[6]) | (fsm_output[4]);
  assign or_1108_nl = (~ (fsm_output[9])) | (fsm_output[6]) | (~ (fsm_output[4]));
  assign mux_1264_nl = MUX_s_1_2_2(or_1109_nl, or_1108_nl, fsm_output[1]);
  assign nor_306_nl = ~((fsm_output[5]) | mux_1264_nl);
  assign mux_1265_nl = MUX_s_1_2_2(nor_305_nl, nor_306_nl, fsm_output[3]);
  assign nand_242_nl = ~((fsm_output[8]) & mux_1265_nl);
  assign or_1400_nl = (fsm_output[8]) | (fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[1])
      | (~ (fsm_output[9])) | (fsm_output[6]) | (~ (fsm_output[4]));
  assign mux_1266_nl = MUX_s_1_2_2(nand_242_nl, or_1400_nl, fsm_output[7]);
  assign COMP_LOOP_mux1h_32_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_3_sva_5_0[4]), modExp_exp_1_1_1_sva,
      modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_3_sva_5_0[5]), {and_dcpl_191 , and_dcpl_177
      , (~ mux_1289_itm) , and_dcpl_192});
  assign and_259_nl = (~ (fsm_output[1])) & (fsm_output[6]) & (fsm_output[9]) & (fsm_output[4])
      & (fsm_output[3]) & (fsm_output[7]) & (~ (fsm_output[5]));
  assign nor_299_nl = ~((fsm_output[6]) | (fsm_output[9]) | (~ (fsm_output[4])) |
      (fsm_output[3]) | (fsm_output[7]) | (~ (fsm_output[5])));
  assign nor_300_nl = ~((fsm_output[9]) | (~ (fsm_output[4])) | (~ (fsm_output[3]))
      | (~ (fsm_output[7])) | (fsm_output[5]));
  assign nor_301_nl = ~((~ (fsm_output[9])) | (fsm_output[4]) | (fsm_output[3]) |
      (fsm_output[7]) | (fsm_output[5]));
  assign mux_1292_nl = MUX_s_1_2_2(nor_300_nl, nor_301_nl, fsm_output[6]);
  assign mux_1293_nl = MUX_s_1_2_2(nor_299_nl, mux_1292_nl, fsm_output[1]);
  assign mux_1294_nl = MUX_s_1_2_2(and_259_nl, mux_1293_nl, fsm_output[8]);
  assign or_1119_nl = (fsm_output[6]) | (~ (fsm_output[9])) | (fsm_output[4]) | (fsm_output[3])
      | (fsm_output[7]) | (fsm_output[5]);
  assign mux_1291_nl = MUX_s_1_2_2(or_1119_nl, nand_82_cse, fsm_output[1]);
  assign nor_302_nl = ~((fsm_output[8]) | mux_1291_nl);
  assign mux_1295_nl = MUX_s_1_2_2(mux_1294_nl, nor_302_nl, fsm_output[2]);
  assign COMP_LOOP_mux1h_46_nl = MUX1HOT_s_1_3_2(modExp_exp_1_3_1_sva, modExp_exp_1_2_1_sva,
      (COMP_LOOP_k_9_3_sva_5_0[0]), {and_dcpl_194 , (~ mux_1289_itm) , and_dcpl_192});
  assign mux_1303_nl = MUX_s_1_2_2(not_tmp_414, or_tmp_966, fsm_output[6]);
  assign mux_1304_nl = MUX_s_1_2_2(mux_1303_nl, mux_tmp_1192, fsm_output[7]);
  assign mux_1305_nl = MUX_s_1_2_2(mux_1304_nl, mux_tmp_1191, fsm_output[1]);
  assign mux_1306_nl = MUX_s_1_2_2(mux_1305_nl, (~ mux_tmp_1277), fsm_output[8]);
  assign mux_1307_nl = MUX_s_1_2_2(mux_1306_nl, mux_tmp_1272, fsm_output[9]);
  assign mux_1308_nl = MUX_s_1_2_2(mux_tmp_1288, mux_1307_nl, fsm_output[0]);
  assign COMP_LOOP_mux1h_48_nl = MUX1HOT_s_1_3_2((COMP_LOOP_k_9_3_sva_5_0[5]), modExp_exp_1_2_1_sva,
      modExp_exp_1_1_1_sva, {and_dcpl_191 , and_dcpl_194 , (~ mux_1308_nl)});
  assign nor_296_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[6]))
      | (fsm_output[0]) | not_tmp_458);
  assign nor_297_nl = ~((fsm_output[5]) | (fsm_output[7]) | (fsm_output[6]) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[4]));
  assign mux_1310_nl = MUX_s_1_2_2(nor_296_nl, nor_297_nl, fsm_output[3]);
  assign nand_192_nl = ~((fsm_output[8]) & mux_1310_nl);
  assign nand_106_nl = ~((fsm_output[6]) & (fsm_output[0]) & (~ (fsm_output[1]))
      & (fsm_output[4]));
  assign or_1140_nl = (fsm_output[6]) | (fsm_output[0]) | not_tmp_458;
  assign mux_1309_nl = MUX_s_1_2_2(nand_106_nl, or_1140_nl, fsm_output[7]);
  assign or_1300_nl = (fsm_output[8]) | (~ (fsm_output[3])) | (fsm_output[5]) | mux_1309_nl;
  assign mux_1311_nl = MUX_s_1_2_2(nand_192_nl, or_1300_nl, fsm_output[2]);
  assign or_1154_nl = (~ (fsm_output[1])) | (fsm_output[7]) | (~ (fsm_output[9]))
      | (fsm_output[4]) | (~((fsm_output[2]) & (fsm_output[6])));
  assign or_1152_nl = (fsm_output[1]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (fsm_output[6]);
  assign mux_1313_nl = MUX_s_1_2_2(or_1154_nl, or_1152_nl, fsm_output[5]);
  assign or_1308_nl = (fsm_output[8]) | mux_1313_nl;
  assign or_1150_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (~((fsm_output[4])
      & (fsm_output[2]) & (fsm_output[6])));
  assign or_1148_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[4]))
      | (fsm_output[2]) | (fsm_output[6]);
  assign mux_1312_nl = MUX_s_1_2_2(or_1150_nl, or_1148_nl, fsm_output[1]);
  assign or_1309_nl = (~ (fsm_output[8])) | (fsm_output[5]) | mux_1312_nl;
  assign mux_1314_nl = MUX_s_1_2_2(or_1308_nl, or_1309_nl, fsm_output[3]);
  assign and_54_nl = (fsm_output[8:7]==2'b11) & or_5_cse;
  assign mux_444_nl = MUX_s_1_2_2(not_tmp_129, and_54_nl, fsm_output[9]);
  assign nor_815_nl = ~((fsm_output[1:0]!=2'b01));
  assign mux_1487_nl = MUX_s_1_2_2(mux_tmp_898, and_312_cse, nor_815_nl);
  assign mux_1488_nl = MUX_s_1_2_2(mux_1487_nl, mux_tmp_1456, fsm_output[8]);
  assign mux_1489_nl = MUX_s_1_2_2(mux_1488_nl, mux_tmp_900, fsm_output[6]);
  assign mux_1484_nl = MUX_s_1_2_2(mux_tmp_898, (~ mux_936_cse), fsm_output[1]);
  assign mux_1485_nl = MUX_s_1_2_2(mux_1484_nl, or_tmp_72, fsm_output[8]);
  assign nor_835_nl = ~((fsm_output[1]) | (~ (fsm_output[9])) | (fsm_output[7]));
  assign or_1473_nl = (fsm_output[1]) | mux_1001_cse;
  assign mux_1483_nl = MUX_s_1_2_2(nor_835_nl, or_1473_nl, fsm_output[8]);
  assign mux_1486_nl = MUX_s_1_2_2(mux_1485_nl, mux_1483_nl, fsm_output[6]);
  assign mux_1490_nl = MUX_s_1_2_2(mux_1489_nl, mux_1486_nl, fsm_output[2]);
  assign mux_1478_nl = MUX_s_1_2_2(and_312_cse, mux_tmp_898, fsm_output[1]);
  assign mux_1479_nl = MUX_s_1_2_2((~ mux_1478_nl), (fsm_output[9]), fsm_output[8]);
  assign nor_836_nl = ~((~ (fsm_output[1])) | (fsm_output[9]) | (~ (fsm_output[7])));
  assign mux_1477_nl = MUX_s_1_2_2(nor_836_nl, or_tmp_783, fsm_output[8]);
  assign mux_1480_nl = MUX_s_1_2_2(mux_1479_nl, mux_1477_nl, fsm_output[6]);
  assign mux_1481_nl = MUX_s_1_2_2(mux_1480_nl, mux_928_cse, fsm_output[2]);
  assign mux_1491_nl = MUX_s_1_2_2(mux_1490_nl, mux_1481_nl, fsm_output[3]);
  assign mux_1470_nl = MUX_s_1_2_2((~ mux_tmp_898), or_tmp_783, or_1470_cse);
  assign mux_1469_nl = MUX_s_1_2_2((fsm_output[9]), and_312_cse, fsm_output[1]);
  assign mux_1471_nl = MUX_s_1_2_2(mux_1470_nl, mux_1469_nl, fsm_output[8]);
  assign mux_1467_nl = MUX_s_1_2_2(or_tmp_783, or_823_cse, fsm_output[1]);
  assign mux_1468_nl = MUX_s_1_2_2((~ or_tmp_72), mux_1467_nl, fsm_output[8]);
  assign mux_1472_nl = MUX_s_1_2_2(mux_1471_nl, mux_1468_nl, fsm_output[6]);
  assign mux_1464_nl = MUX_s_1_2_2(or_823_cse, mux_tmp_898, fsm_output[1]);
  assign and_720_nl = ((fsm_output[1]) | (fsm_output[9])) & (fsm_output[7]);
  assign mux_1465_nl = MUX_s_1_2_2(mux_1464_nl, and_720_nl, fsm_output[8]);
  assign mux_1463_nl = MUX_s_1_2_2(nor_tmp_273, mux_tmp_898, fsm_output[8]);
  assign mux_1466_nl = MUX_s_1_2_2(mux_1465_nl, mux_1463_nl, fsm_output[6]);
  assign mux_1473_nl = MUX_s_1_2_2(mux_1472_nl, mux_1466_nl, fsm_output[2]);
  assign mux_1476_nl = MUX_s_1_2_2(mux_928_cse, mux_1473_nl, fsm_output[3]);
  assign mux_1492_nl = MUX_s_1_2_2(mux_1491_nl, mux_1476_nl, fsm_output[4]);
  assign mux_1458_nl = MUX_s_1_2_2(mux_tmp_1456, (fsm_output[7]), fsm_output[8]);
  assign mux_1455_nl = MUX_s_1_2_2(mux_tmp_898, or_tmp_72, or_1470_cse);
  assign mux_1456_nl = MUX_s_1_2_2(mux_tmp_898, mux_1455_nl, fsm_output[8]);
  assign mux_1459_nl = MUX_s_1_2_2(mux_1458_nl, mux_1456_nl, fsm_output[6]);
  assign mux_1461_nl = MUX_s_1_2_2(mux_1460_cse, mux_1459_nl, and_721_cse);
  assign mux_1452_nl = MUX_s_1_2_2((~ (fsm_output[7])), nor_tmp_273, fsm_output[8]);
  assign mux_1450_nl = MUX_s_1_2_2(mux_936_cse, and_312_cse, fsm_output[1]);
  assign mux_1448_nl = MUX_s_1_2_2(or_tmp_72, (fsm_output[9]), fsm_output[1]);
  assign mux_1451_nl = MUX_s_1_2_2((~ mux_1450_nl), mux_1448_nl, fsm_output[8]);
  assign mux_1453_nl = MUX_s_1_2_2(mux_1452_nl, mux_1451_nl, fsm_output[6]);
  assign mux_1454_nl = MUX_s_1_2_2(mux_1453_nl, mux_1447_cse, or_1516_cse);
  assign mux_1462_nl = MUX_s_1_2_2(mux_1461_nl, mux_1454_nl, fsm_output[4]);
  assign mux_1493_nl = MUX_s_1_2_2(mux_1492_nl, mux_1462_nl, fsm_output[5]);
  assign nor_828_nl = ~((fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[0])) |
      (fsm_output[9]));
  assign and_715_nl = (fsm_output[6]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & (fsm_output[8])
      & (fsm_output[0]) & (fsm_output[9]);
  assign mux_1515_nl = MUX_s_1_2_2(nor_828_nl, and_715_nl, fsm_output[1]);
  assign nor_829_nl = ~((fsm_output[6]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[8]) | not_tmp_621);
  assign nor_830_nl = ~((~ (fsm_output[6])) | (fsm_output[8]) | (fsm_output[0]) |
      (~ (fsm_output[9])));
  assign mux_1514_nl = MUX_s_1_2_2(nor_829_nl, nor_830_nl, fsm_output[1]);
  assign mux_1516_nl = MUX_s_1_2_2(mux_1515_nl, mux_1514_nl, fsm_output[2]);
  assign or_1504_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[8])
      | (~ (fsm_output[0])) | (fsm_output[9]);
  assign mux_1513_nl = MUX_s_1_2_2(or_tmp_1267, or_1504_nl, fsm_output[6]);
  assign and_716_nl = (fsm_output[2:1]==2'b11) & (~ mux_1513_nl);
  assign mux_1517_nl = MUX_s_1_2_2(mux_1516_nl, and_716_nl, fsm_output[7]);
  assign mux_1509_nl = MUX_s_1_2_2((~ (fsm_output[9])), (fsm_output[9]), fsm_output[0]);
  assign mux_1510_nl = MUX_s_1_2_2(mux_1509_nl, or_tmp_1262, fsm_output[8]);
  assign and_717_nl = (fsm_output[6]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  assign mux_1511_nl = MUX_s_1_2_2(or_750_cse, mux_1510_nl, and_717_nl);
  assign or_1502_nl = (fsm_output[6]) | or_tmp_1269;
  assign mux_1512_nl = MUX_s_1_2_2(mux_1511_nl, or_1502_nl, fsm_output[1]);
  assign nor_831_nl = ~((fsm_output[7]) | (fsm_output[2]) | mux_1512_nl);
  assign mux_1518_nl = MUX_s_1_2_2(mux_1517_nl, nor_831_nl, fsm_output[3]);
  assign nand_268_nl = ~((fsm_output[1]) & (fsm_output[8]) & (~ (fsm_output[0]))
      & (fsm_output[9]));
  assign or_1498_nl = (fsm_output[1]) | (fsm_output[6]) | nor_820_cse | (fsm_output[0])
      | (~ (fsm_output[9]));
  assign mux_1507_nl = MUX_s_1_2_2(nand_268_nl, or_1498_nl, fsm_output[2]);
  assign or_1494_nl = (~ (fsm_output[6])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[8]) | not_tmp_621;
  assign mux_1505_nl = MUX_s_1_2_2(or_1494_nl, or_tmp_1274, fsm_output[1]);
  assign or_1492_nl = ((~((fsm_output[6]) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm))
      & (fsm_output[8])) | (fsm_output[0]) | (fsm_output[9]);
  assign mux_1504_nl = MUX_s_1_2_2(or_tmp_1273, or_1492_nl, fsm_output[1]);
  assign mux_1506_nl = MUX_s_1_2_2(mux_1505_nl, mux_1504_nl, fsm_output[2]);
  assign mux_1508_nl = MUX_s_1_2_2(mux_1507_nl, mux_1506_nl, fsm_output[7]);
  assign and_718_nl = (fsm_output[3]) & (~ mux_1508_nl);
  assign mux_1519_nl = MUX_s_1_2_2(mux_1518_nl, and_718_nl, fsm_output[4]);
  assign nor_832_nl = ~((~ (fsm_output[7])) | (fsm_output[2]) | (fsm_output[1]) |
      (fsm_output[6]) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[8])
      | (fsm_output[0]) | (fsm_output[9]));
  assign nor_833_nl = ~((fsm_output[7]) | (~ (fsm_output[2])) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[8])
      | not_tmp_621);
  assign mux_1502_nl = MUX_s_1_2_2(nor_832_nl, nor_833_nl, fsm_output[3]);
  assign mux_1499_nl = MUX_s_1_2_2(or_tmp_1274, or_tmp_1273, fsm_output[1]);
  assign or_1484_nl = (fsm_output[8]) | (fsm_output[0]) | (fsm_output[9]);
  assign mux_1497_nl = MUX_s_1_2_2(or_1484_nl, or_1483_cse, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1498_nl = MUX_s_1_2_2(mux_1497_nl, or_tmp_1269, fsm_output[6]);
  assign or_1485_nl = (fsm_output[1]) | mux_1498_nl;
  assign mux_1500_nl = MUX_s_1_2_2(mux_1499_nl, or_1485_nl, fsm_output[2]);
  assign or_1476_nl = (fsm_output[0]) | (~ (fsm_output[9]));
  assign mux_1494_nl = MUX_s_1_2_2(or_1476_nl, or_tmp_1262, fsm_output[8]);
  assign mux_1495_nl = MUX_s_1_2_2(or_750_cse, mux_1494_nl, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign or_1478_nl = (fsm_output[6]) | mux_1495_nl;
  assign mux_1496_nl = MUX_s_1_2_2(or_tmp_1267, or_1478_nl, fsm_output[1]);
  assign or_1481_nl = (fsm_output[2]) | mux_1496_nl;
  assign mux_1501_nl = MUX_s_1_2_2(mux_1500_nl, or_1481_nl, fsm_output[7]);
  assign nor_834_nl = ~((fsm_output[3]) | mux_1501_nl);
  assign mux_1503_nl = MUX_s_1_2_2(mux_1502_nl, nor_834_nl, fsm_output[4]);
  assign or_845_nl = (fsm_output[9:7]!=3'b000) | mux_1014_cse;
  assign or_841_nl = (~ (fsm_output[7])) | (~ (fsm_output[8])) | (~ (fsm_output[9]))
      | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[1]) | (fsm_output[4]) | (fsm_output[5]);
  assign mux_1015_nl = MUX_s_1_2_2(or_845_nl, or_841_nl, fsm_output[2]);
  assign or_1460_nl = mux_1015_nl | (fsm_output[6]);
  assign nor_825_nl = ~((fsm_output[7]) | (fsm_output[2]) | (fsm_output[9]) | mux_1014_cse);
  assign nor_826_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[2])) | (~ (fsm_output[9]))
      | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[1]) | (fsm_output[4]) | (fsm_output[5]));
  assign mux_1522_nl = MUX_s_1_2_2(nor_825_nl, nor_826_nl, fsm_output[8]);
  assign nor_827_nl = ~((~ (fsm_output[8])) | (fsm_output[7]) | (~ (fsm_output[2]))
      | (~ (fsm_output[9])) | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[1])
      | (fsm_output[4]) | (fsm_output[5]));
  assign and_286_nl = (fsm_output[3:0]==4'b1110);
  assign mux_1029_nl = MUX_s_1_2_2(nor_tmp_21, mux_tmp_229, and_286_nl);
  assign mux_1034_nl = MUX_s_1_2_2(mux_1026_cse, mux_1029_nl, fsm_output[4]);
  assign or_864_nl = (fsm_output[6:5]!=2'b00);
  assign mux_1035_nl = MUX_s_1_2_2(mux_1034_nl, nor_tmp_21, or_864_nl);
  assign nor_327_nl = ~((fsm_output[9:1]!=9'b000011011));
  assign or_982_nl = (~ (fsm_output[1])) | (fsm_output[9]) | not_tmp_29;
  assign or_980_nl = (fsm_output[1]) | (~ (fsm_output[9])) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_1131_nl = MUX_s_1_2_2(or_982_nl, or_980_nl, fsm_output[7]);
  assign nor_329_nl = ~((~ (fsm_output[4])) | (fsm_output[2]) | mux_1131_nl);
  assign mux_1132_nl = MUX_s_1_2_2(nor_365_cse, nor_329_nl, fsm_output[5]);
  assign nor_721_nl = ~((fsm_output[9]) | not_tmp_29);
  assign nor_722_nl = ~((fsm_output[9]) | (fsm_output[6]) | (fsm_output[8]));
  assign mux_55_nl = MUX_s_1_2_2(nor_721_nl, nor_722_nl, fsm_output[1]);
  assign nand_238_nl = ~((fsm_output[7]) & mux_55_nl);
  assign mux_56_nl = MUX_s_1_2_2(or_29_cse, nand_238_nl, fsm_output[2]);
  assign mux_57_nl = MUX_s_1_2_2(or_1161_cse, mux_56_nl, fsm_output[4]);
  assign nor_330_nl = ~((fsm_output[5]) | mux_57_nl);
  assign mux_1133_nl = MUX_s_1_2_2(mux_1132_nl, nor_330_nl, fsm_output[3]);
  assign mux_1134_nl = MUX_s_1_2_2(nor_327_nl, mux_1133_nl, fsm_output[0]);
  assign COMP_LOOP_COMP_LOOP_and_2_nl = (VEC_LOOP_j_sva_11_0[2:0]==3'b011);
  assign nl_COMP_LOOP_1_acc_nl = ({(z_out_8[6:0]) , 3'b000}) + ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))})
      + 10'b0000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[9:0];
  assign nor_808_nl = ~((fsm_output[9]) | (fsm_output[7]) | (fsm_output[6]) | ((fsm_output[5:4]==2'b11)
      & or_1516_cse));
  assign or_1266_nl = (fsm_output[5]) | ((fsm_output[4:3]==2'b11) & or_722_cse);
  assign or_1025_nl = (fsm_output[3]) | and_316_cse;
  assign mux_1153_nl = MUX_s_1_2_2(or_1025_nl, or_1516_cse, fsm_output[0]);
  assign nor_323_nl = ~((fsm_output[5:4]!=2'b00) | mux_1153_nl);
  assign mux_1154_nl = MUX_s_1_2_2(or_1266_nl, nor_323_nl, fsm_output[6]);
  assign or_1021_nl = (fsm_output[3:1]!=3'b000);
  assign mux_1152_nl = MUX_s_1_2_2(or_1516_cse, or_1021_nl, fsm_output[0]);
  assign or_1023_nl = (fsm_output[6:4]!=3'b000) | mux_1152_nl;
  assign mux_1155_nl = MUX_s_1_2_2(mux_1154_nl, or_1023_nl, fsm_output[7]);
  assign and_714_nl = (fsm_output[9]) & mux_1155_nl;
  assign or_1032_nl = (fsm_output[7]) | ((fsm_output[6]) & or_tmp_966);
  assign mux_1157_nl = MUX_s_1_2_2(not_tmp_390, or_1032_nl, fsm_output[8]);
  assign nand_112_nl = ~((fsm_output[6:5]==2'b11) & nor_tmp_12);
  assign mux_1159_nl = MUX_s_1_2_2(or_tmp_970, nand_112_nl, fsm_output[7]);
  assign mux_1158_nl = MUX_s_1_2_2(or_tmp_970, (~ and_433_cse), fsm_output[7]);
  assign mux_1160_nl = MUX_s_1_2_2(mux_1159_nl, mux_1158_nl, fsm_output[1]);
  assign and_208_nl = (fsm_output[7:6]==2'b11) & or_dcpl_39;
  assign and_207_nl = (fsm_output[7:6]==2'b11) & or_tmp_60;
  assign mux_1161_nl = MUX_s_1_2_2(and_208_nl, and_207_nl, fsm_output[1]);
  assign mux_1162_nl = MUX_s_1_2_2(not_tmp_390, mux_1161_nl, fsm_output[8]);
  assign or_1038_nl = (fsm_output[8:6]!=3'b000) | and_292_cse;
  assign nl_COMP_LOOP_acc_1_cse_6_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_3_sva_5_0
      , 3'b101});
  assign and_211_nl = (fsm_output[7]) & ((fsm_output[6:5]!=2'b00) | and_dcpl_75);
  assign and_210_nl = (fsm_output[7]) & ((fsm_output[6:5]!=2'b00) | and_398_cse);
  assign mux_1164_nl = MUX_s_1_2_2(and_211_nl, and_210_nl, fsm_output[1]);
  assign or_1043_nl = (fsm_output[8]) | mux_1164_nl;
  assign and_212_nl = (fsm_output[8]) & ((fsm_output[7:2]!=6'b000000));
  assign nl_COMP_LOOP_acc_1_cse_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_3_sva_5_0
      , 3'b111});
  assign or_1046_nl = (fsm_output[7]) | and_433_cse;
  assign or_1045_nl = (fsm_output[7]) | ((fsm_output[6:5]==2'b11) & or_tmp_63);
  assign mux_1167_nl = MUX_s_1_2_2(or_1046_nl, or_1045_nl, fsm_output[1]);
  assign and_214_nl = (fsm_output[8]) & mux_1167_nl;
  assign COMP_LOOP_or_15_nl = (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_191) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & tmp_10_lpi_4_dfm_mx0c1) | (COMP_LOOP_COMP_LOOP_and_5_itm & tmp_10_lpi_4_dfm_mx0c2)
      | (COMP_LOOP_COMP_LOOP_and_4_itm & tmp_10_lpi_4_dfm_mx0c3) | (COMP_LOOP_COMP_LOOP_and_32_itm
      & tmp_10_lpi_4_dfm_mx0c4) | (COMP_LOOP_COMP_LOOP_and_2_itm & tmp_10_lpi_4_dfm_mx0c5)
      | (COMP_LOOP_COMP_LOOP_and_30_itm & tmp_10_lpi_4_dfm_mx0c6) | (COMP_LOOP_COMP_LOOP_and_58_itm
      & tmp_10_lpi_4_dfm_mx0c7);
  assign COMP_LOOP_or_16_nl = (COMP_LOOP_COMP_LOOP_and_58_itm & and_dcpl_191) | (COMP_LOOP_COMP_LOOP_nor_itm
      & tmp_10_lpi_4_dfm_mx0c1) | (COMP_LOOP_COMP_LOOP_and_6_itm & tmp_10_lpi_4_dfm_mx0c2)
      | (COMP_LOOP_COMP_LOOP_and_5_itm & tmp_10_lpi_4_dfm_mx0c3) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & tmp_10_lpi_4_dfm_mx0c4) | (COMP_LOOP_COMP_LOOP_and_32_itm & tmp_10_lpi_4_dfm_mx0c5)
      | (COMP_LOOP_COMP_LOOP_and_2_itm & tmp_10_lpi_4_dfm_mx0c6) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & tmp_10_lpi_4_dfm_mx0c7);
  assign COMP_LOOP_or_17_nl = (COMP_LOOP_COMP_LOOP_and_30_itm & and_dcpl_191) | (COMP_LOOP_COMP_LOOP_and_58_itm
      & tmp_10_lpi_4_dfm_mx0c1) | (COMP_LOOP_COMP_LOOP_nor_itm & tmp_10_lpi_4_dfm_mx0c2)
      | (COMP_LOOP_COMP_LOOP_and_6_itm & tmp_10_lpi_4_dfm_mx0c3) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & tmp_10_lpi_4_dfm_mx0c4) | (COMP_LOOP_COMP_LOOP_and_4_itm & tmp_10_lpi_4_dfm_mx0c5)
      | (COMP_LOOP_COMP_LOOP_and_32_itm & tmp_10_lpi_4_dfm_mx0c6) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & tmp_10_lpi_4_dfm_mx0c7);
  assign COMP_LOOP_or_18_nl = (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_191) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & tmp_10_lpi_4_dfm_mx0c1) | (COMP_LOOP_COMP_LOOP_and_58_itm & tmp_10_lpi_4_dfm_mx0c2)
      | (COMP_LOOP_COMP_LOOP_nor_itm & tmp_10_lpi_4_dfm_mx0c3) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & tmp_10_lpi_4_dfm_mx0c4) | (COMP_LOOP_COMP_LOOP_and_5_itm & tmp_10_lpi_4_dfm_mx0c5)
      | (COMP_LOOP_COMP_LOOP_and_4_itm & tmp_10_lpi_4_dfm_mx0c6) | (COMP_LOOP_COMP_LOOP_and_32_itm
      & tmp_10_lpi_4_dfm_mx0c7);
  assign COMP_LOOP_or_19_nl = (COMP_LOOP_COMP_LOOP_and_32_itm & and_dcpl_191) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & tmp_10_lpi_4_dfm_mx0c1) | (COMP_LOOP_COMP_LOOP_and_30_itm & tmp_10_lpi_4_dfm_mx0c2)
      | (COMP_LOOP_COMP_LOOP_and_58_itm & tmp_10_lpi_4_dfm_mx0c3) | (COMP_LOOP_COMP_LOOP_nor_itm
      & tmp_10_lpi_4_dfm_mx0c4) | (COMP_LOOP_COMP_LOOP_and_6_itm & tmp_10_lpi_4_dfm_mx0c5)
      | (COMP_LOOP_COMP_LOOP_and_5_itm & tmp_10_lpi_4_dfm_mx0c6) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & tmp_10_lpi_4_dfm_mx0c7);
  assign COMP_LOOP_or_20_nl = (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_191) | (COMP_LOOP_COMP_LOOP_and_32_itm
      & tmp_10_lpi_4_dfm_mx0c1) | (COMP_LOOP_COMP_LOOP_and_2_itm & tmp_10_lpi_4_dfm_mx0c2)
      | (COMP_LOOP_COMP_LOOP_and_30_itm & tmp_10_lpi_4_dfm_mx0c3) | (COMP_LOOP_COMP_LOOP_and_58_itm
      & tmp_10_lpi_4_dfm_mx0c4) | (COMP_LOOP_COMP_LOOP_nor_itm & tmp_10_lpi_4_dfm_mx0c5)
      | (COMP_LOOP_COMP_LOOP_and_6_itm & tmp_10_lpi_4_dfm_mx0c6) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & tmp_10_lpi_4_dfm_mx0c7);
  assign COMP_LOOP_or_21_nl = (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_191) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & tmp_10_lpi_4_dfm_mx0c1) | (COMP_LOOP_COMP_LOOP_and_32_itm & tmp_10_lpi_4_dfm_mx0c2)
      | (COMP_LOOP_COMP_LOOP_and_2_itm & tmp_10_lpi_4_dfm_mx0c3) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & tmp_10_lpi_4_dfm_mx0c4) | (COMP_LOOP_COMP_LOOP_and_58_itm & tmp_10_lpi_4_dfm_mx0c5)
      | (COMP_LOOP_COMP_LOOP_nor_itm & tmp_10_lpi_4_dfm_mx0c6) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & tmp_10_lpi_4_dfm_mx0c7);
  assign COMP_LOOP_or_22_nl = (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_191) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & tmp_10_lpi_4_dfm_mx0c1) | (COMP_LOOP_COMP_LOOP_and_4_itm & tmp_10_lpi_4_dfm_mx0c2)
      | (COMP_LOOP_COMP_LOOP_and_32_itm & tmp_10_lpi_4_dfm_mx0c3) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & tmp_10_lpi_4_dfm_mx0c4) | (COMP_LOOP_COMP_LOOP_and_30_itm & tmp_10_lpi_4_dfm_mx0c5)
      | (COMP_LOOP_COMP_LOOP_and_58_itm & tmp_10_lpi_4_dfm_mx0c6) | (COMP_LOOP_COMP_LOOP_nor_itm
      & tmp_10_lpi_4_dfm_mx0c7);
  assign COMP_LOOP_or_26_nl = ((~ (modulo_result_rem_cmp_z[63])) & and_243_m1c) |
      (not_tmp_496 & (fsm_output[0]) & (~ (modulo_result_rem_cmp_z[63])));
  assign COMP_LOOP_or_27_nl = ((modulo_result_rem_cmp_z[63]) & and_243_m1c) | (not_tmp_496
      & (fsm_output[0]) & (modulo_result_rem_cmp_z[63]));
  assign COMP_LOOP_or_7_nl = (COMP_LOOP_COMP_LOOP_nor_1_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_nor_1_itm
      & and_250_m1c);
  assign COMP_LOOP_or_8_nl = (COMP_LOOP_COMP_LOOP_and_211 & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_211
      & and_250_m1c);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_COMP_LOOP_and_213 & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_213
      & and_250_m1c);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_COMP_LOOP_and_125_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_250_m1c);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_COMP_LOOP_and_215 & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_215
      & and_250_m1c);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_COMP_LOOP_and_11_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_250_m1c);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_COMP_LOOP_and_12_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_124_itm
      & and_250_m1c);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_COMP_LOOP_and_124_itm & and_244_m1c) | (COMP_LOOP_COMP_LOOP_and_125_itm
      & and_250_m1c);
  assign or_1391_nl = (~ (fsm_output[5])) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[8])
      | (~ (fsm_output[6]));
  assign or_1392_nl = (fsm_output[5]) | (fsm_output[1]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[6]);
  assign mux_71_nl = MUX_s_1_2_2(or_1391_nl, or_1392_nl, fsm_output[3]);
  assign or_1393_nl = (~ (fsm_output[3])) | (fsm_output[5]) | (~ (fsm_output[1]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_72_nl = MUX_s_1_2_2(mux_71_nl, or_1393_nl, fsm_output[7]);
  assign or_1394_nl = (fsm_output[7]) | (fsm_output[3]) | (~ (fsm_output[5])) | (~
      (fsm_output[1])) | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_73_nl = MUX_s_1_2_2(mux_72_nl, or_1394_nl, fsm_output[4]);
  assign or_1395_nl = (fsm_output[7]) | (fsm_output[3]) | (fsm_output[5]) | (~((fsm_output[1])
      & (fsm_output[9]) & (fsm_output[8]) & (fsm_output[6])));
  assign or_1396_nl = (fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[1]) | (fsm_output[9])
      | (~ (fsm_output[8])) | (fsm_output[6]);
  assign or_56_nl = (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign or_54_nl = (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[6]);
  assign mux_68_nl = MUX_s_1_2_2(or_56_nl, or_54_nl, fsm_output[1]);
  assign or_1397_nl = (~ (fsm_output[3])) | (fsm_output[5]) | mux_68_nl;
  assign mux_69_nl = MUX_s_1_2_2(or_1396_nl, or_1397_nl, fsm_output[7]);
  assign mux_70_nl = MUX_s_1_2_2(or_1395_nl, mux_69_nl, fsm_output[4]);
  assign mux_74_nl = MUX_s_1_2_2(mux_73_nl, mux_70_nl, fsm_output[2]);
  assign nor_746_nl = ~(mux_74_nl | (fsm_output[0]));
  assign mux_1379_nl = MUX_s_1_2_2((~ and_293_cse), (fsm_output[6]), fsm_output[9]);
  assign mux_1380_nl = MUX_s_1_2_2(mux_1379_nl, or_tmp_5, fsm_output[8]);
  assign mux_1381_nl = MUX_s_1_2_2(mux_1380_nl, mux_tmp_1341, fsm_output[4]);
  assign mux_1375_nl = MUX_s_1_2_2(or_tmp_1142, or_tmp_5, fsm_output[1]);
  assign mux_1376_nl = MUX_s_1_2_2(mux_1375_nl, (~ (fsm_output[6])), fsm_output[9]);
  assign mux_1377_nl = MUX_s_1_2_2(mux_1376_nl, or_119_cse, fsm_output[8]);
  assign mux_1372_nl = MUX_s_1_2_2(or_tmp_1128, or_tmp_1142, fsm_output[1]);
  assign mux_1373_nl = MUX_s_1_2_2(mux_tmp_1353, mux_1372_nl, fsm_output[9]);
  assign mux_1371_nl = MUX_s_1_2_2((~ mux_tmp_1355), or_857_cse, fsm_output[9]);
  assign mux_1374_nl = MUX_s_1_2_2(mux_1373_nl, mux_1371_nl, fsm_output[8]);
  assign mux_1378_nl = MUX_s_1_2_2(mux_1377_nl, mux_1374_nl, fsm_output[4]);
  assign mux_1382_nl = MUX_s_1_2_2(mux_1381_nl, mux_1378_nl, fsm_output[5]);
  assign and_253_nl = (fsm_output[1]) & (fsm_output[7]) & (fsm_output[0]) & (fsm_output[6]);
  assign mux_1367_nl = MUX_s_1_2_2(and_253_nl, mux_tmp_1345, fsm_output[9]);
  assign mux_1368_nl = MUX_s_1_2_2((~ mux_1367_nl), mux_tmp_1348, fsm_output[8]);
  assign or_1207_nl = (fsm_output[7]) | (fsm_output[0]) | (fsm_output[6]);
  assign mux_1364_nl = MUX_s_1_2_2((~ mux_tmp_1329), or_1207_nl, fsm_output[1]);
  assign mux_1365_nl = MUX_s_1_2_2((~ and_293_cse), mux_1364_nl, fsm_output[9]);
  assign or_1206_nl = (fsm_output[7]) | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_1362_nl = MUX_s_1_2_2(or_tmp_1137, or_1206_nl, fsm_output[1]);
  assign mux_1363_nl = MUX_s_1_2_2(or_tmp_13, mux_1362_nl, fsm_output[9]);
  assign mux_1366_nl = MUX_s_1_2_2(mux_1365_nl, mux_1363_nl, fsm_output[8]);
  assign mux_1369_nl = MUX_s_1_2_2(mux_1368_nl, mux_1366_nl, fsm_output[4]);
  assign mux_1361_nl = MUX_s_1_2_2(mux_tmp_1351, mux_tmp_1332, fsm_output[4]);
  assign mux_1370_nl = MUX_s_1_2_2(mux_1369_nl, mux_1361_nl, fsm_output[5]);
  assign mux_1383_nl = MUX_s_1_2_2(mux_1382_nl, mux_1370_nl, fsm_output[3]);
  assign mux_1356_nl = MUX_s_1_2_2(and_293_cse, mux_tmp_1355, fsm_output[9]);
  assign or_1201_nl = (~ (fsm_output[1])) | (fsm_output[7]) | nand_240_cse;
  assign mux_1354_nl = MUX_s_1_2_2(mux_tmp_1353, or_1201_nl, fsm_output[9]);
  assign mux_1357_nl = MUX_s_1_2_2((~ mux_1356_nl), mux_1354_nl, fsm_output[8]);
  assign mux_1358_nl = MUX_s_1_2_2(mux_1357_nl, mux_tmp_1341, fsm_output[4]);
  assign mux_1346_nl = MUX_s_1_2_2((~ mux_tmp_1345), or_857_cse, fsm_output[9]);
  assign mux_1349_nl = MUX_s_1_2_2(mux_tmp_1348, mux_1346_nl, fsm_output[8]);
  assign mux_1352_nl = MUX_s_1_2_2(mux_tmp_1351, mux_1349_nl, fsm_output[4]);
  assign mux_1359_nl = MUX_s_1_2_2(mux_1358_nl, mux_1352_nl, fsm_output[5]);
  assign or_1196_nl = (~ (fsm_output[7])) | (fsm_output[0]) | (~ (fsm_output[6]));
  assign mux_1337_nl = MUX_s_1_2_2(or_1196_nl, or_tmp_1128, fsm_output[1]);
  assign nand_98_nl = ~(((fsm_output[1]) | (~ (fsm_output[7])) | (fsm_output[0]))
      & (fsm_output[6]));
  assign mux_1338_nl = MUX_s_1_2_2(mux_1337_nl, nand_98_nl, fsm_output[9]);
  assign nand_99_nl = ~((fsm_output[7]) & (fsm_output[0]) & (fsm_output[6]));
  assign or_1191_nl = nor_400_cse | (fsm_output[6]);
  assign mux_1336_nl = MUX_s_1_2_2(nand_99_nl, or_1191_nl, fsm_output[1]);
  assign or_1192_nl = (fsm_output[9]) | mux_1336_nl;
  assign mux_1339_nl = MUX_s_1_2_2(mux_1338_nl, or_1192_nl, fsm_output[8]);
  assign mux_1342_nl = MUX_s_1_2_2(mux_tmp_1341, mux_1339_nl, fsm_output[4]);
  assign nand_183_nl = ~((~((fsm_output[1]) & (fsm_output[7]) & (fsm_output[0])))
      & (fsm_output[6]));
  assign mux_1333_nl = MUX_s_1_2_2(or_tmp_5, nand_183_nl, fsm_output[9]);
  assign mux_1334_nl = MUX_s_1_2_2(mux_1333_nl, or_119_cse, fsm_output[8]);
  assign mux_1335_nl = MUX_s_1_2_2(mux_1334_nl, mux_tmp_1332, fsm_output[4]);
  assign mux_1343_nl = MUX_s_1_2_2(mux_1342_nl, mux_1335_nl, fsm_output[5]);
  assign mux_1360_nl = MUX_s_1_2_2(mux_1359_nl, mux_1343_nl, fsm_output[3]);
  assign mux_1038_nl = MUX_s_1_2_2(mux_tmp_1037, mux_tmp_81, fsm_output[1]);
  assign and_725_nl = and_dcpl_223 & and_dcpl_218 & (~ (fsm_output[4])) & (fsm_output[0]);
  assign and_726_nl = and_dcpl_223 & and_dcpl_218 & nor_379_cse;
  assign modExp_while_mux1h_3_nl = MUX1HOT_v_64_4_2(modExp_base_sva, modExp_result_sva,
      COMP_LOOP_1_mul_mut, operator_64_false_acc_mut_63_0, {and_725_nl , and_726_nl
      , not_tmp_519 , not_tmp_524});
  assign modExp_while_or_2_nl = not_tmp_519 | not_tmp_524;
  assign modExp_while_mux_1_nl = MUX_v_64_2_2(modExp_base_sva, COMP_LOOP_1_mul_mut,
      modExp_while_or_2_nl);
  assign nl_z_out = modExp_while_mux1h_3_nl * modExp_while_mux_1_nl;
  assign z_out = nl_z_out[63:0];
  assign and_727_nl = (fsm_output[9:7]==3'b111) & nor_797_cse & (~ (fsm_output[4]))
      & (fsm_output[2]) & (~ (fsm_output[1])) & and_dcpl_313;
  assign COMP_LOOP_mux_45_nl = MUX_v_10_2_2(({1'b0 , COMP_LOOP_k_9_3_sva_5_0 , 3'b011}),
      STAGE_LOOP_lshift_psp_sva, and_727_nl);
  assign nl_z_out_1 = conv_u2u_12_13(VEC_LOOP_j_sva_11_0) + conv_u2u_10_13(COMP_LOOP_mux_45_nl);
  assign z_out_1 = nl_z_out_1[12:0];
  assign COMP_LOOP_mux_46_nl = MUX_v_56_2_2((tmp_10_lpi_4_dfm[63:8]), (p_sva[63:8]),
      and_dcpl_256);
  assign COMP_LOOP_COMP_LOOP_or_6_nl = MUX_v_56_2_2(COMP_LOOP_mux_46_nl, 56'b11111111111111111111111111111111111111111111111111111111,
      COMP_LOOP_or_39_itm);
  assign COMP_LOOP_mux1h_268_nl = MUX1HOT_s_1_4_2((tmp_10_lpi_4_dfm[7]), (~ modExp_exp_1_7_1_sva),
      (p_sva[7]), (~ modExp_exp_1_1_1_sva), {and_dcpl_246 , and_dcpl_247 , and_dcpl_256
      , and_dcpl_262});
  assign COMP_LOOP_mux1h_269_nl = MUX1HOT_s_1_4_2((tmp_10_lpi_4_dfm[6]), (~ modExp_exp_1_6_1_sva),
      (p_sva[6]), (~ modExp_exp_1_7_1_sva), {and_dcpl_246 , and_dcpl_247 , and_dcpl_256
      , and_dcpl_262});
  assign COMP_LOOP_mux1h_270_nl = MUX1HOT_s_1_4_2((tmp_10_lpi_4_dfm[5]), (~ modExp_exp_1_5_1_sva),
      (p_sva[5]), (~ modExp_exp_1_6_1_sva), {and_dcpl_246 , and_dcpl_247 , and_dcpl_256
      , and_dcpl_262});
  assign COMP_LOOP_mux1h_271_nl = MUX1HOT_s_1_4_2((tmp_10_lpi_4_dfm[4]), (~ modExp_exp_1_4_1_sva),
      (p_sva[4]), (~ modExp_exp_1_5_1_sva), {and_dcpl_246 , and_dcpl_247 , and_dcpl_256
      , and_dcpl_262});
  assign COMP_LOOP_mux1h_272_nl = MUX1HOT_s_1_4_2((tmp_10_lpi_4_dfm[3]), (~ modExp_exp_1_3_1_sva),
      (p_sva[3]), (~ modExp_exp_1_4_1_sva), {and_dcpl_246 , and_dcpl_247 , and_dcpl_256
      , and_dcpl_262});
  assign COMP_LOOP_mux1h_273_nl = MUX1HOT_s_1_4_2((tmp_10_lpi_4_dfm[2]), (~ modExp_exp_1_2_1_sva),
      (p_sva[2]), (~ modExp_exp_1_3_1_sva), {and_dcpl_246 , and_dcpl_247 , and_dcpl_256
      , and_dcpl_262});
  assign COMP_LOOP_mux1h_274_nl = MUX1HOT_s_1_4_2((tmp_10_lpi_4_dfm[1]), (~ modExp_exp_1_1_1_sva),
      (p_sva[1]), (~ modExp_exp_1_2_1_sva), {and_dcpl_246 , and_dcpl_247 , and_dcpl_256
      , and_dcpl_262});
  assign COMP_LOOP_mux1h_275_nl = MUX1HOT_s_1_3_2((tmp_10_lpi_4_dfm[0]), (~ modExp_exp_1_0_1_sva_1),
      (p_sva[0]), {and_dcpl_246 , COMP_LOOP_or_39_itm , and_dcpl_256});
  assign COMP_LOOP_or_48_nl = (~(and_dcpl_247 | and_dcpl_256 | and_dcpl_262)) | and_dcpl_246;
  assign COMP_LOOP_mux_47_nl = MUX_v_64_2_2(modulo_result_mux_1_cse, 64'b1111111111111111111111111111111111111111111111111111111111111110,
      COMP_LOOP_or_39_itm);
  assign COMP_LOOP_not_199_nl = ~ and_dcpl_256;
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nand_1_nl = ~(MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
      COMP_LOOP_mux_47_nl, COMP_LOOP_not_199_nl));
  assign nl_acc_1_nl = conv_u2u_65_66({COMP_LOOP_COMP_LOOP_or_6_nl , COMP_LOOP_mux1h_268_nl
      , COMP_LOOP_mux1h_269_nl , COMP_LOOP_mux1h_270_nl , COMP_LOOP_mux1h_271_nl
      , COMP_LOOP_mux1h_272_nl , COMP_LOOP_mux1h_273_nl , COMP_LOOP_mux1h_274_nl
      , COMP_LOOP_mux1h_275_nl , COMP_LOOP_or_48_nl}) + conv_s2u_65_66({COMP_LOOP_COMP_LOOP_COMP_LOOP_nand_1_nl
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[65:0];
  assign z_out_2 = readslicef_66_65_1(acc_1_nl);
  assign operator_64_false_1_operator_64_false_1_or_2_nl = operator_64_false_1_nor_1_itm
      | and_dcpl_277;
  assign operator_64_false_1_mux_1_nl = MUX_s_1_2_2((~ (STAGE_LOOP_lshift_psp_sva[9])),
      (STAGE_LOOP_lshift_psp_sva[9]), and_dcpl_289);
  assign operator_64_false_1_operator_64_false_1_or_3_nl = operator_64_false_1_mux_1_nl
      | and_dcpl_271 | and_dcpl_284;
  assign operator_64_false_1_mux1h_3_nl = MUX1HOT_v_6_4_2((~ COMP_LOOP_k_9_3_sva_5_0),
      (~ (STAGE_LOOP_lshift_psp_sva[8:3])), (~ (STAGE_LOOP_lshift_psp_sva[9:4])),
      (STAGE_LOOP_lshift_psp_sva[8:3]), {and_dcpl_271 , and_dcpl_277 , and_dcpl_284
      , and_dcpl_289});
  assign operator_64_false_1_or_4_nl = (~(and_dcpl_271 | and_dcpl_289)) | and_dcpl_277
      | and_dcpl_284;
  assign operator_64_false_1_operator_64_false_1_and_1_nl = (COMP_LOOP_k_9_3_sva_5_0[5])
      & operator_64_false_1_nor_1_itm;
  assign operator_64_false_1_or_5_nl = and_dcpl_284 | and_dcpl_289;
  assign operator_64_false_1_mux1h_4_nl = MUX1HOT_v_6_3_2(6'b000001, ({(COMP_LOOP_k_9_3_sva_5_0[4:0])
      , 1'b0}), COMP_LOOP_k_9_3_sva_5_0, {and_dcpl_271 , and_dcpl_277 , operator_64_false_1_or_5_nl});
  assign nl_acc_2_nl = ({operator_64_false_1_operator_64_false_1_or_2_nl , operator_64_false_1_operator_64_false_1_or_3_nl
      , operator_64_false_1_mux1h_3_nl , operator_64_false_1_or_4_nl}) + conv_u2u_8_9({operator_64_false_1_operator_64_false_1_and_1_nl
      , operator_64_false_1_mux1h_4_nl , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[8:0];
  assign z_out_3 = readslicef_9_8_1(acc_2_nl);
  assign COMP_LOOP_COMP_LOOP_or_7_nl = (VEC_LOOP_j_sva_11_0[11]) | and_dcpl_305 |
      and_dcpl_312 | and_dcpl_318 | and_dcpl_326 | and_dcpl_330;
  assign COMP_LOOP_COMP_LOOP_mux_9_nl = MUX_v_9_2_2((VEC_LOOP_j_sva_11_0[10:2]),
      (~ (STAGE_LOOP_lshift_psp_sva[9:1])), COMP_LOOP_or_43_itm);
  assign COMP_LOOP_or_49_nl = (~ and_dcpl_298) | and_dcpl_305 | and_dcpl_312 | and_dcpl_318
      | and_dcpl_326 | and_dcpl_330;
  assign COMP_LOOP_COMP_LOOP_mux_10_nl = MUX_v_6_2_2(({2'b00 , (COMP_LOOP_k_9_3_sva_5_0[5:2])}),
      COMP_LOOP_k_9_3_sva_5_0, COMP_LOOP_or_43_itm);
  assign COMP_LOOP_COMP_LOOP_or_8_nl = ((COMP_LOOP_k_9_3_sva_5_0[1]) & (~(and_dcpl_305
      | and_dcpl_312))) | and_dcpl_318 | and_dcpl_326 | and_dcpl_330;
  assign COMP_LOOP_COMP_LOOP_or_9_nl = ((COMP_LOOP_k_9_3_sva_5_0[0]) & (~(and_dcpl_305
      | and_dcpl_318 | and_dcpl_326))) | and_dcpl_312 | and_dcpl_330;
  assign COMP_LOOP_COMP_LOOP_or_10_nl = (~(and_dcpl_312 | and_dcpl_318 | and_dcpl_330))
      | and_dcpl_298 | and_dcpl_305 | and_dcpl_326;
  assign nl_acc_3_nl = ({COMP_LOOP_COMP_LOOP_or_7_nl , COMP_LOOP_COMP_LOOP_mux_9_nl
      , COMP_LOOP_or_49_nl}) + conv_u2u_10_11({COMP_LOOP_COMP_LOOP_mux_10_nl , COMP_LOOP_COMP_LOOP_or_8_nl
      , COMP_LOOP_COMP_LOOP_or_9_nl , COMP_LOOP_COMP_LOOP_or_10_nl , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[10:0];
  assign z_out_4 = readslicef_11_10_1(acc_3_nl);
  assign and_728_nl = (fsm_output[9:7]==3'b001) & and_dcpl_280 & (~ (fsm_output[2]))
      & (~ (fsm_output[4])) & (~ (fsm_output[1])) & and_dcpl_278;
  assign and_729_nl = and_dcpl_91 & (~ (fsm_output[7])) & and_dcpl_267 & and_dcpl_342
      & and_dcpl_313;
  assign and_730_nl = and_dcpl_91 & (fsm_output[7]) & and_dcpl_280 & (fsm_output[2])
      & (fsm_output[4]) & (~ (fsm_output[1])) & and_dcpl_313;
  assign and_731_nl = and_dcpl_360 & nor_797_cse & and_dcpl_355 & (fsm_output[1])
      & and_dcpl_313;
  assign and_732_nl = and_dcpl_360 & and_dcpl_267 & and_dcpl_291 & (~ (fsm_output[1]))
      & and_dcpl_278;
  assign and_733_nl = and_dcpl_359 & (fsm_output[7]) & and_dcpl_280 & and_dcpl_342
      & and_dcpl_278;
  assign COMP_LOOP_mux1h_276_nl = MUX1HOT_v_3_6_2(3'b001, 3'b010, 3'b011, 3'b100,
      3'b101, 3'b110, {and_728_nl , and_729_nl , and_730_nl , and_731_nl , and_732_nl
      , and_733_nl});
  assign and_734_nl = (fsm_output[9:7]==3'b110) & nor_797_cse & and_dcpl_355 & (~
      (fsm_output[1])) & and_dcpl_278;
  assign COMP_LOOP_or_50_nl = MUX_v_3_2_2(COMP_LOOP_mux1h_276_nl, 3'b111, and_734_nl);
  assign nl_COMP_LOOP_acc_59_nl = STAGE_LOOP_lshift_psp_sva + conv_u2u_9_10({COMP_LOOP_k_9_3_sva_5_0
      , COMP_LOOP_or_50_nl});
  assign COMP_LOOP_acc_59_nl = nl_COMP_LOOP_acc_59_nl[9:0];
  assign COMP_LOOP_or_51_nl = (and_dcpl_309 & (~ (fsm_output[8])) & and_dcpl_280
      & (~((fsm_output[2]) | (fsm_output[4]) | (fsm_output[1]))) & and_dcpl_278)
      | ((fsm_output[9:7]==3'b010) & and_dcpl_267 & and_dcpl_342 & and_dcpl_313)
      | and_dcpl_318 | (and_dcpl_411 & nor_797_cse & and_dcpl_355 & (fsm_output[1])
      & and_dcpl_313) | (and_dcpl_411 & and_dcpl_267 & and_dcpl_291 & (~ (fsm_output[1]))
      & and_dcpl_278) | ((fsm_output[9:7]==3'b101) & and_dcpl_280 & and_dcpl_342
      & and_dcpl_278) | (and_dcpl_410 & (fsm_output[8]) & nor_797_cse & and_dcpl_355
      & (~ (fsm_output[1])) & and_dcpl_278);
  assign COMP_LOOP_COMP_LOOP_mux_11_nl = MUX_v_10_2_2(({(z_out_3[6:0]) , (STAGE_LOOP_lshift_psp_sva[2:0])}),
      COMP_LOOP_acc_59_nl, COMP_LOOP_or_51_nl);
  assign nl_COMP_LOOP_acc_58_nl = conv_u2u_12_13(VEC_LOOP_j_sva_11_0) + conv_u2u_10_13(COMP_LOOP_COMP_LOOP_mux_11_nl);
  assign COMP_LOOP_acc_58_nl = nl_COMP_LOOP_acc_58_nl[12:0];
  assign z_out_6_12_1 = readslicef_13_12_1(COMP_LOOP_acc_58_nl);
  assign COMP_LOOP_not_200_nl = ~ and_dcpl_442;
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_2_nl = ~(MUX_v_53_2_2((operator_66_true_div_cmp_z[63:11]),
      53'b11111111111111111111111111111111111111111111111111111, COMP_LOOP_not_200_nl));
  assign COMP_LOOP_mux_48_nl = MUX_v_11_2_2((VEC_LOOP_j_sva_11_0[11:1]), (~ (operator_66_true_div_cmp_z[10:0])),
      and_dcpl_442);
  assign not_2902_nl = ~ and_dcpl_442;
  assign COMP_LOOP_COMP_LOOP_and_220_nl = MUX_v_6_2_2(6'b000000, COMP_LOOP_k_9_3_sva_5_0,
      not_2902_nl);
  assign nl_z_out_7 = ({and_dcpl_442 , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_2_nl , COMP_LOOP_mux_48_nl})
      + conv_u2u_8_65({COMP_LOOP_COMP_LOOP_and_220_nl , (~ and_dcpl_442) , 1'b1});
  assign z_out_7 = nl_z_out_7[64:0];
  assign COMP_LOOP_COMP_LOOP_or_11_nl = (~(and_dcpl_451 | and_dcpl_460)) | and_dcpl_467;
  assign COMP_LOOP_or_52_nl = and_dcpl_451 | and_dcpl_460;
  assign COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_3_nl = ~(MUX_v_52_2_2((operator_64_false_slc_modExp_exp_63_1_itm[62:11]),
      52'b1111111111111111111111111111111111111111111111111111, COMP_LOOP_or_52_nl));
  assign COMP_LOOP_mux1h_277_nl = MUX1HOT_v_11_3_2((VEC_LOOP_j_sva_11_0[11:1]), ({5'b00000
      , COMP_LOOP_k_9_3_sva_5_0}), (~ (operator_64_false_slc_modExp_exp_63_1_itm[10:0])),
      {and_dcpl_451 , and_dcpl_460 , and_dcpl_467});
  assign COMP_LOOP_nor_109_nl = ~(and_dcpl_460 | and_dcpl_467);
  assign COMP_LOOP_COMP_LOOP_and_221_nl = MUX_v_6_2_2(6'b000000, COMP_LOOP_k_9_3_sva_5_0,
      COMP_LOOP_nor_109_nl);
  assign nl_z_out_8 = ({COMP_LOOP_COMP_LOOP_or_11_nl , COMP_LOOP_COMP_LOOP_COMP_LOOP_nor_3_nl
      , COMP_LOOP_mux1h_277_nl}) + conv_u2u_8_64({COMP_LOOP_COMP_LOOP_and_221_nl
      , 2'b01});
  assign z_out_8 = nl_z_out_8[63:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_6_2;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [5:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    result = result | ( input_4 & {3{sel[4]}});
    result = result | ( input_5 & {3{sel[5]}});
    MUX1HOT_v_3_6_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_12_2;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [11:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    MUX1HOT_v_64_12_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_5_2;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [4:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    MUX1HOT_v_64_5_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_8_2;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [7:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    MUX1HOT_v_64_8_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_11_2;
    input [8:0] input_10;
    input [8:0] input_9;
    input [8:0] input_8;
    input [8:0] input_7;
    input [8:0] input_6;
    input [8:0] input_5;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [10:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    result = result | ( input_4 & {9{sel[4]}});
    result = result | ( input_5 & {9{sel[5]}});
    result = result | ( input_6 & {9{sel[6]}});
    result = result | ( input_7 & {9{sel[7]}});
    result = result | ( input_8 & {9{sel[8]}});
    result = result | ( input_9 & {9{sel[9]}});
    result = result | ( input_10 & {9{sel[10]}});
    MUX1HOT_v_9_11_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [51:0] MUX_v_52_2_2;
    input [51:0] input_0;
    input [51:0] input_1;
    input [0:0] sel;
    reg [51:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_52_2_2 = result;
  end
  endfunction


  function automatic [52:0] MUX_v_53_2_2;
    input [52:0] input_0;
    input [52:0] input_1;
    input [0:0] sel;
    reg [52:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_53_2_2 = result;
  end
  endfunction


  function automatic [55:0] MUX_v_56_2_2;
    input [55:0] input_0;
    input [55:0] input_1;
    input [0:0] sel;
    reg [55:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_56_2_2 = result;
  end
  endfunction


  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [64:0] readslicef_66_65_1;
    input [65:0] vector;
    reg [65:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_66_65_1 = tmp[64:0];
  end
  endfunction


  function automatic [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction


  function automatic [65:0] conv_s2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_s2u_65_66 = {vector[64], vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_6_9 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_9 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [63:0] conv_u2u_8_64 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_64 = {{56{1'b0}}, vector};
  end
  endfunction


  function automatic [64:0] conv_u2u_8_65 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_65 = {{57{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_10_13 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_13 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [65:0] conv_u2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_u2u_65_66 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      vec_rsc_0_2_adra, vec_rsc_0_2_da, vec_rsc_0_2_wea, vec_rsc_0_2_qa, vec_rsc_triosy_0_2_lz,
      vec_rsc_0_3_adra, vec_rsc_0_3_da, vec_rsc_0_3_wea, vec_rsc_0_3_qa, vec_rsc_triosy_0_3_lz,
      vec_rsc_0_4_adra, vec_rsc_0_4_da, vec_rsc_0_4_wea, vec_rsc_0_4_qa, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_adra, vec_rsc_0_5_da, vec_rsc_0_5_wea, vec_rsc_0_5_qa, vec_rsc_triosy_0_5_lz,
      vec_rsc_0_6_adra, vec_rsc_0_6_da, vec_rsc_0_6_wea, vec_rsc_0_6_qa, vec_rsc_triosy_0_6_lz,
      vec_rsc_0_7_adra, vec_rsc_0_7_da, vec_rsc_0_7_wea, vec_rsc_0_7_qa, vec_rsc_triosy_0_7_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [8:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [8:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  output [8:0] vec_rsc_0_2_adra;
  output [63:0] vec_rsc_0_2_da;
  output vec_rsc_0_2_wea;
  input [63:0] vec_rsc_0_2_qa;
  output vec_rsc_triosy_0_2_lz;
  output [8:0] vec_rsc_0_3_adra;
  output [63:0] vec_rsc_0_3_da;
  output vec_rsc_0_3_wea;
  input [63:0] vec_rsc_0_3_qa;
  output vec_rsc_triosy_0_3_lz;
  output [8:0] vec_rsc_0_4_adra;
  output [63:0] vec_rsc_0_4_da;
  output vec_rsc_0_4_wea;
  input [63:0] vec_rsc_0_4_qa;
  output vec_rsc_triosy_0_4_lz;
  output [8:0] vec_rsc_0_5_adra;
  output [63:0] vec_rsc_0_5_da;
  output vec_rsc_0_5_wea;
  input [63:0] vec_rsc_0_5_qa;
  output vec_rsc_triosy_0_5_lz;
  output [8:0] vec_rsc_0_6_adra;
  output [63:0] vec_rsc_0_6_da;
  output vec_rsc_0_6_wea;
  input [63:0] vec_rsc_0_6_qa;
  output vec_rsc_triosy_0_6_lz;
  output [8:0] vec_rsc_0_7_adra;
  output [63:0] vec_rsc_0_7_da;
  output vec_rsc_0_7_wea;
  input [63:0] vec_rsc_0_7_qa;
  output vec_rsc_triosy_0_7_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_qa_d;
  wire vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_qa_d;
  wire vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_qa_d;
  wire vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_qa_d;
  wire vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_qa_d;
  wire vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_qa_d;
  wire vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [8:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;
  wire vec_rsc_0_2_i_wea_d_iff;
  wire vec_rsc_0_3_i_wea_d_iff;
  wire vec_rsc_0_4_i_wea_d_iff;
  wire vec_rsc_0_5_i_wea_d_iff;
  wire vec_rsc_0_6_i_wea_d_iff;
  wire vec_rsc_0_7_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_9_64_512_512_64_1_gen vec_rsc_0_0_i
      (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_9_64_512_512_64_1_gen vec_rsc_0_1_i
      (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_9_64_512_512_64_1_gen vec_rsc_0_2_i
      (
      .qa(vec_rsc_0_2_qa),
      .wea(vec_rsc_0_2_wea),
      .da(vec_rsc_0_2_da),
      .adra(vec_rsc_0_2_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_2_i_qa_d),
      .wea_d(vec_rsc_0_2_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_9_64_512_512_64_1_gen vec_rsc_0_3_i
      (
      .qa(vec_rsc_0_3_qa),
      .wea(vec_rsc_0_3_wea),
      .da(vec_rsc_0_3_da),
      .adra(vec_rsc_0_3_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_3_i_qa_d),
      .wea_d(vec_rsc_0_3_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_9_64_512_512_64_1_gen vec_rsc_0_4_i
      (
      .qa(vec_rsc_0_4_qa),
      .wea(vec_rsc_0_4_wea),
      .da(vec_rsc_0_4_da),
      .adra(vec_rsc_0_4_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_4_i_qa_d),
      .wea_d(vec_rsc_0_4_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_9_64_512_512_64_1_gen vec_rsc_0_5_i
      (
      .qa(vec_rsc_0_5_qa),
      .wea(vec_rsc_0_5_wea),
      .da(vec_rsc_0_5_da),
      .adra(vec_rsc_0_5_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_5_i_qa_d),
      .wea_d(vec_rsc_0_5_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_9_64_512_512_64_1_gen
      vec_rsc_0_6_i (
      .qa(vec_rsc_0_6_qa),
      .wea(vec_rsc_0_6_wea),
      .da(vec_rsc_0_6_da),
      .adra(vec_rsc_0_6_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_6_i_qa_d),
      .wea_d(vec_rsc_0_6_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_9_64_512_512_64_1_gen
      vec_rsc_0_7_i (
      .qa(vec_rsc_0_7_qa),
      .wea(vec_rsc_0_7_wea),
      .da(vec_rsc_0_7_da),
      .adra(vec_rsc_0_7_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_7_i_qa_d),
      .wea_d(vec_rsc_0_7_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_wea_d_iff)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_qa_d(vec_rsc_0_2_i_qa_d),
      .vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_qa_d(vec_rsc_0_3_i_qa_d),
      .vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_qa_d(vec_rsc_0_4_i_qa_d),
      .vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_qa_d(vec_rsc_0_5_i_qa_d),
      .vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_qa_d(vec_rsc_0_6_i_qa_d),
      .vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_qa_d(vec_rsc_0_7_i_qa_d),
      .vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff),
      .vec_rsc_0_2_i_wea_d_pff(vec_rsc_0_2_i_wea_d_iff),
      .vec_rsc_0_3_i_wea_d_pff(vec_rsc_0_3_i_wea_d_iff),
      .vec_rsc_0_4_i_wea_d_pff(vec_rsc_0_4_i_wea_d_iff),
      .vec_rsc_0_5_i_wea_d_pff(vec_rsc_0_5_i_wea_d_iff),
      .vec_rsc_0_6_i_wea_d_pff(vec_rsc_0_6_i_wea_d_iff),
      .vec_rsc_0_7_i_wea_d_pff(vec_rsc_0_7_i_wea_d_iff)
    );
endmodule



